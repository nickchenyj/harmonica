module harmonica(phi,
                   AluDivFinish,
                   AluDivQ,
                   AluDivR,
                   FpuBasicFinish,
                   FpuBasicRes,
                   FpuMultFinish,
                   FpuMultRes,
                   AluDivA,
                   AluDivB,
                   AluDivStall,
                   AluDivValid,
                   FpuBasicA,
                   FpuBasicB,
                   FpuBasicOp,
                   FpuBasicStall,
                   FpuBasicValid,
                   FpuMultA,
                   FpuMultB,
                   FpuMultOp,
                   FpuMultStall,
                   FpuMultValid,
                   char_out,
                   char_out_val,
                   reg00,
                   reg01,
                   reg02,
                   reg03,
                   reg04,
                   reg05,
                   reg06,
                   reg07);
  input phi;
  input AluDivFinish;
  input [127:0] AluDivQ;
  input [127:0] AluDivR;
  input FpuBasicFinish;
  input [127:0] FpuBasicRes;
  input FpuMultFinish;
  input [127:0] FpuMultRes;
  output [127:0] AluDivA;
  output [127:0] AluDivB;
  output AluDivStall;
  output AluDivValid;
  output [127:0] FpuBasicA;
  output [127:0] FpuBasicB;
  output [5:0] FpuBasicOp;
  output FpuBasicStall;
  output FpuBasicValid;
  output [127:0] FpuMultA;
  output [127:0] FpuMultB;
  output [5:0] FpuMultOp;
  output FpuMultStall;
  output FpuMultValid;
  output char_out;
  output [6:0] char_out_val;
  output [31:0] reg00;
  output [31:0] reg01;
  output [31:0] reg02;
  output [31:0] reg03;
  output [31:0] reg04;
  output [31:0] reg05;
  output [31:0] reg06;
  output [31:0] reg07;

  reg [31:0] ram_array0[255:0];
  reg [31:0] ram_array1[255:0];
  reg [31:0] ram_array2[255:0];
  reg [31:0] ram_array3[255:0];
  reg x58, x59, x60, x61, x62, x63, x602, x603;
  reg x604, x605, x606, x607, x608, x609, x610, x611;
  reg x612, x613, x614, x615, x616, x617, x618, x619;
  reg x620, x621, x622, x623, x624, x625, x626, x627;
  reg x628, x629, x630, x631, x632, x633, x674, x675;
  reg x676, x677, x1232, x1238, x1244, x1250, x1256, x1262;
  reg x1268, x1274, x1281, x1288, x1294, x1300, x1306, x1312;
  reg x1318, x1324, x1330, x1336, x1342, x1348, x1354, x1360;
  reg x1366, x1372, x1379, x1386, x1392, x1398, x1404, x1410;
  reg x1416, x1422, x1758, x1768, x1778, x1788, x1798, x1808;
  reg x1818, x1828, x1914, x1918, x1922, x1926, x1930, x1934;
  reg x1940, x1944, x1948, x1952, x1956, x1960, x1966, x1970;
  reg x1974, x1978, x1982, x1986, x1992, x1996, x2000, x2004;
  reg x2008, x2012, x2018, x2022, x2026, x2030, x2034, x2038;
  reg x2044, x2048, x2052, x2056, x2060, x2064, x2070, x2074;
  reg x2078, x2082, x2086, x2090, x2096, x2100, x2104, x2108;
  reg x2112, x2116, x2317, x2321, x2325, x2329, x2333, x2337;
  reg x2341, x2345, x2349, x2353, x2357, x2361, x2365, x2369;
  reg x2373, x2377, x2381, x2385, x2389, x2393, x2397, x2401;
  reg x2405, x2409, x2413, x2417, x2421, x2425, x2429, x2433;
  reg x2437, x2441, x2447, x2451, x2455, x2459, x2463, x2467;
  reg x2471, x2475, x2479, x2483, x2487, x2491, x2495, x2499;
  reg x2503, x2507, x2511, x2515, x2519, x2523, x2527, x2531;
  reg x2535, x2539, x2543, x2547, x2551, x2555, x2559, x2563;
  reg x2567, x2571, x2577, x2581, x2585, x2589, x2593, x2597;
  reg x2601, x2605, x2609, x2613, x2617, x2621, x2625, x2629;
  reg x2633, x2637, x2641, x2645, x2649, x2653, x2657, x2661;
  reg x2665, x2669, x2673, x2677, x2681, x2685, x2689, x2693;
  reg x2697, x2701, x2707, x2711, x2715, x2719, x2723, x2727;
  reg x2731, x2735, x2739, x2743, x2747, x2751, x2755, x2759;
  reg x2763, x2767, x2771, x2775, x2779, x2783, x2787, x2791;
  reg x2795, x2799, x2803, x2807, x2811, x2815, x2819, x2823;
  reg x2827, x2831, x2837, x2841, x2845, x2849, x2853, x2857;
  reg x2861, x2865, x2869, x2873, x2877, x2881, x2885, x2889;
  reg x2893, x2897, x2901, x2905, x2909, x2913, x2917, x2921;
  reg x2925, x2929, x2933, x2937, x2941, x2945, x2949, x2953;
  reg x2957, x2961, x2967, x2971, x2975, x2979, x2983, x2987;
  reg x2991, x2995, x2999, x3003, x3007, x3011, x3015, x3019;
  reg x3023, x3027, x3031, x3035, x3039, x3043, x3047, x3051;
  reg x3055, x3059, x3063, x3067, x3071, x3075, x3079, x3083;
  reg x3087, x3091, x3097, x3101, x3105, x3109, x3113, x3117;
  reg x3121, x3125, x3129, x3133, x3137, x3141, x3145, x3149;
  reg x3153, x3157, x3161, x3165, x3169, x3173, x3177, x3181;
  reg x3185, x3189, x3193, x3197, x3201, x3205, x3209, x3213;
  reg x3217, x3221, x3227, x3231, x3235, x3239, x3243, x3247;
  reg x3251, x3255, x3259, x3263, x3267, x3271, x3275, x3279;
  reg x3283, x3287, x3291, x3295, x3299, x3303, x3307, x3311;
  reg x3315, x3319, x3323, x3327, x3331, x3335, x3339, x3343;
  reg x3347, x3351, x3358, x3363, x3367, x3371, x3375, x3379;
  reg x3383, x3387, x3391, x3395, x3399, x3403, x3407, x3411;
  reg x3415, x3419, x3423, x3427, x3431, x3435, x3439, x3443;
  reg x3447, x3451, x3455, x3459, x3463, x3467, x3471, x3475;
  reg x3479, x3483, x3489, x3493, x3497, x3501, x3505, x3509;
  reg x3513, x3517, x3521, x3525, x3529, x3533, x3537, x3541;
  reg x3545, x3549, x3553, x3557, x3561, x3565, x3569, x3573;
  reg x3577, x3581, x3585, x3589, x3593, x3597, x3601, x3605;
  reg x3609, x3613, x3619, x3623, x3627, x3631, x3635, x3639;
  reg x3643, x3647, x3651, x3655, x3659, x3663, x3667, x3671;
  reg x3675, x3679, x3683, x3687, x3691, x3695, x3699, x3703;
  reg x3707, x3711, x3715, x3719, x3723, x3727, x3731, x3735;
  reg x3739, x3743, x3749, x3753, x3757, x3761, x3765, x3769;
  reg x3773, x3777, x3781, x3785, x3789, x3793, x3797, x3801;
  reg x3805, x3809, x3813, x3817, x3821, x3825, x3829, x3833;
  reg x3837, x3841, x3845, x3849, x3853, x3857, x3861, x3865;
  reg x3869, x3873, x3879, x3883, x3887, x3891, x3895, x3899;
  reg x3903, x3907, x3911, x3915, x3919, x3923, x3927, x3931;
  reg x3935, x3939, x3943, x3947, x3951, x3955, x3959, x3963;
  reg x3967, x3971, x3975, x3979, x3983, x3987, x3991, x3995;
  reg x3999, x4003, x4009, x4013, x4017, x4021, x4025, x4029;
  reg x4033, x4037, x4041, x4045, x4049, x4053, x4057, x4061;
  reg x4065, x4069, x4073, x4077, x4081, x4085, x4089, x4093;
  reg x4097, x4101, x4105, x4109, x4113, x4117, x4121, x4125;
  reg x4129, x4133, x4139, x4143, x4147, x4151, x4155, x4159;
  reg x4163, x4167, x4171, x4175, x4179, x4183, x4187, x4191;
  reg x4195, x4199, x4203, x4207, x4211, x4215, x4219, x4223;
  reg x4227, x4231, x4235, x4239, x4243, x4247, x4251, x4255;
  reg x4259, x4263, x4269, x4273, x4277, x4281, x4285, x4289;
  reg x4293, x4297, x4301, x4305, x4309, x4313, x4317, x4321;
  reg x4325, x4329, x4333, x4337, x4341, x4345, x4349, x4353;
  reg x4357, x4361, x4365, x4369, x4373, x4377, x4381, x4385;
  reg x4389, x4393, x4399, x4404, x4409, x4413, x4417, x4421;
  reg x4425, x4429, x4433, x4437, x4441, x4445, x4449, x4453;
  reg x4457, x4461, x4465, x4469, x4473, x4477, x4481, x4485;
  reg x4489, x4493, x4497, x4501, x4505, x4509, x4513, x4517;
  reg x4521, x4525, x4531, x4535, x4539, x4543, x4547, x4551;
  reg x4555, x4559, x4563, x4567, x4571, x4575, x4579, x4583;
  reg x4587, x4591, x4595, x4599, x4603, x4607, x4611, x4615;
  reg x4619, x4623, x4627, x4631, x4635, x4639, x4643, x4647;
  reg x4651, x4655, x4661, x4665, x4669, x4673, x4677, x4681;
  reg x4685, x4689, x4693, x4697, x4701, x4705, x4709, x4713;
  reg x4717, x4721, x4725, x4729, x4733, x4737, x4741, x4745;
  reg x4749, x4753, x4757, x4761, x4765, x4769, x4773, x4777;
  reg x4781, x4785, x4791, x4795, x4799, x4803, x4807, x4811;
  reg x4815, x4819, x4823, x4827, x4831, x4835, x4839, x4843;
  reg x4847, x4851, x4855, x4859, x4863, x4867, x4871, x4875;
  reg x4879, x4883, x4887, x4891, x4895, x4899, x4903, x4907;
  reg x4911, x4915, x4921, x4925, x4929, x4933, x4937, x4941;
  reg x4945, x4949, x4953, x4957, x4961, x4965, x4969, x4973;
  reg x4977, x4981, x4985, x4989, x4993, x4997, x5001, x5005;
  reg x5009, x5013, x5017, x5021, x5025, x5029, x5033, x5037;
  reg x5041, x5045, x5051, x5055, x5059, x5063, x5067, x5071;
  reg x5075, x5079, x5083, x5087, x5091, x5095, x5099, x5103;
  reg x5107, x5111, x5115, x5119, x5123, x5127, x5131, x5135;
  reg x5139, x5143, x5147, x5151, x5155, x5159, x5163, x5167;
  reg x5171, x5175, x5181, x5185, x5189, x5193, x5197, x5201;
  reg x5205, x5209, x5213, x5217, x5221, x5225, x5229, x5233;
  reg x5237, x5241, x5245, x5249, x5253, x5257, x5261, x5265;
  reg x5269, x5273, x5277, x5281, x5285, x5289, x5293, x5297;
  reg x5301, x5305, x5311, x5315, x5319, x5323, x5327, x5331;
  reg x5335, x5339, x5343, x5347, x5351, x5355, x5359, x5363;
  reg x5367, x5371, x5375, x5379, x5383, x5387, x5391, x5395;
  reg x5399, x5403, x5407, x5411, x5415, x5419, x5423, x5427;
  reg x5431, x5435, x5442, x5448, x5453, x5457, x5461, x5465;
  reg x5469, x5473, x5477, x5481, x5485, x5489, x5493, x5497;
  reg x5501, x5505, x5509, x5513, x5517, x5521, x5525, x5529;
  reg x5533, x5537, x5541, x5545, x5549, x5553, x5557, x5561;
  reg x5565, x5569, x5575, x5579, x5583, x5587, x5591, x5595;
  reg x5599, x5603, x5607, x5611, x5615, x5619, x5623, x5627;
  reg x5631, x5635, x5639, x5643, x5647, x5651, x5655, x5659;
  reg x5663, x5667, x5671, x5675, x5679, x5683, x5687, x5691;
  reg x5695, x5699, x5705, x5709, x5713, x5717, x5721, x5725;
  reg x5729, x5733, x5737, x5741, x5745, x5749, x5753, x5757;
  reg x5761, x5765, x5769, x5773, x5777, x5781, x5785, x5789;
  reg x5793, x5797, x5801, x5805, x5809, x5813, x5817, x5821;
  reg x5825, x5829, x5835, x5839, x5843, x5847, x5851, x5855;
  reg x5859, x5863, x5867, x5871, x5875, x5879, x5883, x5887;
  reg x5891, x5895, x5899, x5903, x5907, x5911, x5915, x5919;
  reg x5923, x5927, x5931, x5935, x5939, x5943, x5947, x5951;
  reg x5955, x5959, x5965, x5969, x5973, x5977, x5981, x5985;
  reg x5989, x5993, x5997, x6001, x6005, x6009, x6013, x6017;
  reg x6021, x6025, x6029, x6033, x6037, x6041, x6045, x6049;
  reg x6053, x6057, x6061, x6065, x6069, x6073, x6077, x6081;
  reg x6085, x6089, x6095, x6099, x6103, x6107, x6111, x6115;
  reg x6119, x6123, x6127, x6131, x6135, x6139, x6143, x6147;
  reg x6151, x6155, x6159, x6163, x6167, x6171, x6175, x6179;
  reg x6183, x6187, x6191, x6195, x6199, x6203, x6207, x6211;
  reg x6215, x6219, x6225, x6229, x6233, x6237, x6241, x6245;
  reg x6249, x6253, x6257, x6261, x6265, x6269, x6273, x6277;
  reg x6281, x6285, x6289, x6293, x6297, x6301, x6305, x6309;
  reg x6313, x6317, x6321, x6325, x6329, x6333, x6337, x6341;
  reg x6345, x6349, x6355, x6359, x6363, x6367, x6371, x6375;
  reg x6379, x6383, x6387, x6391, x6395, x6399, x6403, x6407;
  reg x6411, x6415, x6419, x6423, x6427, x6431, x6435, x6439;
  reg x6443, x6447, x6451, x6455, x6459, x6463, x6467, x6471;
  reg x6475, x6479, x14598, x14608, x14618, x14628, x14638, x14648;
  reg x14658, x14668, x14767, x14771, x14775, x14779, x14783, x14787;
  reg x14793, x14797, x14801, x14805, x14809, x14813, x14819, x14823;
  reg x14827, x14831, x14835, x14839, x14845, x14849, x14853, x14857;
  reg x14861, x14865, x14871, x14875, x14879, x14883, x14887, x14891;
  reg x14897, x14901, x14905, x14909, x14913, x14917, x14923, x14927;
  reg x14931, x14935, x14939, x14943, x14949, x14953, x14957, x14961;
  reg x14965, x14969, x27755, x27759, x27763, x27767, x27771, x27775;
  reg x27779, x27783, x27787, x27791, x27795, x27799, x27803, x27807;
  reg x27811, x27815, x27819, x27823, x27827, x27831, x27835, x27839;
  reg x27843, x27847, x27851, x27855, x27859, x27863, x27867, x27871;
  reg x27875, x27879, x38722, x38726, x38730, x38734, x38738, x38742;
  reg x38746, x38750, x38754, x38758, x38762, x38766, x38770, x38774;
  reg x38778, x38782, x38786, x38790, x38794, x38798, x38802, x38806;
  reg x38810, x38814, x38818, x38822, x38826, x38830, x38834, x38838;
  reg x38842, x38846, x49689, x49693, x49697, x49701, x49705, x49709;
  reg x49713, x49717, x49721, x49725, x49729, x49733, x49737, x49741;
  reg x49745, x49749, x49753, x49757, x49761, x49765, x49769, x49773;
  reg x49777, x49781, x49785, x49789, x49793, x49797, x49801, x49805;
  reg x49809, x49813, x60656, x60660, x60664, x60668, x60672, x60676;
  reg x60680, x60684, x60688, x60692, x60696, x60700, x60704, x60708;
  reg x60712, x60716, x60720, x60724, x60728, x60732, x60736, x60740;
  reg x60744, x60748, x60752, x60756, x60760, x60764, x60768, x60772;
  reg x60776, x60780, x60784, x60788, x60792, x60796, x60800, x60804;
  reg x60808, x60812, x60816, x60820, x60824, x60828, x60832, x60836;
  reg x60840, x60976, x61105, x61234, x61363, x61367, x61371, x61375;
  reg x61379, x61383, x61387, x61391, x61395, x61399, x61403, x61407;
  reg x61411, x61415, x61419, x61423, x61981, x61988, x61995, x62002;
  reg x62009, x62016, x62023, x62030, x62037, x62044, x62051, x62058;
  reg x62065, x62072, x62079, x62086, x62093, x62100, x62107, x62114;
  reg x62121, x62128, x62135, x62142, x62149, x62156, x62163, x62170;
  reg x62177, x62184, x62191, x62198, x62205, x62212, x62219, x62226;
  reg x62233, x62240, x62247, x62254, x62261, x62268, x62275, x62282;
  reg x62289, x62296, x62303, x62310, x62317, x62324, x62331, x62338;
  reg x62345, x62352, x62359, x62366, x62373, x62380, x62387, x62394;
  reg x62401, x62408, x62415, x62422, x62429, x62436, x62443, x62450;
  reg x62457, x62464, x62471, x62478, x62485, x62492, x62499, x62506;
  reg x62513, x62520, x62527, x62534, x62541, x62548, x62555, x62562;
  reg x62569, x62576, x62583, x62590, x62597, x62604, x62611, x62618;
  reg x62625, x62632, x62639, x62646, x62653, x62660, x62667, x62674;
  reg x62681, x62688, x62695, x62702, x62709, x62716, x62723, x62730;
  reg x62737, x62744, x62751, x62758, x62765, x62772, x62779, x62786;
  reg x62793, x62800, x62807, x62814, x62821, x62828, x62835, x62842;
  reg x62849, x62856, x62863, x62870, x62873, x62877, x62881, x62885;
  reg x62889, x62893, x62897, x62901, x62905, x62909, x62913, x62917;
  reg x62921, x62925, x62929, x63908, x63909, x63910, x63911, x63912;
  reg x64640, x64641, x64642, x64643, x64644, x65310, x65311, x65312;
  reg x65313, x65314, x65980, x65981, x65982, x65983, x65984, x66413;
  reg x66417, x66421, x66425, x66429, x66433, x66437, x66441, x66445;
  reg x66449, x66453, x66457, x66461, x66465, x66469, x66894, x66898;
  reg x66902, x66906, x66910, x66914, x66918, x66922, x66926, x66930;
  reg x66934, x66938, x66942, x66946, x66950, x66954, x66958, x66962;
  reg x66966, x66970, x66974, x66978, x66982, x66986, x66990, x66994;
  reg x66998, x67002, x67006, x67010, x67014, x67018, x67022, x67026;
  reg x67030, x67034, x67038, x67042, x67046, x67050, x67054, x67058;
  reg x67062, x67066, x67070, x67074, x67078, x67082, x67086, x67090;
  reg x67094, x67098, x67102, x67106, x67110, x67114, x67118, x67122;
  reg x67126, x67130, x67134, x67138, x67142, x67146, x67150, x67154;
  reg x67158, x67162, x67166, x67170, x67174, x67178, x67182, x67186;
  reg x67190, x67194, x67198, x67202, x67206, x67210, x67214, x67218;
  reg x67222, x67226, x67230, x67234, x67238, x67242, x67246, x67250;
  reg x67254, x67258, x67262, x67266, x67270, x67274, x67278, x67282;
  reg x67286, x67290, x67294, x67298, x67302, x67306, x67310, x67314;
  reg x67318, x67322, x67326, x67330, x67334, x67338, x67342, x67346;
  reg x67350, x67354, x67358, x67362, x67366, x67370, x67374, x67378;
  reg x67382, x67386, x67390, x67394, x67398, x67402, x67405, x67409;
  reg x67413, x67417, x67421, x67425, x67429, x67433, x67437, x67441;
  reg x67445, x67449, x67453, x67457, x67461, x67887, x67891, x67895;
  reg x67899, x67903, x67907, x67911, x67915, x67919, x67923, x67927;
  reg x67931, x67935, x67939, x67943, x67947, x67951, x67955, x67959;
  reg x67963, x67967, x67971, x67975, x67979, x67983, x67987, x67991;
  reg x67995, x67999, x68003, x68007, x68011, x68015, x68019, x68023;
  reg x68027, x68031, x68035, x68039, x68043, x68047, x68051, x68055;
  reg x68059, x68063, x68067, x68071, x68075, x68079, x68083, x68087;
  reg x68091, x68095, x68099, x68103, x68107, x68111, x68115, x68119;
  reg x68123, x68127, x68131, x68135, x68139, x68143, x68147, x68151;
  reg x68155, x68159, x68163, x68167, x68171, x68175, x68179, x68183;
  reg x68187, x68191, x68195, x68199, x68203, x68207, x68211, x68215;
  reg x68219, x68223, x68227, x68231, x68235, x68239, x68243, x68247;
  reg x68251, x68255, x68259, x68263, x68267, x68271, x68275, x68279;
  reg x68283, x68287, x68291, x68295, x68299, x68303, x68307, x68311;
  reg x68315, x68319, x68323, x68327, x68331, x68335, x68339, x68343;
  reg x68347, x68351, x68355, x68359, x68363, x68367, x68371, x68375;
  reg x68379, x68383, x68387, x68391, x68395, x68398, x68402, x68406;
  reg x68410, x68414, x68418, x68422, x68426, x68430, x68434, x68438;
  reg x68442, x68446, x68450, x68454, x68618, x68619, x68620, x68621;
  reg x68622, x68623, x71147, x71152, x71157, x71162, x71167, x71172;
  reg x71177, x71182, x71185, x71188, x71191, x71194, x71197, x71202;
  reg x71205, x71210, x71215, x71220, x71225, x71230, x71235, x71240;
  reg x71245, x71250, x71255, x71260, x71265, x71270, x71275, x71277;
  reg x71279, x71284, x71289, x71294, x71299, x71304, x71309, x71314;
  reg x71319, x71324, x71329, x71334, x71339, x71344, x71349, x71354;
  reg x71359, x71364, x71369, x71374, x71379, x71384, x71389, x71394;
  reg x71399, x71404, x71409, x71414, x71419, x71424, x71429, x71434;
  reg x71439, x71444, x71449, x71454, x71459, x71464, x71469, x71474;
  reg x71479, x71482, x71485, x71490, x71495, x71500, x71505, x71510;
  reg x71515, x71520, x71525, x71530, x71535, x71540, x71545, x71550;
  reg x71555, x71560, x71565, x71570, x71575, x71580, x71585, x71590;
  reg x71595, x71600, x71605, x71610, x71615, x71620, x71625, x71630;
  reg x71635, x71642, x71647, x71652, x71657, x71662, x71667, x71672;
  reg x71677, x71682, x71687, x71692, x71697, x71702, x71707, x71712;
  reg x71717, x71722, x71727, x71732, x71737, x71742, x71747, x71752;
  reg x71757, x71762, x71767, x71772, x71777, x71782, x71787, x71792;
  reg x71797, x71802, x71807, x71812, x71817, x71822, x71827, x71832;
  reg x71837, x71842, x71847, x71852, x71857, x71862, x71867, x71872;
  reg x71877, x71882, x71887, x71892, x71897, x71902, x71907, x71910;
  reg x71913, x71916, x71919, x71922, x71925, x71928, x71931, x71934;
  reg x71937, x71942, x71947, x71952, x71957, x71962, x71967, x71972;
  reg x71977, x71982, x71987, x71992, x71997, x72002, x72007, x72012;
  reg x72017, x72022, x72027, x72032, x72037, x72042, x72047, x72052;
  reg x72057, x72062, x72067, x72072, x72077, x72082, x72087, x72092;
  reg x72097, x72102, x72107, x72112, x72117, x72122, x72127, x72132;
  reg x72137, x72142, x72147, x72152, x72157, x72162, x72167, x72172;
  reg x72177, x72182, x72187, x72192, x72197, x72202, x72207, x72212;
  reg x72217, x72222, x72227, x72232, x72237, x72242, x72247, x72252;
  reg x72257, x72262, x72267, x72272, x72277, x72282, x72287, x72292;
  reg x72297, x72302, x72307, x72312, x72317, x72322, x72327, x72332;
  reg x72337, x72342, x72347, x72352, x72357, x72362, x72367, x72372;
  reg x72377, x72382, x72387, x72392, x72397, x72402, x72407, x72412;
  reg x72417, x72422, x72427, x72432, x72437, x72442, x72447, x72452;
  reg x72457, x72462, x72467, x72472, x72477, x72482, x72487, x72492;
  reg x72497, x72502, x72507, x72512, x72517, x72522, x72527, x72532;
  reg x72537, x72542, x72547, x72552, x72557, x72562, x72567, x72572;
  reg x72577, x72582, x72587, x72592, x72597, x72602, x72607, x72612;
  reg x72617, x72622, x72627, x72632, x72637, x72642, x72647, x72652;
  reg x72657, x72662, x72667, x72672, x72677, x72682, x72687, x72692;
  reg x72697, x72702, x72707, x72712, x72717, x72722, x72727, x72732;
  reg x72737, x72742, x72747, x72752, x72757, x72762, x72767, x72772;
  reg x72777, x72782, x72787, x72792, x72797, x72802, x72807, x72812;
  reg x72817, x72822, x72827, x72832, x72837, x72842, x72847, x72852;
  reg x72857, x72862, x72867, x72872, x72877, x72882, x72887, x72892;
  reg x72897, x72902, x72907, x72912, x72917, x72922, x72927, x72932;
  reg x72937, x72942, x72947, x72952, x72957, x72962, x72967, x72972;
  reg x72977, x72982, x72987, x72992, x72997, x73002, x73007, x73012;
  reg x73017, x73022, x73027, x73032, x73037, x73042, x73047, x73052;
  reg x73057, x73062, x73067, x73072, x73077, x73082, x73087, x73092;
  reg x73097, x73102, x73107, x73112, x73117, x73122, x73127, x73132;
  reg x73137, x73142, x73147, x73152, x73157, x73162, x73167, x73172;
  reg x73177, x73182, x73187, x73192, x73197, x73202, x73207, x73212;
  reg x73217, x73222, x73227, x73232, x73237, x73242, x73247, x73252;
  reg x73257, x73262, x73267, x73272, x73277, x73282, x73287, x73292;
  reg x73297, x73302, x73307, x73312, x73317, x73322, x73327, x73332;
  reg x73337, x73342, x73347, x73352, x73357, x73362, x73367, x73372;
  reg x73377, x73382, x73387, x73392, x73397, x73402, x73407, x73412;
  reg x73417, x73422, x73427, x73432, x73437, x73442, x73447, x73452;
  reg x73457, x73462, x73467, x73472, x73477, x73482, x73487, x73492;
  reg x73497, x73502, x73507, x73512, x73517, x73522, x73527, x73532;
  reg x73537, x73542, x73547, x73552, x73557, x73562, x73567, x73572;
  reg x73577, x73582, x73587, x73592, x73597, x73602, x73607, x73612;
  reg x73617, x73622, x73627, x73632, x73637, x73642, x73647, x73652;
  reg x73657, x73662, x73667, x73672, x73677, x73682, x73687, x73692;
  reg x73697, x73702, x73707, x73712, x73717, x73722, x73727, x73732;
  reg x73737, x73742, x73747, x73752, x73757, x73762, x73767, x73772;
  reg x73777, x73782, x73787, x73792, x73797, x73802, x73807, x73812;
  reg x73817, x73822, x73827, x73832, x73837, x73842, x73847, x73852;
  reg x73857, x73862, x73867, x73872, x73877, x73882, x73887, x73892;
  reg x73897, x73902, x73907, x73912, x73917, x73922, x73927, x73932;
  reg x73937, x73942, x73947, x73952, x73957, x73962, x73967, x73972;
  reg x73977, x73982, x73987, x73992, x73997, x74002, x74005, x74008;
  reg x74011, x74014, x74017, x74020, x74023, x74026, x74029, x74032;
  reg x74035, x74038, x74041, x74044, x74047, x74050, x74053, x74056;
  reg x74059, x74062, x74065, x74068, x74071, x74074, x74077, x74080;
  reg x74083, x74086, x74089, x74092, x74095, x74098, x74101, x74104;
  reg x74107, x74110, x74113, x74116, x74119, x74122, x74125, x74128;
  reg x74131, x74134, x74137, x74140, x74143, x74146, x74149, x74152;
  reg x74155, x74158, x74161, x74164, x74167, x74170, x74173, x74176;
  reg x74179, x74182, x74185, x74188, x74191, x74194, x74197, x74200;
  reg x74203, x74206, x74209, x74212, x74215, x74218, x74221, x74224;
  reg x74227, x74230, x74233, x74236, x74239, x74242, x74245, x74248;
  reg x74251, x74254, x74257, x74260, x74263, x74266, x74269, x74272;
  reg x74275, x74278, x74281, x74284, x74287, x74290, x74293, x74296;
  reg x74299, x74302, x74305, x74308, x74311, x74314, x74317, x74320;
  reg x74323, x74326, x74329, x74332, x74335, x74338, x74341, x74344;
  reg x74347, x74350, x74353, x74356, x74359, x74362, x74365, x74368;
  reg x74371, x74374, x74377, x74380, x74383, x74386, x74389, x74392;
  reg x74395, x74398, x74401, x74404, x74407, x74410, x74413, x74416;
  reg x74419, x74422, x74425, x74428, x74431, x74434, x74437, x74440;
  reg x74443, x74446, x74449, x74452, x74455, x74458, x74461, x74464;
  reg x74467, x74470, x74473, x74476, x74479, x74482, x74485, x74488;
  reg x74491, x74494, x74497, x74500, x74503, x74506, x74509, x74512;
  reg x74515, x74518, x74521, x74524, x74527, x74530, x74533, x74536;
  reg x74539, x74542, x74545, x74548, x74551, x74554, x74557, x74560;
  reg x74563, x74566, x74569, x74572, x74575, x74578, x74581, x74584;
  reg x74587, x74590, x74593, x74596, x74599, x74602, x74605, x74608;
  reg x74611, x74614, x74617, x74620, x74623, x74626, x74629, x74632;
  reg x74635, x74638, x74641, x74644, x74647, x74650, x74653, x74656;
  reg x74659, x74662, x74665, x74668, x74671, x74674, x74677, x74680;
  reg x74683, x74686, x74689, x74692, x74695, x74698, x74701, x74704;
  reg x74707, x74710, x74713, x74716, x74719, x74722, x74725, x74728;
  reg x74731, x74734, x74737, x74740, x74743, x74746, x74749, x74752;
  reg x74755, x74758, x74761, x74764, x74767, x74770, x74773, x74776;
  reg x74779, x74782, x74785, x74788, x74791, x74794, x74797, x74800;
  reg x74803, x74806, x74809, x74812, x74815, x74818, x74821, x74824;
  reg x74827, x74830, x74833, x74836, x74839, x74842, x74845, x74848;
  reg x74851, x74854, x74857, x74860, x74863, x74866, x74869, x74872;
  reg x74875, x74878, x74881, x74884, x74887, x74890, x74893, x74896;
  reg x74899, x74902, x74905, x74908, x74911, x74914, x74917, x74920;
  reg x74923, x74926, x74929, x74932, x74935, x74938, x74941, x74944;
  reg x74947, x74950, x74953, x74956, x74959, x74962, x74965, x74968;
  reg x74971, x74974, x74977, x74980, x74983, x74986, x74989, x74992;
  reg x74995, x74998, x75001, x75004, x75007, x75010, x75013, x75016;
  reg x75019, x75022, x75025, x75028, x75031, x75034, x75037, x75040;
  reg x75043, x75046, x75049, x75052, x75055, x75058, x75061, x75064;
  reg x75067, x75070, x75073, x75076, x75079, x75082, x75085, x75088;
  reg x75091, x75094, x75097, x75100, x75103, x75106, x75109, x75112;
  reg x75115, x75118, x75121, x75124, x75127, x75130, x75133, x75136;
  reg x75139, x75142, x75145, x75148, x75151, x75154, x75157, x75160;
  reg x75163, x75166, x75169, x75172, x75175, x75178, x75181, x75184;
  reg x75187, x75190, x75193, x75196, x75199, x75202, x75205, x75208;
  reg x75211, x75214, x75217, x75220, x75223, x75226, x75229, x75232;
  reg x75235, x75238, x75241, x75244, x75247, x75250, x75253, x75256;
  reg x75259, x75262, x75265, x75268, x75271, x75274, x75277, x75280;
  reg x75283, x75286, x75289, x75292, x75295, x75298, x75301, x75304;
  reg x75307, x75310, x75313, x75316, x75319, x75322, x75325, x75328;
  reg x75331, x75334, x75337, x75340, x75343, x75346, x75349, x75352;
  reg x75355, x75358, x75361, x75364, x75367, x75370, x75373, x75376;
  reg x75379, x75382, x75385, x75388, x75391, x75394, x75397, x75400;
  reg x75403, x75406, x75409, x75412, x75415, x75418, x75421, x75424;
  reg x75427, x75430, x75433, x75436, x75439, x75442, x75445, x75448;
  reg x75451, x75454, x75457, x75460, x75463, x75466, x75469, x75472;
  reg x75475, x75478, x75481, x75484, x75487, x75490, x75493, x75496;
  reg x75499, x75502, x75505, x75508, x75511, x75514, x75517, x75520;
  reg x75523, x75526, x75529, x75532, x75535, x75538, x75541, x75544;
  reg x75547, x75550, x75553, x75556, x75559, x75562, x75565, x75568;
  reg x75571, x75574, x75577, x75580, x75583, x75586, x75589, x75592;
  reg x75595, x75598, x75601, x75604, x75607, x75610, x75613, x75616;
  reg x75619, x75622, x75625, x75628, x75631, x75634, x75637, x75640;
  reg x75643, x75646, x75649, x75652, x75655, x75658, x75661, x75664;
  reg x75667, x75670, x75673, x75676, x75679, x75682, x75685, x75688;
  reg x75691, x75694, x75697, x75700, x75703, x75706, x75709, x75712;
  reg x75715, x75718, x75721, x75724, x75727, x75730, x75733, x75736;
  reg x75739, x75742, x75745, x75748, x75751, x75754, x75757, x75760;
  reg x75763, x75766, x75769, x75772, x75775, x75778, x75781, x75784;
  reg x75787, x75790, x75793, x75796, x75799, x75802, x75805, x75808;
  reg x75811, x75814, x75817, x75820, x75823, x75826, x75829, x75832;
  reg x75835, x75838, x75841, x75844, x75847, x75850, x75853, x75856;
  reg x75859, x75862, x75865, x75868, x75871, x75874, x75877, x75880;
  reg x75883, x75886, x75889, x75892, x75895, x75898, x75901, x75904;
  reg x75907, x75910, x75913, x75916, x75919, x75922, x75925, x75928;
  reg x75931, x75934, x75937, x75940, x75943, x75946, x75949, x75952;
  reg x75955, x75958, x75961, x75964, x75967, x75970, x75973, x75976;
  reg x75979, x75982, x75985, x75988, x75991, x75994, x75997, x76000;
  reg x76003, x76006, x76009, x76012, x76015, x76018, x76021, x76024;
  reg x76027, x76030, x76033, x76036, x76039, x76042, x76045, x76048;
  reg x76051, x76054, x76057, x76060, x76063, x76066, x76069, x76072;
  reg x76075, x76078, x76081, x76084, x76087, x76090, x76093, x76096;
  reg x76099, x76102, x76105, x76108, x76111, x76114, x76117, x76120;
  reg x76123, x76126, x76129, x76132, x76135, x76138, x76141, x76144;
  reg x76147, x76150, x76153, x76156, x76159, x76162, x76165, x76168;
  reg x76171, x76174, x76177, x76180, x76183, x76186, x76189, x76192;
  reg x76195, x76198, x76201, x76204, x76207, x76210, x76213, x76216;
  reg x76219, x76222, x76225, x76228, x76231, x76234, x76237, x76240;
  reg x76243, x76246, x76249, x76252, x76255, x76258, x76261, x76264;
  reg x76267, x76270, x76273, x76276, x76279, x76282, x76285, x76288;
  reg x76291, x76294, x76297, x76300, x76303, x76306, x76309, x76312;
  reg x76315, x76318, x76321, x76324, x76327, x76330, x76333, x76336;
  reg x76339, x76342, x76345, x76348, x76351, x76354, x76357, x76360;
  reg x76363, x76366, x76369, x76372, x76375, x76378, x76381, x76384;
  reg x76387, x76390, x76393, x76396, x76399, x76402, x76405, x76408;
  reg x76411, x76414, x76417, x76420, x76423, x76426, x76429, x76432;
  reg x76435, x76438, x76441, x76444, x76447, x76450, x76453, x76456;
  reg x76459, x76462, x76465, x76468, x76471, x76474, x76477, x76480;
  reg x76483, x76486, x76489, x76492, x76495, x76498, x76501, x76504;
  reg x76507, x76510, x76513, x76516, x76519, x76522, x76525, x76528;
  reg x76531, x76534, x76537, x76540, x76543, x76546, x76549, x76552;
  reg x76555, x76558, x76561, x76564, x76567, x76570, x76573, x76576;
  reg x76579, x76582, x76585, x76588, x76591, x76594, x76597, x76600;
  reg x76603, x76606, x76609, x76612, x76615, x76618, x76621, x76624;
  reg x76627, x76630, x76633, x76636, x76639, x76642, x76645, x76648;
  reg x76651, x76654, x76657, x76660, x76663, x76666, x76669, x76672;
  reg x76675, x76678, x76681, x76684, x76687, x76690, x76693, x76696;
  reg x76699, x76702, x76705, x76708, x76711, x76714, x76717, x76720;
  reg x76723, x76726, x76729, x76732, x76735, x76738, x76741, x76744;
  reg x76747, x76750, x76753, x76756, x76759, x76762, x76765, x76768;
  reg x76771, x76774, x76777, x76780, x76783, x76786, x76789, x76792;
  reg x76795, x76798, x76801, x76804, x76807, x76810, x76813, x76816;
  reg x76819, x76822, x76825, x76828, x76831, x76834, x76837, x76840;
  reg x76843, x76846, x76849, x76852, x76855, x76858, x76861, x76864;
  reg x76867, x76870, x76873, x76876, x76879, x76882, x76885, x76888;
  reg x76891, x76894, x76897, x76900, x76903, x76906, x76909, x76912;
  reg x76915, x76918, x76921, x76924, x76927, x76930, x76933, x76936;
  reg x76939, x76942, x76945, x76948, x76951, x76954, x76957, x76960;
  reg x76963, x76966, x76969, x76972, x76975, x76978, x76981, x76984;
  reg x76987, x76990, x76993, x76996, x76999, x77002, x77005, x77008;
  reg x77011, x77014, x77017, x77020, x77023, x77026, x77029, x77032;
  reg x77035, x77038, x77041, x77044, x77047, x77050, x77053, x77056;
  reg x77059, x77062, x77065, x77068, x77071, x77074, x77077, x77080;
  reg x77083, x77086, x77089, x77092, x77095, x77098, x77101, x77104;
  reg x77107, x77110, x77113, x77116, x77119, x77122, x77125, x77128;
  reg x77131, x77134, x77137, x77140, x77143, x77146, x77149, x77152;
  reg x77155, x77158, x77161, x77164, x77167, x77170, x77173, x77176;
  reg x77179, x77182, x77185, x77188, x77191, x77194, x77197, x77200;
  reg x77203, x77206, x77209, x77212, x77215, x77218, x77221, x77224;
  reg x77227, x77230, x77233, x77236, x77239, x77242, x77245, x77248;
  reg x77251, x77254, x77257, x77260, x77263, x77266, x77269, x77272;
  reg x77275, x77278, x77281, x77284, x77287, x77290, x77293, x77296;
  reg x77299, x77302, x77305, x77308, x77311, x77314, x77317, x77320;
  reg x77323, x77326, x77329, x77332, x77335, x77338, x77341, x77344;
  reg x77347, x77350, x77353, x77356, x77359, x77362, x77365, x77368;
  reg x77371, x77374, x77377, x77380, x77383, x77386, x77389, x77392;
  reg x77395, x77398, x77401, x77404, x77407, x77410, x77413, x77416;
  reg x77419, x77422, x77425, x77428, x77431, x77434, x77437, x77440;
  reg x77443, x77446, x77449, x77452, x77455, x77458, x77461, x77464;
  reg x77467, x77470, x77473, x77476, x77479, x77482, x77485, x77488;
  reg x77491, x77494, x77497, x77500, x77503, x77506, x77509, x77512;
  reg x77515, x77518, x77521, x77524, x77527, x77530, x77533, x77536;
  reg x77539, x77542, x77545, x77548, x77551, x77554, x77557, x77560;
  reg x77563, x77566, x77569, x77572, x77575, x77578, x77581, x77584;
  reg x77587, x77590, x77593, x77596, x77599, x77602, x77605, x77608;
  reg x77611, x77614, x77617, x77620, x77623, x77626, x77629, x77632;
  reg x77635, x77638, x77641, x77644, x77647, x77650, x77653, x77656;
  reg x77659, x77662, x77665, x77668, x77671, x77674, x77677, x77680;
  reg x77683, x77686, x77689, x77692, x77695, x77698, x77701, x77704;
  reg x77707, x77710, x77713, x77716, x77719, x77722, x77725, x77728;
  reg x77731, x77734, x77737, x77740, x77743, x77746, x77749, x77752;
  reg x77755, x77758, x77761, x77764, x77767, x77770, x77773, x77776;
  reg x77779, x77782, x77785, x77788, x77791, x77794, x77797, x77800;
  reg x77803, x77806, x77809, x77812, x77815, x77818, x77821, x77824;
  reg x77827, x77830, x77833, x77836, x77839, x77842, x77845, x77848;
  reg x77851, x77854, x77857, x77860, x77863, x77866, x77869, x77872;
  reg x77875, x77878, x77881, x77884, x77887, x77890, x77893, x77896;
  reg x77899, x77902, x77905, x77908, x77911, x77914, x77917, x77920;
  reg x77923, x77926, x77929, x77932, x77935, x77938, x77941, x77944;
  reg x77947, x77950, x77953, x77956, x77959, x77962, x77965, x77968;
  reg x77971, x77974, x77977, x77980, x77983, x77986, x77989, x77992;
  reg x77995, x77998, x78001, x78004, x78007, x78010, x78013, x78016;
  reg x78019, x78022, x78025, x78028, x78031, x78034, x78037, x78040;
  reg x78043, x78046, x78049, x78052, x78055, x78058, x78061, x78064;
  reg x78067, x78070, x78073, x78076, x78079, x78082, x78085, x78088;
  reg x78091, x78094, x78097, x78100, x78103, x78106, x78109, x78112;
  reg x78115, x78118, x78121, x78124, x78127, x78130, x78133, x78136;
  reg x78139, x78142, x78145, x78148, x78151, x78154, x78157, x78160;
  reg x78163, x78166, x78169, x78172, x78175, x78178, x78181, x78184;
  reg x78187, x78190, x78193, x78196, x78199, x78202, x78205, x78208;
  reg x78211, x78214, x78217, x78220, x78223, x78226, x78229, x78232;
  reg x78235, x78238, x78241, x78244, x78247, x78250, x78253, x78256;
  reg x78259, x78262, x78265, x78268, x78271, x78274, x78277, x78280;
  reg x78283, x78286, x78289, x78292, x78295, x78298, x78301, x78304;
  reg x78307, x78310, x78313, x78316, x78319, x78322, x78325, x78328;
  reg x78331, x78334, x78337, x78340, x78343, x78346, x78349, x78352;
  reg x78355, x78358, x78361, x78364, x78367, x78370, x78373, x78376;
  reg x78379, x78382, x78385, x78388, x78391, x78394, x78397, x78400;
  reg x78403, x78406, x78409, x78412, x78415, x78418, x78421, x78424;
  reg x78427, x78430, x78433, x78436, x78439, x78442, x78445, x78448;
  reg x78451, x78454, x78457, x78460, x78463, x78466, x78469, x78472;
  reg x78475, x78478, x78481, x78484, x78487, x78490, x78493, x78496;
  reg x78499, x78502, x78505, x78508, x78511, x78514, x78517, x78520;
  reg x78523, x78526, x78529, x78532, x78535, x78538, x78541, x78544;
  reg x78547, x78550, x78553, x78556, x78559, x78562, x78565, x78568;
  reg x78571, x78574, x78577, x78580, x78583, x78586, x78589, x78592;
  reg x78595, x78598, x78601, x78604, x78607, x78610, x78613, x78616;
  reg x78619, x78622, x78625, x78628, x78631, x78634, x78637, x78640;
  reg x78643, x78646, x78649, x78652, x78655, x78658, x78661, x78664;
  reg x78667, x78670, x78673, x78676, x78679, x78682, x78685, x78688;
  reg x78691, x78694, x78697, x78700, x78703, x78706, x78709, x78712;
  reg x78715, x78718, x78721, x78724, x78727, x78730, x78733, x78736;
  reg x78739, x78742, x78745, x78748, x78751, x78754, x78757, x78760;
  reg x78763, x78766, x78769, x78772, x78775, x78778, x78781, x78784;
  reg x78787, x78790, x78793, x78796, x78799, x78802, x78805, x78808;
  reg x78811, x78814, x78817, x78820, x78823, x78826, x78829, x78832;
  reg x78835, x78838, x78841, x78844, x78847, x78850, x78853, x78856;
  reg x78859, x78862, x78865, x78868, x78871, x78874, x78877, x78880;
  reg x78883, x78886, x78889, x78892, x78895, x78898, x78901, x78904;
  reg x78907, x78910, x78913, x78916, x78919, x78922, x78925, x78928;
  reg x78931, x78934, x78937, x78940, x78943, x78946, x78949, x78952;
  reg x78955, x78958, x78961, x78964, x78967, x78970, x78973, x78976;
  reg x78979, x78982, x78985, x78988, x78991, x78994, x78997, x79000;
  reg x79003, x79006, x79009, x79012, x79015, x79018, x79021, x79024;
  reg x79027, x79030, x79033, x79036, x79039, x79042, x79045, x79048;
  reg x79051, x79054, x79057, x79060, x79063, x79066, x79069, x79072;
  reg x79075, x79078, x79081, x79084, x79087, x79090, x79093, x79096;
  reg x79099, x79102, x79105, x79108, x79111, x79114, x79117, x79120;
  reg x79123, x79126, x79129, x79132, x79135, x79138, x79141, x79144;
  reg x79147, x79150, x79153, x79156, x79159, x79162, x79165, x79168;
  reg x79171, x79174, x79177, x79180, x79183, x79186, x79189, x79192;
  reg x79195, x79198, x79201, x79204, x79207, x79210, x79213, x79216;
  reg x79219, x79222, x79225, x79228, x79231, x79234, x79237, x79240;
  reg x79243, x79246, x79249, x79252, x79255, x79258, x79261, x79264;
  reg x79267, x79270, x79273, x79276, x79279, x79282, x79285, x79288;
  reg x79291, x79294, x79297, x79300, x79303, x79306, x79309, x79312;
  reg x79315, x79318, x79321, x79324, x79327, x79330, x79333, x79336;
  reg x79339, x79342, x79345, x79348, x79351, x79354, x79357, x79360;
  reg x79363, x79366, x79369, x79372, x79375, x79378, x79381, x79384;
  reg x79387, x79390, x79393, x79396, x79399, x79402, x79405, x79408;
  reg x79411, x79414, x79417, x79420, x79423, x79426, x79429, x79432;
  reg x79435, x79438, x79441, x79444, x79447, x79450, x79453, x79456;
  reg x79459, x79462, x79465, x79468, x79471, x79474, x79477, x79480;
  reg x79483, x79486, x79489, x79492, x79495, x79498, x79501, x79504;
  reg x79507, x79510, x79513, x79516, x79519, x79522, x79525, x79528;
  reg x79531, x79534, x79537, x79540, x79543, x79546, x79549, x79552;
  reg x79555, x79558, x79561, x79564, x79567, x79570, x79573, x79576;
  reg x79579, x79582, x79585, x79588, x79591, x79594, x79597, x79600;
  reg x79603, x79606, x79609, x79612, x79615, x79618, x79621, x79624;
  reg x79627, x79630, x79633, x79636, x79639, x79642, x79645, x79648;
  reg x79651, x79654, x79657, x79660, x79663, x79666, x79669, x79672;
  reg x79675, x79678, x79681, x79684, x79687, x79690, x79693, x79696;
  reg x79699, x79702, x79705, x79708, x79711, x79714, x79717, x79720;
  reg x79723, x79726, x79729, x79732, x79735, x79738, x79741, x79744;
  reg x79747, x79750, x79753, x79756, x79759, x79762, x79765, x79768;
  reg x79771, x79774, x79777, x79780, x79783, x79786, x79789, x79792;
  reg x79795, x79798, x79801, x79804, x79807, x79810, x79813, x79816;
  reg x79819, x79822, x79825, x79828, x79831, x79834, x79837, x79840;
  reg x79843, x79846, x79849, x79852, x79855, x79858, x79861, x79864;
  reg x79867, x79870, x79873, x79876, x79879, x79882, x79885, x79888;
  reg x79891, x79894, x79897, x79900, x79903, x79906, x79909, x79912;
  reg x79915, x79918, x79921, x79924, x79927, x79930, x79933, x79936;
  reg x79939, x79942, x79945, x79948, x79951, x79954, x79957, x79960;
  reg x79963, x79966, x79969, x79972, x79975, x79978, x79981, x79984;
  reg x79987, x79990, x79993, x79996, x79999, x80002, x80005, x80008;
  reg x80011, x80014, x80017, x80020, x80023, x80026, x80029, x80032;
  reg x80035, x80038, x80041, x80044, x80047, x80050, x80053, x80056;
  reg x80059, x80062, x80065, x80068, x80071, x80074, x80077, x80080;
  reg x80083, x80086, x80089, x80092, x80095, x80098, x80101, x80104;
  reg x80107, x80110, x80113, x80116, x80119, x80122, x80125, x80128;
  reg x80131, x80134, x80137, x80140, x80143, x80146, x80149, x80152;
  reg x80155, x80158, x80161, x80164, x80167, x80170, x80173, x80176;
  reg x80179, x80182, x80185, x80188, x80191, x80194, x80197, x80200;
  reg x80203, x80206, x80209, x80212, x80215, x80218, x80221, x80224;
  reg x80227, x80230, x80233, x80236, x80239, x80242, x80245, x80248;
  reg x80251, x80254, x80257, x80260, x80263, x80266, x80269, x80272;
  reg x80275, x80278, x80281, x80284, x80287, x80290, x80293, x80296;
  reg x80299, x80302, x80305, x80308, x80311, x80314, x80317, x80320;
  reg x80323, x80326, x80329, x80332, x80335, x80338, x80341, x80344;
  reg x80347, x80350, x80353, x80356, x80359, x80362, x80365, x80368;
  reg x80371, x80374, x80377, x80380, x80383, x80386, x80389, x80392;
  reg x80395, x80398, x80401, x80404, x80407, x80410, x80413, x80416;
  reg x80419, x80422, x80425, x80428, x80431, x80434, x80437, x80440;
  reg x80443, x80446, x80449, x80452, x80455, x80458, x80461, x80464;
  reg x80467, x80470, x80473, x80476, x80479, x80482, x80485, x80488;
  reg x80491, x80494, x80497, x80500, x80503, x80506, x80509, x80512;
  reg x80515, x80518, x80521, x80524, x80527, x80530, x80533, x80536;
  reg x80539, x80542, x80545, x80548, x80551, x80554, x80557, x80560;
  reg x80563, x80566, x80569, x80572, x80575, x80578, x80581, x80584;
  reg x80587, x80590, x80593, x80596, x80599, x80602, x80605, x80608;
  reg x80611, x80614, x80617, x80620, x80623, x80626, x80629, x80632;
  reg x80635, x80638, x80641, x80644, x80647, x80650, x80653, x80656;
  reg x80659, x80662, x80665, x80668, x80671, x80674, x80677, x80680;
  reg x80683, x80686, x80689, x80692, x80695, x80698, x80701, x80704;
  reg x80707, x80710, x80713, x80716, x80719, x80722, x80725, x80728;
  reg x80731, x80734, x80737, x80740, x80743, x80746, x80749, x80752;
  reg x80755, x80758, x80761, x80764, x80767, x80770, x80773, x80776;
  reg x80779, x80782, x80785, x80788, x80791, x80794, x80797, x80800;
  reg x80803, x80806, x80809, x80812, x80815, x80818, x80821, x80824;
  reg x80827, x80830, x80833, x80836, x80839, x80842, x80845, x80848;
  reg x80851, x80854, x80857, x80860, x80863, x80866, x80869, x80872;
  reg x80875, x80878, x80881, x80884, x80887, x80890, x80893, x80896;
  reg x80899, x80902, x80905, x80908, x80911, x80914, x80917, x80920;
  reg x80923, x80926, x80929, x80932, x80935, x80938, x80941, x80944;
  reg x80947, x80950, x80953, x80956, x80959, x80962, x80965, x80968;
  reg x80971, x80974, x80977, x80980, x80983, x80986, x80989, x80992;
  reg x80995, x80998, x81001, x81004, x81007, x81010, x81013, x81016;
  reg x81019, x81022, x81025, x81028, x81031, x81034, x81037, x81040;
  reg x81043, x81046, x81049, x81052, x81055, x81058, x81061, x81064;
  reg x81067, x81070, x81073, x81076, x81079, x81082, x81085, x81088;
  reg x81091, x81094, x81097, x81100, x81103, x81106, x81109, x81112;
  reg x81115, x81118, x81121, x81124, x81127, x81130, x81133, x81136;
  reg x81139, x81142, x81145, x81148, x81151, x81154, x81157, x81160;
  reg x81163, x81166, x81169, x81172, x81175, x81178, x81181, x81184;
  reg x81187, x81190, x81193, x81196, x81199, x81202, x81205, x81208;
  reg x81211, x81214, x81217, x81220, x81223, x81226, x81229, x81232;
  reg x81235, x81238, x81241, x81244, x81247, x81250, x81253, x81256;
  reg x81259, x81262, x81265, x81268, x81271, x81274, x81277, x81280;
  reg x81283, x81286, x81289, x81292, x81295, x81298, x81301, x81304;
  reg x81307, x81310, x81313, x81316, x81319, x81322, x81325, x81328;
  reg x81331, x81334, x81337, x81340, x81343, x81346, x81349, x81352;
  reg x81355, x81358, x81361, x81364, x81367, x81370, x81373, x81376;
  reg x81379, x81382, x81385, x81388, x81391, x81394, x81397, x81400;
  reg x81403, x81406, x81409, x81412, x81415, x81418, x81421, x81424;
  reg x81427, x81430, x81433, x81436, x81439, x81442, x81445, x81448;
  reg x81451, x81454, x81457, x81460, x81463, x81466, x81469, x81472;
  reg x81475, x81478, x81481, x81484, x81487, x81490, x81493, x81496;
  reg x81499, x81502, x81505, x81508, x81511, x81514, x81517, x81520;
  reg x81523, x81526, x81529, x81532, x81535, x81538, x81541, x81544;
  reg x81547, x81550, x81553, x81556, x81559, x81562, x81565, x81568;
  reg x81571, x81574, x81577, x81580, x81583, x81586, x81589, x81592;
  reg x81595, x81598, x81601, x81604, x81607, x81610, x81613, x81616;
  reg x81619, x81622, x81625, x81628, x81631, x81634, x81637, x81640;
  reg x81643, x81646, x81649, x81652, x81655, x81658, x81661, x81664;
  reg x81667, x81670, x81673, x81676, x81679, x81682, x81685, x81688;
  reg x81691, x81694, x81697, x81700, x81703, x81706, x81709, x81712;
  reg x81715, x81718, x81721, x81724, x81727, x81730, x81733, x81736;
  reg x81739, x81742, x81745, x81748, x81751, x81754, x81757, x81760;
  reg x81763, x81766, x81769, x81772, x81775, x81778, x81781, x81784;
  reg x81787, x81790, x81793, x81796, x81799, x81802, x81805, x81808;
  reg x81811, x81814, x81817, x81820, x81823, x81826, x81829, x81832;
  reg x81835, x81838, x81841, x81844, x81847, x81850, x81853, x81856;
  reg x81859, x81862, x81865, x81868, x81871, x81874, x81877, x81880;
  reg x81883, x81886, x81889, x81892, x81895, x81898, x81901, x81904;
  reg x81907, x81910, x81913, x81916, x81919, x81922, x81925, x81928;
  reg x81931, x81934, x81937, x81940, x81943, x81946, x81949, x81952;
  reg x81955, x81958, x81961, x81964, x81967, x81970, x81973, x81976;
  reg x81979, x81982, x81985, x81988, x81991, x81994, x81997, x82000;
  reg x82003, x82006, x82009, x82012, x82015, x82018, x82021, x82024;
  reg x82027, x82030, x82033, x82036, x82039, x82042, x82045, x82048;
  reg x82051, x82054, x82057, x82060, x82063, x82066, x82069, x82072;
  reg x82075, x82078, x82081, x82084, x82087, x82090, x82093, x82096;
  reg x82099, x82102, x82105, x82108, x82111, x82114, x82117, x82120;
  reg x82123, x82126, x82129, x82132, x82135, x82138, x82141, x82144;
  reg x82147, x82150, x82153, x82156, x82159, x82162, x82165, x82168;
  reg x82171, x82174, x82177, x82180, x82183, x82186, x82189, x82192;
  reg x82195, x82198, x82201, x82204, x82207, x82210, x82213, x82216;
  reg x82219, x82222, x82225, x82228, x82231, x82234, x82237, x82240;
  reg x82243, x82246, x82249, x82252, x82255, x82258, x82261, x82264;
  reg x82267, x82270, x82273, x82276, x82279, x82282, x82285, x82288;
  reg x82291, x82294, x82297, x82300, x82303, x82306, x82309, x82312;
  reg x82315, x82318, x82321, x82324, x82327, x82330, x82333, x82336;
  reg x82339, x82342, x82345, x82348, x82351, x82354, x82357, x82360;
  reg x82363, x82366, x82369, x82372, x82375, x82378, x82381, x82384;
  reg x82387, x82390, x82393, x82396, x82399, x82402, x82405, x82408;
  reg x82411, x82414, x82417, x82420, x82423, x82426, x82429, x82432;
  reg x82435, x82438, x82441, x82444, x82447, x82450, x82453, x82456;
  reg x82459, x82462, x82465, x82468, x82471, x82474, x82477, x82480;
  reg x82483, x82486, x82489, x82492, x82495, x82498, x82501, x82504;
  reg x82507, x82510, x82513, x82516, x82519, x82522, x82525, x82528;
  reg x82531, x82534, x82537, x82540, x82543, x82546, x82549, x82552;
  reg x82555, x82558, x82561, x82564, x82567, x82570, x82573, x82576;
  reg x82579, x82582, x82585, x82588, x82591, x82594, x82597, x82600;
  reg x82603, x82606, x82609, x82612, x82615, x82618, x82621, x82624;
  reg x82627, x82630, x82633, x82636, x82639, x82642, x82645, x82648;
  reg x82651, x82654, x82657, x82660, x82663, x82666, x82669, x82672;
  reg x82675, x82678, x82681, x82684, x82687, x82690, x82693, x82696;
  reg x82699, x82702, x82705, x82708, x82711, x82714, x82717, x82720;
  reg x82723, x82726, x82729, x82732, x82735, x82738, x82741, x82744;
  reg x82747, x82750, x82753, x82756, x82759, x82762, x82765, x82768;
  reg x82771, x82774, x82777, x82780, x82783, x82786, x82789, x82792;
  reg x82795, x82798, x82801, x82804, x82807, x82810, x82813, x82816;
  reg x82819, x82822, x82825, x82828, x82831, x82834, x82837, x82840;
  reg x82843, x82846, x82849, x82852, x82855, x82858, x82861, x82864;
  reg x82867, x82870, x82873, x82876, x82879, x82882, x82885, x82888;
  reg x82891, x82894, x82897, x82900, x82903, x82906, x82909, x82912;
  reg x82915, x82918, x82921, x82924, x82927, x82930, x82933, x82936;
  reg x82939, x82942, x82945, x82948, x82951, x82954, x82957, x82960;
  reg x82963, x82966, x82969, x82972, x82975, x82978, x82981, x82984;
  reg x82987, x82990, x82993, x82996, x82999, x83002, x83005, x83008;
  reg x83011, x83014, x83017, x83020, x83023, x83026, x83029, x83032;
  reg x83035, x83038, x83041, x83044, x83047, x83050, x83053, x83056;
  reg x83059, x83062, x83065, x83068, x83071, x83074, x83077, x83080;
  reg x83083, x83086, x83089, x83092, x83095, x83098, x83101, x83104;
  reg x83107, x83110, x83113, x83116, x83119, x83122, x83125, x83128;
  reg x83131, x83134, x83137, x83140, x83143, x83146, x83149, x83152;
  reg x83155, x83158, x83161, x83164, x83167, x83170, x83173, x83176;
  reg x83179, x83182, x83185, x83188, x83191, x83194, x83197, x83200;
  reg x83203, x83206, x83209, x83212, x83215, x83218, x83221, x83224;
  reg x83227, x83230, x83233, x83236, x83239, x83242, x83245, x83248;
  reg x83251, x83254, x83257, x83260, x83263, x83266, x83269, x83272;
  reg x83275, x83278, x83281, x83284, x83287, x83290, x83293, x83296;
  reg x83299, x83302, x83305, x83308, x83311, x83314, x83317, x83320;
  reg x83323, x83326, x83329, x83332, x83335, x83338, x83341, x83344;
  reg x83347, x83352, x83357, x83362, x83367, x83372, x83377, x83382;

  wire x61684;
  wire x61428;
  wire x61429;
  wire x61430;
  wire x61431;
  wire x61432;
  wire x61433;
  wire x61434;
  wire x61435;
  wire x61436;
  wire x61437;
  wire x61438;
  wire x61439;
  wire x61440;
  wire x61441;
  wire x61442;
  wire x61443;
  wire x61444;
  wire x61445;
  wire x61446;
  wire x61447;
  wire x61448;
  wire x61449;
  wire x61450;
  wire x61451;
  wire x61452;
  wire x61453;
  wire x61454;
  wire x61455;
  wire x61456;
  wire x61457;
  wire x61458;
  wire x61459;
  wire x61460;
  wire x61461;
  wire x61462;
  wire x61463;
  wire x61464;
  wire x61465;
  wire x61466;
  wire x61467;
  wire x61468;
  wire x61469;
  wire x61470;
  wire x61471;
  wire x61472;
  wire x61473;
  wire x61474;
  wire x61475;
  wire x61476;
  wire x61477;
  wire x61478;
  wire x61479;
  wire x61480;
  wire x61481;
  wire x61482;
  wire x61483;
  wire x61484;
  wire x61485;
  wire x61486;
  wire x61487;
  wire x61488;
  wire x61489;
  wire x61490;
  wire x61491;
  wire x61492;
  wire x61493;
  wire x61494;
  wire x61495;
  wire x61496;
  wire x61497;
  wire x61498;
  wire x61499;
  wire x61500;
  wire x61501;
  wire x61502;
  wire x61503;
  wire x61504;
  wire x61505;
  wire x61506;
  wire x61507;
  wire x61508;
  wire x61509;
  wire x61510;
  wire x61511;
  wire x61512;
  wire x61513;
  wire x61514;
  wire x61515;
  wire x61516;
  wire x61517;
  wire x61518;
  wire x61519;
  wire x61520;
  wire x61521;
  wire x61522;
  wire x61523;
  wire x61524;
  wire x61525;
  wire x61526;
  wire x61527;
  wire x61528;
  wire x61529;
  wire x61530;
  wire x61531;
  wire x61532;
  wire x61533;
  wire x61534;
  wire x61535;
  wire x61536;
  wire x61537;
  wire x61538;
  wire x61539;
  wire x61540;
  wire x61541;
  wire x61542;
  wire x61543;
  wire x61544;
  wire x61545;
  wire x61546;
  wire x61547;
  wire x61548;
  wire x61549;
  wire x61550;
  wire x61551;
  wire x61552;
  wire x61553;
  wire x61554;
  wire x61555;
  wire x61556;
  wire x61557;
  wire x61558;
  wire x61559;
  wire x61560;
  wire x61561;
  wire x61562;
  wire x61563;
  wire x61564;
  wire x61565;
  wire x61566;
  wire x61567;
  wire x61568;
  wire x61569;
  wire x61570;
  wire x61571;
  wire x61572;
  wire x61573;
  wire x61574;
  wire x61575;
  wire x61576;
  wire x61577;
  wire x61578;
  wire x61579;
  wire x61580;
  wire x61581;
  wire x61582;
  wire x61583;
  wire x61584;
  wire x61585;
  wire x61586;
  wire x61587;
  wire x61588;
  wire x61589;
  wire x61590;
  wire x61591;
  wire x61592;
  wire x61593;
  wire x61594;
  wire x61595;
  wire x61596;
  wire x61597;
  wire x61598;
  wire x61599;
  wire x61600;
  wire x61601;
  wire x61602;
  wire x61603;
  wire x61604;
  wire x61605;
  wire x61606;
  wire x61607;
  wire x61608;
  wire x61609;
  wire x61610;
  wire x61611;
  wire x61612;
  wire x61613;
  wire x61614;
  wire x61615;
  wire x61616;
  wire x61617;
  wire x61618;
  wire x61619;
  wire x61620;
  wire x61621;
  wire x61622;
  wire x61623;
  wire x61624;
  wire x61625;
  wire x61626;
  wire x61627;
  wire x61628;
  wire x61629;
  wire x61630;
  wire x61631;
  wire x61632;
  wire x61633;
  wire x61634;
  wire x61635;
  wire x61636;
  wire x61637;
  wire x61638;
  wire x61639;
  wire x61640;
  wire x61641;
  wire x61642;
  wire x61643;
  wire x61644;
  wire x61645;
  wire x61646;
  wire x61647;
  wire x61648;
  wire x61649;
  wire x61650;
  wire x61651;
  wire x61652;
  wire x61653;
  wire x61654;
  wire x61655;
  wire x61656;
  wire x61657;
  wire x61658;
  wire x61659;
  wire x61660;
  wire x61661;
  wire x61662;
  wire x61663;
  wire x61664;
  wire x61665;
  wire x61666;
  wire x61667;
  wire x61668;
  wire x61669;
  wire x61670;
  wire x61671;
  wire x61672;
  wire x61673;
  wire x61674;
  wire x61675;
  wire x61676;
  wire x61677;
  wire x61678;
  wire x61679;
  wire x61680;
  wire x61681;
  wire x61682;
  wire x61683;
  wire x66601;
  wire x66473;
  wire x66474;
  wire x66475;
  wire x66476;
  wire x66477;
  wire x66478;
  wire x66479;
  wire x66480;
  wire x66481;
  wire x66482;
  wire x66483;
  wire x66484;
  wire x66485;
  wire x66486;
  wire x66487;
  wire x66488;
  wire x66489;
  wire x66490;
  wire x66491;
  wire x66492;
  wire x66493;
  wire x66494;
  wire x66495;
  wire x66496;
  wire x66497;
  wire x66498;
  wire x66499;
  wire x66500;
  wire x66501;
  wire x66502;
  wire x66503;
  wire x66504;
  wire x66505;
  wire x66506;
  wire x66507;
  wire x66508;
  wire x66509;
  wire x66510;
  wire x66511;
  wire x66512;
  wire x66513;
  wire x66514;
  wire x66515;
  wire x66516;
  wire x66517;
  wire x66518;
  wire x66519;
  wire x66520;
  wire x66521;
  wire x66522;
  wire x66523;
  wire x66524;
  wire x66525;
  wire x66526;
  wire x66527;
  wire x66528;
  wire x66529;
  wire x66530;
  wire x66531;
  wire x66532;
  wire x66533;
  wire x66534;
  wire x66535;
  wire x66536;
  wire x66537;
  wire x66538;
  wire x66539;
  wire x66540;
  wire x66541;
  wire x66542;
  wire x66543;
  wire x66544;
  wire x66545;
  wire x66546;
  wire x66547;
  wire x66548;
  wire x66549;
  wire x66550;
  wire x66551;
  wire x66552;
  wire x66553;
  wire x66554;
  wire x66555;
  wire x66556;
  wire x66557;
  wire x66558;
  wire x66559;
  wire x66560;
  wire x66561;
  wire x66562;
  wire x66563;
  wire x66564;
  wire x66565;
  wire x66566;
  wire x66567;
  wire x66568;
  wire x66569;
  wire x66570;
  wire x66571;
  wire x66572;
  wire x66573;
  wire x66574;
  wire x66575;
  wire x66576;
  wire x66577;
  wire x66578;
  wire x66579;
  wire x66580;
  wire x66581;
  wire x66582;
  wire x66583;
  wire x66584;
  wire x66585;
  wire x66586;
  wire x66587;
  wire x66588;
  wire x66589;
  wire x66590;
  wire x66591;
  wire x66592;
  wire x66593;
  wire x66594;
  wire x66595;
  wire x66596;
  wire x66597;
  wire x66598;
  wire x66599;
  wire x66600;
  wire x67594;
  wire x67466;
  wire x67467;
  wire x67468;
  wire x67469;
  wire x67470;
  wire x67471;
  wire x67472;
  wire x67473;
  wire x67474;
  wire x67475;
  wire x67476;
  wire x67477;
  wire x67478;
  wire x67479;
  wire x67480;
  wire x67481;
  wire x67482;
  wire x67483;
  wire x67484;
  wire x67485;
  wire x67486;
  wire x67487;
  wire x67488;
  wire x67489;
  wire x67490;
  wire x67491;
  wire x67492;
  wire x67493;
  wire x67494;
  wire x67495;
  wire x67496;
  wire x67497;
  wire x67498;
  wire x67499;
  wire x67500;
  wire x67501;
  wire x67502;
  wire x67503;
  wire x67504;
  wire x67505;
  wire x67506;
  wire x67507;
  wire x67508;
  wire x67509;
  wire x67510;
  wire x67511;
  wire x67512;
  wire x67513;
  wire x67514;
  wire x67515;
  wire x67516;
  wire x67517;
  wire x67518;
  wire x67519;
  wire x67520;
  wire x67521;
  wire x67522;
  wire x67523;
  wire x67524;
  wire x67525;
  wire x67526;
  wire x67527;
  wire x67528;
  wire x67529;
  wire x67530;
  wire x67531;
  wire x67532;
  wire x67533;
  wire x67534;
  wire x67535;
  wire x67536;
  wire x67537;
  wire x67538;
  wire x67539;
  wire x67540;
  wire x67541;
  wire x67542;
  wire x67543;
  wire x67544;
  wire x67545;
  wire x67546;
  wire x67547;
  wire x67548;
  wire x67549;
  wire x67550;
  wire x67551;
  wire x67552;
  wire x67553;
  wire x67554;
  wire x67555;
  wire x67556;
  wire x67557;
  wire x67558;
  wire x67559;
  wire x67560;
  wire x67561;
  wire x67562;
  wire x67563;
  wire x67564;
  wire x67565;
  wire x67566;
  wire x67567;
  wire x67568;
  wire x67569;
  wire x67570;
  wire x67571;
  wire x67572;
  wire x67573;
  wire x67574;
  wire x67575;
  wire x67576;
  wire x67577;
  wire x67578;
  wire x67579;
  wire x67580;
  wire x67581;
  wire x67582;
  wire x67583;
  wire x67584;
  wire x67585;
  wire x67586;
  wire x67587;
  wire x67588;
  wire x67589;
  wire x67590;
  wire x67591;
  wire x67592;
  wire x67593;

  wire ram_w0;
  wire [7:0] ram_qa0;
  reg  [31:0] ram_q0;
  wire [7:0] ram_da0;
  wire [31:0] ram_d0;
  wire ram_w1;
  wire [7:0] ram_qa1;
  reg  [31:0] ram_q1;
  wire [7:0] ram_da1;
  wire [31:0] ram_d1;
  wire ram_w2;
  wire [7:0] ram_qa2;
  reg  [31:0] ram_q2;
  wire [7:0] ram_da2;
  wire [31:0] ram_d2;
  wire ram_w3;
  wire [7:0] ram_qa3;
  reg  [31:0] ram_q3;
  wire [7:0] ram_da3;
  wire [31:0] ram_d3;

  wire x2, x9, x10, x12, x14, x16, x17, x18;
  wire x20, x21, x22, x24, x25, x26, x28, x29;
  wire x30, x32, x33, x34, x36, x37, x38, x40;
  wire x41, x42, x43, x44, x45, x46, x47, x48;
  wire x49, x50, x51, x52, x53, x54, x55, x56;
  wire x57, x94, x95, x97, x99, x101, x103, x105;
  wire x107, x109, x111, x113, x115, x117, x119, x121;
  wire x123, x125, x127, x129, x131, x133, x135, x137;
  wire x139, x141, x143, x145, x147, x149, x150, x151;
  wire x153, x155, x157, x159, x161, x163, x165, x167;
  wire x169, x171, x173, x175, x177, x179, x181, x183;
  wire x185, x187, x189, x191, x193, x195, x197, x199;
  wire x201, x202, x203, x204, x205, x207, x209, x211;
  wire x213, x215, x217, x219, x221, x223, x225, x227;
  wire x229, x231, x233, x235, x237, x239, x241, x243;
  wire x245, x247, x248, x249, x250, x251, x252, x253;
  wire x254, x255, x257, x259, x261, x263, x265, x267;
  wire x269, x271, x273, x275, x277, x279, x281, x282;
  wire x283, x284, x285, x286, x287, x288, x289, x290;
  wire x291, x292, x293, x294, x295, x297, x298, x299;
  wire x301, x302, x303, x305, x306, x307, x309, x310;
  wire x311, x313, x314, x315, x317, x318, x319, x321;
  wire x322, x323, x325, x326, x327, x329, x330, x331;
  wire x333, x334, x335, x337, x338, x339, x341, x342;
  wire x343, x345, x346, x347, x349, x350, x351, x353;
  wire x354, x355, x357, x358, x359, x361, x362, x363;
  wire x365, x366, x367, x369, x370, x371, x373, x374;
  wire x375, x377, x378, x379, x381, x382, x383, x385;
  wire x386, x387, x389, x390, x391, x393, x394, x395;
  wire x397, x398, x399, x401, x402, x403, x405, x406;
  wire x407, x409, x411, x412, x413, x414, x415, x416;
  wire x417, x418, x419, x420, x421, x422, x423, x424;
  wire x425, x426, x427, x428, x429, x430, x431, x432;
  wire x433, x434, x435, x436, x437, x438, x439, x440;
  wire x441, x442, x443, x444, x445, x446, x447, x448;
  wire x449, x450, x451, x452, x453, x454, x455, x456;
  wire x457, x458, x459, x460, x461, x462, x463, x464;
  wire x465, x466, x467, x468, x469, x470, x471, x472;
  wire x473, x474, x475, x476, x477, x478, x479, x480;
  wire x481, x482, x483, x484, x485, x486, x487, x488;
  wire x489, x490, x491, x492, x493, x494, x495, x496;
  wire x497, x498, x499, x500, x501, x502, x503, x504;
  wire x505, x506, x507, x508, x509, x510, x511, x512;
  wire x513, x514, x515, x516, x517, x518, x519, x520;
  wire x521, x522, x523, x524, x525, x526, x527, x528;
  wire x529, x530, x531, x532, x533, x534, x535, x536;
  wire x537, x538, x539, x540, x541, x542, x543, x544;
  wire x545, x546, x547, x548, x549, x550, x551, x552;
  wire x553, x554, x555, x556, x557, x558, x559, x560;
  wire x561, x562, x563, x564, x565, x566, x567, x568;
  wire x569, x570, x571, x572, x573, x574, x575, x576;
  wire x577, x578, x579, x580, x581, x582, x583, x584;
  wire x585, x586, x587, x588, x589, x590, x591, x592;
  wire x593, x594, x595, x596, x597, x598, x599, x600;
  wire x601, x638, x639, x641, x642, x643, x645, x646;
  wire x647, x649, x650, x651, x653, x655, x657, x658;
  wire x659, x660, x661, x662, x663, x664, x665, x666;
  wire x667, x668, x669, x670, x671, x672, x673, x679;
  wire x680, x681, x682, x683, x684, x685, x686, x687;
  wire x688, x689, x690, x691, x692, x693, x694, x695;
  wire x696, x697, x698, x699, x700, x701, x702, x703;
  wire x704, x705, x706, x707, x708, x709, x710, x711;
  wire x712, x713, x714, x715, x716, x717, x718, x719;
  wire x720, x721, x722, x723, x724, x725, x726, x727;
  wire x728, x729, x730, x731, x732, x733, x734, x735;
  wire x736, x737, x738, x739, x740, x741, x742, x743;
  wire x744, x745, x746, x747, x748, x749, x750, x751;
  wire x752, x753, x754, x755, x756, x757, x758, x759;
  wire x760, x761, x762, x763, x764, x765, x766, x767;
  wire x768, x769, x770, x771, x772, x773, x774, x775;
  wire x776, x777, x778, x779, x780, x781, x782, x783;
  wire x784, x785, x786, x787, x788, x789, x790, x791;
  wire x792, x793, x794, x795, x796, x797, x798, x799;
  wire x800, x801, x802, x803, x804, x805, x806, x807;
  wire x808, x809, x810, x811, x812, x813, x814, x815;
  wire x816, x817, x818, x819, x820, x821, x822, x823;
  wire x824, x825, x826, x827, x828, x829, x830, x831;
  wire x832, x833, x834, x835, x836, x837, x838, x839;
  wire x840, x841, x842, x843, x844, x845, x846, x847;
  wire x848, x849, x850, x851, x852, x853, x854, x855;
  wire x856, x857, x858, x859, x860, x861, x862, x863;
  wire x864, x865, x866, x867, x868, x869, x870, x871;
  wire x872, x873, x874, x875, x876, x877, x878, x879;
  wire x880, x881, x882, x883, x884, x885, x886, x887;
  wire x888, x889, x890, x891, x892, x893, x894, x895;
  wire x896, x897, x898, x899, x900, x901, x902, x903;
  wire x904, x905, x906, x907, x908, x909, x910, x911;
  wire x912, x913, x914, x915, x916, x917, x918, x919;
  wire x920, x921, x922, x923, x924, x925, x926, x927;
  wire x928, x929, x930, x931, x932, x933, x934, x935;
  wire x936, x937, x938, x939, x940, x941, x942, x943;
  wire x944, x945, x946, x947, x948, x949, x950, x951;
  wire x952, x953, x954, x955, x956, x957, x958, x959;
  wire x960, x961, x962, x963, x964, x965, x966, x967;
  wire x968, x969, x970, x971, x972, x973, x974, x975;
  wire x976, x977, x978, x979, x980, x981, x982, x983;
  wire x984, x985, x986, x987, x988, x989, x990, x991;
  wire x992, x993, x994, x995, x996, x997, x998, x999;
  wire x1002, x1004, x1006, x1008, x1010, x1013, x1015, x1017;
  wire x1019, x1021, x1023, x1025, x1027, x1029, x1030, x1032;
  wire x1034, x1036, x1037, x1039, x1041, x1043, x1044, x1045;
  wire x1047, x1049, x1051, x1053, x1054, x1055, x1056, x1057;
  wire x1058, x1060, x1061, x1063, x1064, x1065, x1066, x1067;
  wire x1069, x1070, x1071, x1072, x1073, x1074, x1076, x1078;
  wire x1080, x1082, x1084, x1086, x1088, x1090, x1092, x1094;
  wire x1096, x1098, x1099, x1100, x1102, x1104, x1105, x1107;
  wire x1108, x1109, x1111, x1112, x1113, x1114, x1115, x1117;
  wire x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1126;
  wire x1128, x1130, x1132, x1134, x1136, x1138, x1140, x1142;
  wire x1143, x1144, x1146, x1147, x1149, x1150, x1151, x1153;
  wire x1154, x1155, x1156, x1157, x1158, x1160, x1165, x1166;
  wire x1167, x1171, x1173, x1174, x1176, x1178, x1182, x1184;
  wire x1185, x1187, x1189, x1191, x1192, x1195, x1197, x1199;
  wire x1202, x1204, x1206, x1208, x1211, x1213, x1215, x1217;
  wire x1219, x1221, x1223, x1225, x1227, x1229, x1230, x1231;
  wire x1233, x1235, x1236, x1237, x1239, x1241, x1242, x1243;
  wire x1245, x1247, x1248, x1249, x1251, x1253, x1254, x1255;
  wire x1257, x1259, x1260, x1261, x1263, x1265, x1266, x1267;
  wire x1269, x1271, x1272, x1273, x1275, x1277, x1278, x1279;
  wire x1283, x1285, x1286, x1287, x1289, x1291, x1292, x1293;
  wire x1295, x1297, x1298, x1299, x1301, x1303, x1304, x1305;
  wire x1307, x1309, x1310, x1311, x1313, x1315, x1316, x1317;
  wire x1319, x1321, x1322, x1323, x1325, x1327, x1328, x1329;
  wire x1331, x1333, x1334, x1335, x1337, x1339, x1340, x1341;
  wire x1343, x1345, x1346, x1347, x1349, x1351, x1352, x1353;
  wire x1355, x1357, x1358, x1359, x1361, x1363, x1364, x1365;
  wire x1367, x1369, x1370, x1371, x1373, x1375, x1376, x1377;
  wire x1381, x1383, x1384, x1385, x1387, x1389, x1390, x1391;
  wire x1393, x1395, x1396, x1397, x1399, x1401, x1402, x1403;
  wire x1405, x1407, x1408, x1409, x1411, x1413, x1414, x1415;
  wire x1417, x1419, x1420, x1421, x1423, x1425, x1426, x1427;
  wire x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435;
  wire x1436, x1438, x1439, x1440, x1441, x1442, x1443, x1445;
  wire x1446, x1447, x1449, x1450, x1451, x1452, x1453, x1454;
  wire x1455, x1456, x1457, x1458, x1459, x1460, x1462, x1463;
  wire x1464, x1465, x1466, x1467, x1469, x1470, x1471, x1473;
  wire x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481;
  wire x1482, x1483, x1484, x1486, x1487, x1488, x1489, x1490;
  wire x1491, x1493, x1494, x1495, x1496, x1497, x1498, x1499;
  wire x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507;
  wire x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515;
  wire x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523;
  wire x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531;
  wire x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539;
  wire x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547;
  wire x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555;
  wire x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563;
  wire x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571;
  wire x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579;
  wire x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587;
  wire x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595;
  wire x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603;
  wire x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611;
  wire x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619;
  wire x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627;
  wire x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635;
  wire x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643;
  wire x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651;
  wire x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659;
  wire x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667;
  wire x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675;
  wire x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683;
  wire x1685, x1687, x1689, x1691, x1692, x1694, x1696, x1698;
  wire x1700, x1702, x1704, x1706, x1708, x1710, x1712, x1713;
  wire x1715, x1716, x1718, x1719, x1720, x1721, x1722, x1723;
  wire x1726, x1728, x1730, x1733, x1735, x1737, x1739, x1742;
  wire x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750;
  wire x1752, x1753, x1755, x1756, x1760, x1762, x1763, x1765;
  wire x1766, x1770, x1772, x1773, x1775, x1776, x1780, x1782;
  wire x1783, x1785, x1786, x1790, x1792, x1793, x1795, x1796;
  wire x1800, x1802, x1803, x1805, x1806, x1810, x1812, x1813;
  wire x1815, x1816, x1820, x1822, x1823, x1825, x1826, x1830;
  wire x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838;
  wire x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846;
  wire x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854;
  wire x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862;
  wire x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870;
  wire x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878;
  wire x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886;
  wire x1887, x1888, x1889, x1890, x1891, x1892, x1894, x1895;
  wire x1898, x1900, x1909, x1911, x1912, x1913, x1915, x1916;
  wire x1917, x1919, x1920, x1921, x1923, x1924, x1925, x1927;
  wire x1928, x1929, x1931, x1932, x1933, x1935, x1937, x1938;
  wire x1939, x1941, x1942, x1943, x1945, x1946, x1947, x1949;
  wire x1950, x1951, x1953, x1954, x1955, x1957, x1958, x1959;
  wire x1961, x1963, x1964, x1965, x1967, x1968, x1969, x1971;
  wire x1972, x1973, x1975, x1976, x1977, x1979, x1980, x1981;
  wire x1983, x1984, x1985, x1987, x1989, x1990, x1991, x1993;
  wire x1994, x1995, x1997, x1998, x1999, x2001, x2002, x2003;
  wire x2005, x2006, x2007, x2009, x2010, x2011, x2013, x2015;
  wire x2016, x2017, x2019, x2020, x2021, x2023, x2024, x2025;
  wire x2027, x2028, x2029, x2031, x2032, x2033, x2035, x2036;
  wire x2037, x2039, x2041, x2042, x2043, x2045, x2046, x2047;
  wire x2049, x2050, x2051, x2053, x2054, x2055, x2057, x2058;
  wire x2059, x2061, x2062, x2063, x2065, x2067, x2068, x2069;
  wire x2071, x2072, x2073, x2075, x2076, x2077, x2079, x2080;
  wire x2081, x2083, x2084, x2085, x2087, x2088, x2089, x2091;
  wire x2093, x2094, x2095, x2097, x2098, x2099, x2101, x2102;
  wire x2103, x2105, x2106, x2107, x2109, x2110, x2111, x2113;
  wire x2114, x2115, x2117, x2118, x2119, x2120, x2121, x2122;
  wire x2123, x2124, x2125, x2126, x2127, x2128, x2129, x2130;
  wire x2131, x2132, x2133, x2134, x2135, x2136, x2137, x2138;
  wire x2139, x2140, x2141, x2142, x2143, x2144, x2145, x2146;
  wire x2147, x2148, x2149, x2150, x2151, x2152, x2153, x2154;
  wire x2155, x2156, x2157, x2158, x2159, x2160, x2161, x2162;
  wire x2163, x2164, x2165, x2166, x2167, x2168, x2169, x2170;
  wire x2171, x2172, x2173, x2174, x2175, x2176, x2177, x2178;
  wire x2179, x2180, x2181, x2182, x2183, x2184, x2185, x2186;
  wire x2187, x2188, x2189, x2190, x2191, x2192, x2193, x2194;
  wire x2195, x2196, x2197, x2198, x2199, x2200, x2201, x2202;
  wire x2203, x2204, x2205, x2206, x2207, x2208, x2209, x2210;
  wire x2211, x2212, x2213, x2214, x2215, x2216, x2217, x2218;
  wire x2219, x2220, x2221, x2222, x2223, x2224, x2225, x2226;
  wire x2227, x2228, x2229, x2230, x2231, x2232, x2233, x2234;
  wire x2235, x2236, x2237, x2238, x2239, x2240, x2241, x2242;
  wire x2243, x2245, x2246, x2248, x2249, x2251, x2252, x2254;
  wire x2255, x2257, x2258, x2259, x2260, x2261, x2262, x2263;
  wire x2264, x2265, x2266, x2268, x2269, x2270, x2271, x2272;
  wire x2273, x2274, x2275, x2276, x2277, x2280, x2282, x2284;
  wire x2287, x2289, x2291, x2293, x2296, x2298, x2300, x2302;
  wire x2304, x2306, x2308, x2310, x2312, x2314, x2315, x2316;
  wire x2318, x2319, x2320, x2322, x2323, x2324, x2326, x2327;
  wire x2328, x2330, x2331, x2332, x2334, x2335, x2336, x2338;
  wire x2339, x2340, x2342, x2343, x2344, x2346, x2347, x2348;
  wire x2350, x2351, x2352, x2354, x2355, x2356, x2358, x2359;
  wire x2360, x2362, x2363, x2364, x2366, x2367, x2368, x2370;
  wire x2371, x2372, x2374, x2375, x2376, x2378, x2379, x2380;
  wire x2382, x2383, x2384, x2386, x2387, x2388, x2390, x2391;
  wire x2392, x2394, x2395, x2396, x2398, x2399, x2400, x2402;
  wire x2403, x2404, x2406, x2407, x2408, x2410, x2411, x2412;
  wire x2414, x2415, x2416, x2418, x2419, x2420, x2422, x2423;
  wire x2424, x2426, x2427, x2428, x2430, x2431, x2432, x2434;
  wire x2435, x2436, x2438, x2439, x2440, x2442, x2444, x2445;
  wire x2446, x2448, x2449, x2450, x2452, x2453, x2454, x2456;
  wire x2457, x2458, x2460, x2461, x2462, x2464, x2465, x2466;
  wire x2468, x2469, x2470, x2472, x2473, x2474, x2476, x2477;
  wire x2478, x2480, x2481, x2482, x2484, x2485, x2486, x2488;
  wire x2489, x2490, x2492, x2493, x2494, x2496, x2497, x2498;
  wire x2500, x2501, x2502, x2504, x2505, x2506, x2508, x2509;
  wire x2510, x2512, x2513, x2514, x2516, x2517, x2518, x2520;
  wire x2521, x2522, x2524, x2525, x2526, x2528, x2529, x2530;
  wire x2532, x2533, x2534, x2536, x2537, x2538, x2540, x2541;
  wire x2542, x2544, x2545, x2546, x2548, x2549, x2550, x2552;
  wire x2553, x2554, x2556, x2557, x2558, x2560, x2561, x2562;
  wire x2564, x2565, x2566, x2568, x2569, x2570, x2572, x2574;
  wire x2575, x2576, x2578, x2579, x2580, x2582, x2583, x2584;
  wire x2586, x2587, x2588, x2590, x2591, x2592, x2594, x2595;
  wire x2596, x2598, x2599, x2600, x2602, x2603, x2604, x2606;
  wire x2607, x2608, x2610, x2611, x2612, x2614, x2615, x2616;
  wire x2618, x2619, x2620, x2622, x2623, x2624, x2626, x2627;
  wire x2628, x2630, x2631, x2632, x2634, x2635, x2636, x2638;
  wire x2639, x2640, x2642, x2643, x2644, x2646, x2647, x2648;
  wire x2650, x2651, x2652, x2654, x2655, x2656, x2658, x2659;
  wire x2660, x2662, x2663, x2664, x2666, x2667, x2668, x2670;
  wire x2671, x2672, x2674, x2675, x2676, x2678, x2679, x2680;
  wire x2682, x2683, x2684, x2686, x2687, x2688, x2690, x2691;
  wire x2692, x2694, x2695, x2696, x2698, x2699, x2700, x2702;
  wire x2704, x2705, x2706, x2708, x2709, x2710, x2712, x2713;
  wire x2714, x2716, x2717, x2718, x2720, x2721, x2722, x2724;
  wire x2725, x2726, x2728, x2729, x2730, x2732, x2733, x2734;
  wire x2736, x2737, x2738, x2740, x2741, x2742, x2744, x2745;
  wire x2746, x2748, x2749, x2750, x2752, x2753, x2754, x2756;
  wire x2757, x2758, x2760, x2761, x2762, x2764, x2765, x2766;
  wire x2768, x2769, x2770, x2772, x2773, x2774, x2776, x2777;
  wire x2778, x2780, x2781, x2782, x2784, x2785, x2786, x2788;
  wire x2789, x2790, x2792, x2793, x2794, x2796, x2797, x2798;
  wire x2800, x2801, x2802, x2804, x2805, x2806, x2808, x2809;
  wire x2810, x2812, x2813, x2814, x2816, x2817, x2818, x2820;
  wire x2821, x2822, x2824, x2825, x2826, x2828, x2829, x2830;
  wire x2832, x2834, x2835, x2836, x2838, x2839, x2840, x2842;
  wire x2843, x2844, x2846, x2847, x2848, x2850, x2851, x2852;
  wire x2854, x2855, x2856, x2858, x2859, x2860, x2862, x2863;
  wire x2864, x2866, x2867, x2868, x2870, x2871, x2872, x2874;
  wire x2875, x2876, x2878, x2879, x2880, x2882, x2883, x2884;
  wire x2886, x2887, x2888, x2890, x2891, x2892, x2894, x2895;
  wire x2896, x2898, x2899, x2900, x2902, x2903, x2904, x2906;
  wire x2907, x2908, x2910, x2911, x2912, x2914, x2915, x2916;
  wire x2918, x2919, x2920, x2922, x2923, x2924, x2926, x2927;
  wire x2928, x2930, x2931, x2932, x2934, x2935, x2936, x2938;
  wire x2939, x2940, x2942, x2943, x2944, x2946, x2947, x2948;
  wire x2950, x2951, x2952, x2954, x2955, x2956, x2958, x2959;
  wire x2960, x2962, x2964, x2965, x2966, x2968, x2969, x2970;
  wire x2972, x2973, x2974, x2976, x2977, x2978, x2980, x2981;
  wire x2982, x2984, x2985, x2986, x2988, x2989, x2990, x2992;
  wire x2993, x2994, x2996, x2997, x2998, x3000, x3001, x3002;
  wire x3004, x3005, x3006, x3008, x3009, x3010, x3012, x3013;
  wire x3014, x3016, x3017, x3018, x3020, x3021, x3022, x3024;
  wire x3025, x3026, x3028, x3029, x3030, x3032, x3033, x3034;
  wire x3036, x3037, x3038, x3040, x3041, x3042, x3044, x3045;
  wire x3046, x3048, x3049, x3050, x3052, x3053, x3054, x3056;
  wire x3057, x3058, x3060, x3061, x3062, x3064, x3065, x3066;
  wire x3068, x3069, x3070, x3072, x3073, x3074, x3076, x3077;
  wire x3078, x3080, x3081, x3082, x3084, x3085, x3086, x3088;
  wire x3089, x3090, x3092, x3094, x3095, x3096, x3098, x3099;
  wire x3100, x3102, x3103, x3104, x3106, x3107, x3108, x3110;
  wire x3111, x3112, x3114, x3115, x3116, x3118, x3119, x3120;
  wire x3122, x3123, x3124, x3126, x3127, x3128, x3130, x3131;
  wire x3132, x3134, x3135, x3136, x3138, x3139, x3140, x3142;
  wire x3143, x3144, x3146, x3147, x3148, x3150, x3151, x3152;
  wire x3154, x3155, x3156, x3158, x3159, x3160, x3162, x3163;
  wire x3164, x3166, x3167, x3168, x3170, x3171, x3172, x3174;
  wire x3175, x3176, x3178, x3179, x3180, x3182, x3183, x3184;
  wire x3186, x3187, x3188, x3190, x3191, x3192, x3194, x3195;
  wire x3196, x3198, x3199, x3200, x3202, x3203, x3204, x3206;
  wire x3207, x3208, x3210, x3211, x3212, x3214, x3215, x3216;
  wire x3218, x3219, x3220, x3222, x3224, x3225, x3226, x3228;
  wire x3229, x3230, x3232, x3233, x3234, x3236, x3237, x3238;
  wire x3240, x3241, x3242, x3244, x3245, x3246, x3248, x3249;
  wire x3250, x3252, x3253, x3254, x3256, x3257, x3258, x3260;
  wire x3261, x3262, x3264, x3265, x3266, x3268, x3269, x3270;
  wire x3272, x3273, x3274, x3276, x3277, x3278, x3280, x3281;
  wire x3282, x3284, x3285, x3286, x3288, x3289, x3290, x3292;
  wire x3293, x3294, x3296, x3297, x3298, x3300, x3301, x3302;
  wire x3304, x3305, x3306, x3308, x3309, x3310, x3312, x3313;
  wire x3314, x3316, x3317, x3318, x3320, x3321, x3322, x3324;
  wire x3325, x3326, x3328, x3329, x3330, x3332, x3333, x3334;
  wire x3336, x3337, x3338, x3340, x3341, x3342, x3344, x3345;
  wire x3346, x3348, x3349, x3350, x3352, x3354, x3355, x3356;
  wire x3360, x3361, x3362, x3364, x3365, x3366, x3368, x3369;
  wire x3370, x3372, x3373, x3374, x3376, x3377, x3378, x3380;
  wire x3381, x3382, x3384, x3385, x3386, x3388, x3389, x3390;
  wire x3392, x3393, x3394, x3396, x3397, x3398, x3400, x3401;
  wire x3402, x3404, x3405, x3406, x3408, x3409, x3410, x3412;
  wire x3413, x3414, x3416, x3417, x3418, x3420, x3421, x3422;
  wire x3424, x3425, x3426, x3428, x3429, x3430, x3432, x3433;
  wire x3434, x3436, x3437, x3438, x3440, x3441, x3442, x3444;
  wire x3445, x3446, x3448, x3449, x3450, x3452, x3453, x3454;
  wire x3456, x3457, x3458, x3460, x3461, x3462, x3464, x3465;
  wire x3466, x3468, x3469, x3470, x3472, x3473, x3474, x3476;
  wire x3477, x3478, x3480, x3481, x3482, x3484, x3486, x3487;
  wire x3488, x3490, x3491, x3492, x3494, x3495, x3496, x3498;
  wire x3499, x3500, x3502, x3503, x3504, x3506, x3507, x3508;
  wire x3510, x3511, x3512, x3514, x3515, x3516, x3518, x3519;
  wire x3520, x3522, x3523, x3524, x3526, x3527, x3528, x3530;
  wire x3531, x3532, x3534, x3535, x3536, x3538, x3539, x3540;
  wire x3542, x3543, x3544, x3546, x3547, x3548, x3550, x3551;
  wire x3552, x3554, x3555, x3556, x3558, x3559, x3560, x3562;
  wire x3563, x3564, x3566, x3567, x3568, x3570, x3571, x3572;
  wire x3574, x3575, x3576, x3578, x3579, x3580, x3582, x3583;
  wire x3584, x3586, x3587, x3588, x3590, x3591, x3592, x3594;
  wire x3595, x3596, x3598, x3599, x3600, x3602, x3603, x3604;
  wire x3606, x3607, x3608, x3610, x3611, x3612, x3614, x3616;
  wire x3617, x3618, x3620, x3621, x3622, x3624, x3625, x3626;
  wire x3628, x3629, x3630, x3632, x3633, x3634, x3636, x3637;
  wire x3638, x3640, x3641, x3642, x3644, x3645, x3646, x3648;
  wire x3649, x3650, x3652, x3653, x3654, x3656, x3657, x3658;
  wire x3660, x3661, x3662, x3664, x3665, x3666, x3668, x3669;
  wire x3670, x3672, x3673, x3674, x3676, x3677, x3678, x3680;
  wire x3681, x3682, x3684, x3685, x3686, x3688, x3689, x3690;
  wire x3692, x3693, x3694, x3696, x3697, x3698, x3700, x3701;
  wire x3702, x3704, x3705, x3706, x3708, x3709, x3710, x3712;
  wire x3713, x3714, x3716, x3717, x3718, x3720, x3721, x3722;
  wire x3724, x3725, x3726, x3728, x3729, x3730, x3732, x3733;
  wire x3734, x3736, x3737, x3738, x3740, x3741, x3742, x3744;
  wire x3746, x3747, x3748, x3750, x3751, x3752, x3754, x3755;
  wire x3756, x3758, x3759, x3760, x3762, x3763, x3764, x3766;
  wire x3767, x3768, x3770, x3771, x3772, x3774, x3775, x3776;
  wire x3778, x3779, x3780, x3782, x3783, x3784, x3786, x3787;
  wire x3788, x3790, x3791, x3792, x3794, x3795, x3796, x3798;
  wire x3799, x3800, x3802, x3803, x3804, x3806, x3807, x3808;
  wire x3810, x3811, x3812, x3814, x3815, x3816, x3818, x3819;
  wire x3820, x3822, x3823, x3824, x3826, x3827, x3828, x3830;
  wire x3831, x3832, x3834, x3835, x3836, x3838, x3839, x3840;
  wire x3842, x3843, x3844, x3846, x3847, x3848, x3850, x3851;
  wire x3852, x3854, x3855, x3856, x3858, x3859, x3860, x3862;
  wire x3863, x3864, x3866, x3867, x3868, x3870, x3871, x3872;
  wire x3874, x3876, x3877, x3878, x3880, x3881, x3882, x3884;
  wire x3885, x3886, x3888, x3889, x3890, x3892, x3893, x3894;
  wire x3896, x3897, x3898, x3900, x3901, x3902, x3904, x3905;
  wire x3906, x3908, x3909, x3910, x3912, x3913, x3914, x3916;
  wire x3917, x3918, x3920, x3921, x3922, x3924, x3925, x3926;
  wire x3928, x3929, x3930, x3932, x3933, x3934, x3936, x3937;
  wire x3938, x3940, x3941, x3942, x3944, x3945, x3946, x3948;
  wire x3949, x3950, x3952, x3953, x3954, x3956, x3957, x3958;
  wire x3960, x3961, x3962, x3964, x3965, x3966, x3968, x3969;
  wire x3970, x3972, x3973, x3974, x3976, x3977, x3978, x3980;
  wire x3981, x3982, x3984, x3985, x3986, x3988, x3989, x3990;
  wire x3992, x3993, x3994, x3996, x3997, x3998, x4000, x4001;
  wire x4002, x4004, x4006, x4007, x4008, x4010, x4011, x4012;
  wire x4014, x4015, x4016, x4018, x4019, x4020, x4022, x4023;
  wire x4024, x4026, x4027, x4028, x4030, x4031, x4032, x4034;
  wire x4035, x4036, x4038, x4039, x4040, x4042, x4043, x4044;
  wire x4046, x4047, x4048, x4050, x4051, x4052, x4054, x4055;
  wire x4056, x4058, x4059, x4060, x4062, x4063, x4064, x4066;
  wire x4067, x4068, x4070, x4071, x4072, x4074, x4075, x4076;
  wire x4078, x4079, x4080, x4082, x4083, x4084, x4086, x4087;
  wire x4088, x4090, x4091, x4092, x4094, x4095, x4096, x4098;
  wire x4099, x4100, x4102, x4103, x4104, x4106, x4107, x4108;
  wire x4110, x4111, x4112, x4114, x4115, x4116, x4118, x4119;
  wire x4120, x4122, x4123, x4124, x4126, x4127, x4128, x4130;
  wire x4131, x4132, x4134, x4136, x4137, x4138, x4140, x4141;
  wire x4142, x4144, x4145, x4146, x4148, x4149, x4150, x4152;
  wire x4153, x4154, x4156, x4157, x4158, x4160, x4161, x4162;
  wire x4164, x4165, x4166, x4168, x4169, x4170, x4172, x4173;
  wire x4174, x4176, x4177, x4178, x4180, x4181, x4182, x4184;
  wire x4185, x4186, x4188, x4189, x4190, x4192, x4193, x4194;
  wire x4196, x4197, x4198, x4200, x4201, x4202, x4204, x4205;
  wire x4206, x4208, x4209, x4210, x4212, x4213, x4214, x4216;
  wire x4217, x4218, x4220, x4221, x4222, x4224, x4225, x4226;
  wire x4228, x4229, x4230, x4232, x4233, x4234, x4236, x4237;
  wire x4238, x4240, x4241, x4242, x4244, x4245, x4246, x4248;
  wire x4249, x4250, x4252, x4253, x4254, x4256, x4257, x4258;
  wire x4260, x4261, x4262, x4264, x4266, x4267, x4268, x4270;
  wire x4271, x4272, x4274, x4275, x4276, x4278, x4279, x4280;
  wire x4282, x4283, x4284, x4286, x4287, x4288, x4290, x4291;
  wire x4292, x4294, x4295, x4296, x4298, x4299, x4300, x4302;
  wire x4303, x4304, x4306, x4307, x4308, x4310, x4311, x4312;
  wire x4314, x4315, x4316, x4318, x4319, x4320, x4322, x4323;
  wire x4324, x4326, x4327, x4328, x4330, x4331, x4332, x4334;
  wire x4335, x4336, x4338, x4339, x4340, x4342, x4343, x4344;
  wire x4346, x4347, x4348, x4350, x4351, x4352, x4354, x4355;
  wire x4356, x4358, x4359, x4360, x4362, x4363, x4364, x4366;
  wire x4367, x4368, x4370, x4371, x4372, x4374, x4375, x4376;
  wire x4378, x4379, x4380, x4382, x4383, x4384, x4386, x4387;
  wire x4388, x4390, x4391, x4392, x4394, x4396, x4397, x4398;
  wire x4400, x4401, x4402, x4406, x4407, x4408, x4410, x4411;
  wire x4412, x4414, x4415, x4416, x4418, x4419, x4420, x4422;
  wire x4423, x4424, x4426, x4427, x4428, x4430, x4431, x4432;
  wire x4434, x4435, x4436, x4438, x4439, x4440, x4442, x4443;
  wire x4444, x4446, x4447, x4448, x4450, x4451, x4452, x4454;
  wire x4455, x4456, x4458, x4459, x4460, x4462, x4463, x4464;
  wire x4466, x4467, x4468, x4470, x4471, x4472, x4474, x4475;
  wire x4476, x4478, x4479, x4480, x4482, x4483, x4484, x4486;
  wire x4487, x4488, x4490, x4491, x4492, x4494, x4495, x4496;
  wire x4498, x4499, x4500, x4502, x4503, x4504, x4506, x4507;
  wire x4508, x4510, x4511, x4512, x4514, x4515, x4516, x4518;
  wire x4519, x4520, x4522, x4523, x4524, x4526, x4528, x4529;
  wire x4530, x4532, x4533, x4534, x4536, x4537, x4538, x4540;
  wire x4541, x4542, x4544, x4545, x4546, x4548, x4549, x4550;
  wire x4552, x4553, x4554, x4556, x4557, x4558, x4560, x4561;
  wire x4562, x4564, x4565, x4566, x4568, x4569, x4570, x4572;
  wire x4573, x4574, x4576, x4577, x4578, x4580, x4581, x4582;
  wire x4584, x4585, x4586, x4588, x4589, x4590, x4592, x4593;
  wire x4594, x4596, x4597, x4598, x4600, x4601, x4602, x4604;
  wire x4605, x4606, x4608, x4609, x4610, x4612, x4613, x4614;
  wire x4616, x4617, x4618, x4620, x4621, x4622, x4624, x4625;
  wire x4626, x4628, x4629, x4630, x4632, x4633, x4634, x4636;
  wire x4637, x4638, x4640, x4641, x4642, x4644, x4645, x4646;
  wire x4648, x4649, x4650, x4652, x4653, x4654, x4656, x4658;
  wire x4659, x4660, x4662, x4663, x4664, x4666, x4667, x4668;
  wire x4670, x4671, x4672, x4674, x4675, x4676, x4678, x4679;
  wire x4680, x4682, x4683, x4684, x4686, x4687, x4688, x4690;
  wire x4691, x4692, x4694, x4695, x4696, x4698, x4699, x4700;
  wire x4702, x4703, x4704, x4706, x4707, x4708, x4710, x4711;
  wire x4712, x4714, x4715, x4716, x4718, x4719, x4720, x4722;
  wire x4723, x4724, x4726, x4727, x4728, x4730, x4731, x4732;
  wire x4734, x4735, x4736, x4738, x4739, x4740, x4742, x4743;
  wire x4744, x4746, x4747, x4748, x4750, x4751, x4752, x4754;
  wire x4755, x4756, x4758, x4759, x4760, x4762, x4763, x4764;
  wire x4766, x4767, x4768, x4770, x4771, x4772, x4774, x4775;
  wire x4776, x4778, x4779, x4780, x4782, x4783, x4784, x4786;
  wire x4788, x4789, x4790, x4792, x4793, x4794, x4796, x4797;
  wire x4798, x4800, x4801, x4802, x4804, x4805, x4806, x4808;
  wire x4809, x4810, x4812, x4813, x4814, x4816, x4817, x4818;
  wire x4820, x4821, x4822, x4824, x4825, x4826, x4828, x4829;
  wire x4830, x4832, x4833, x4834, x4836, x4837, x4838, x4840;
  wire x4841, x4842, x4844, x4845, x4846, x4848, x4849, x4850;
  wire x4852, x4853, x4854, x4856, x4857, x4858, x4860, x4861;
  wire x4862, x4864, x4865, x4866, x4868, x4869, x4870, x4872;
  wire x4873, x4874, x4876, x4877, x4878, x4880, x4881, x4882;
  wire x4884, x4885, x4886, x4888, x4889, x4890, x4892, x4893;
  wire x4894, x4896, x4897, x4898, x4900, x4901, x4902, x4904;
  wire x4905, x4906, x4908, x4909, x4910, x4912, x4913, x4914;
  wire x4916, x4918, x4919, x4920, x4922, x4923, x4924, x4926;
  wire x4927, x4928, x4930, x4931, x4932, x4934, x4935, x4936;
  wire x4938, x4939, x4940, x4942, x4943, x4944, x4946, x4947;
  wire x4948, x4950, x4951, x4952, x4954, x4955, x4956, x4958;
  wire x4959, x4960, x4962, x4963, x4964, x4966, x4967, x4968;
  wire x4970, x4971, x4972, x4974, x4975, x4976, x4978, x4979;
  wire x4980, x4982, x4983, x4984, x4986, x4987, x4988, x4990;
  wire x4991, x4992, x4994, x4995, x4996, x4998, x4999, x5000;
  wire x5002, x5003, x5004, x5006, x5007, x5008, x5010, x5011;
  wire x5012, x5014, x5015, x5016, x5018, x5019, x5020, x5022;
  wire x5023, x5024, x5026, x5027, x5028, x5030, x5031, x5032;
  wire x5034, x5035, x5036, x5038, x5039, x5040, x5042, x5043;
  wire x5044, x5046, x5048, x5049, x5050, x5052, x5053, x5054;
  wire x5056, x5057, x5058, x5060, x5061, x5062, x5064, x5065;
  wire x5066, x5068, x5069, x5070, x5072, x5073, x5074, x5076;
  wire x5077, x5078, x5080, x5081, x5082, x5084, x5085, x5086;
  wire x5088, x5089, x5090, x5092, x5093, x5094, x5096, x5097;
  wire x5098, x5100, x5101, x5102, x5104, x5105, x5106, x5108;
  wire x5109, x5110, x5112, x5113, x5114, x5116, x5117, x5118;
  wire x5120, x5121, x5122, x5124, x5125, x5126, x5128, x5129;
  wire x5130, x5132, x5133, x5134, x5136, x5137, x5138, x5140;
  wire x5141, x5142, x5144, x5145, x5146, x5148, x5149, x5150;
  wire x5152, x5153, x5154, x5156, x5157, x5158, x5160, x5161;
  wire x5162, x5164, x5165, x5166, x5168, x5169, x5170, x5172;
  wire x5173, x5174, x5176, x5178, x5179, x5180, x5182, x5183;
  wire x5184, x5186, x5187, x5188, x5190, x5191, x5192, x5194;
  wire x5195, x5196, x5198, x5199, x5200, x5202, x5203, x5204;
  wire x5206, x5207, x5208, x5210, x5211, x5212, x5214, x5215;
  wire x5216, x5218, x5219, x5220, x5222, x5223, x5224, x5226;
  wire x5227, x5228, x5230, x5231, x5232, x5234, x5235, x5236;
  wire x5238, x5239, x5240, x5242, x5243, x5244, x5246, x5247;
  wire x5248, x5250, x5251, x5252, x5254, x5255, x5256, x5258;
  wire x5259, x5260, x5262, x5263, x5264, x5266, x5267, x5268;
  wire x5270, x5271, x5272, x5274, x5275, x5276, x5278, x5279;
  wire x5280, x5282, x5283, x5284, x5286, x5287, x5288, x5290;
  wire x5291, x5292, x5294, x5295, x5296, x5298, x5299, x5300;
  wire x5302, x5303, x5304, x5306, x5308, x5309, x5310, x5312;
  wire x5313, x5314, x5316, x5317, x5318, x5320, x5321, x5322;
  wire x5324, x5325, x5326, x5328, x5329, x5330, x5332, x5333;
  wire x5334, x5336, x5337, x5338, x5340, x5341, x5342, x5344;
  wire x5345, x5346, x5348, x5349, x5350, x5352, x5353, x5354;
  wire x5356, x5357, x5358, x5360, x5361, x5362, x5364, x5365;
  wire x5366, x5368, x5369, x5370, x5372, x5373, x5374, x5376;
  wire x5377, x5378, x5380, x5381, x5382, x5384, x5385, x5386;
  wire x5388, x5389, x5390, x5392, x5393, x5394, x5396, x5397;
  wire x5398, x5400, x5401, x5402, x5404, x5405, x5406, x5408;
  wire x5409, x5410, x5412, x5413, x5414, x5416, x5417, x5418;
  wire x5420, x5421, x5422, x5424, x5425, x5426, x5428, x5429;
  wire x5430, x5432, x5433, x5434, x5436, x5438, x5439, x5440;
  wire x5444, x5445, x5446, x5450, x5451, x5452, x5454, x5455;
  wire x5456, x5458, x5459, x5460, x5462, x5463, x5464, x5466;
  wire x5467, x5468, x5470, x5471, x5472, x5474, x5475, x5476;
  wire x5478, x5479, x5480, x5482, x5483, x5484, x5486, x5487;
  wire x5488, x5490, x5491, x5492, x5494, x5495, x5496, x5498;
  wire x5499, x5500, x5502, x5503, x5504, x5506, x5507, x5508;
  wire x5510, x5511, x5512, x5514, x5515, x5516, x5518, x5519;
  wire x5520, x5522, x5523, x5524, x5526, x5527, x5528, x5530;
  wire x5531, x5532, x5534, x5535, x5536, x5538, x5539, x5540;
  wire x5542, x5543, x5544, x5546, x5547, x5548, x5550, x5551;
  wire x5552, x5554, x5555, x5556, x5558, x5559, x5560, x5562;
  wire x5563, x5564, x5566, x5567, x5568, x5570, x5572, x5573;
  wire x5574, x5576, x5577, x5578, x5580, x5581, x5582, x5584;
  wire x5585, x5586, x5588, x5589, x5590, x5592, x5593, x5594;
  wire x5596, x5597, x5598, x5600, x5601, x5602, x5604, x5605;
  wire x5606, x5608, x5609, x5610, x5612, x5613, x5614, x5616;
  wire x5617, x5618, x5620, x5621, x5622, x5624, x5625, x5626;
  wire x5628, x5629, x5630, x5632, x5633, x5634, x5636, x5637;
  wire x5638, x5640, x5641, x5642, x5644, x5645, x5646, x5648;
  wire x5649, x5650, x5652, x5653, x5654, x5656, x5657, x5658;
  wire x5660, x5661, x5662, x5664, x5665, x5666, x5668, x5669;
  wire x5670, x5672, x5673, x5674, x5676, x5677, x5678, x5680;
  wire x5681, x5682, x5684, x5685, x5686, x5688, x5689, x5690;
  wire x5692, x5693, x5694, x5696, x5697, x5698, x5700, x5702;
  wire x5703, x5704, x5706, x5707, x5708, x5710, x5711, x5712;
  wire x5714, x5715, x5716, x5718, x5719, x5720, x5722, x5723;
  wire x5724, x5726, x5727, x5728, x5730, x5731, x5732, x5734;
  wire x5735, x5736, x5738, x5739, x5740, x5742, x5743, x5744;
  wire x5746, x5747, x5748, x5750, x5751, x5752, x5754, x5755;
  wire x5756, x5758, x5759, x5760, x5762, x5763, x5764, x5766;
  wire x5767, x5768, x5770, x5771, x5772, x5774, x5775, x5776;
  wire x5778, x5779, x5780, x5782, x5783, x5784, x5786, x5787;
  wire x5788, x5790, x5791, x5792, x5794, x5795, x5796, x5798;
  wire x5799, x5800, x5802, x5803, x5804, x5806, x5807, x5808;
  wire x5810, x5811, x5812, x5814, x5815, x5816, x5818, x5819;
  wire x5820, x5822, x5823, x5824, x5826, x5827, x5828, x5830;
  wire x5832, x5833, x5834, x5836, x5837, x5838, x5840, x5841;
  wire x5842, x5844, x5845, x5846, x5848, x5849, x5850, x5852;
  wire x5853, x5854, x5856, x5857, x5858, x5860, x5861, x5862;
  wire x5864, x5865, x5866, x5868, x5869, x5870, x5872, x5873;
  wire x5874, x5876, x5877, x5878, x5880, x5881, x5882, x5884;
  wire x5885, x5886, x5888, x5889, x5890, x5892, x5893, x5894;
  wire x5896, x5897, x5898, x5900, x5901, x5902, x5904, x5905;
  wire x5906, x5908, x5909, x5910, x5912, x5913, x5914, x5916;
  wire x5917, x5918, x5920, x5921, x5922, x5924, x5925, x5926;
  wire x5928, x5929, x5930, x5932, x5933, x5934, x5936, x5937;
  wire x5938, x5940, x5941, x5942, x5944, x5945, x5946, x5948;
  wire x5949, x5950, x5952, x5953, x5954, x5956, x5957, x5958;
  wire x5960, x5962, x5963, x5964, x5966, x5967, x5968, x5970;
  wire x5971, x5972, x5974, x5975, x5976, x5978, x5979, x5980;
  wire x5982, x5983, x5984, x5986, x5987, x5988, x5990, x5991;
  wire x5992, x5994, x5995, x5996, x5998, x5999, x6000, x6002;
  wire x6003, x6004, x6006, x6007, x6008, x6010, x6011, x6012;
  wire x6014, x6015, x6016, x6018, x6019, x6020, x6022, x6023;
  wire x6024, x6026, x6027, x6028, x6030, x6031, x6032, x6034;
  wire x6035, x6036, x6038, x6039, x6040, x6042, x6043, x6044;
  wire x6046, x6047, x6048, x6050, x6051, x6052, x6054, x6055;
  wire x6056, x6058, x6059, x6060, x6062, x6063, x6064, x6066;
  wire x6067, x6068, x6070, x6071, x6072, x6074, x6075, x6076;
  wire x6078, x6079, x6080, x6082, x6083, x6084, x6086, x6087;
  wire x6088, x6090, x6092, x6093, x6094, x6096, x6097, x6098;
  wire x6100, x6101, x6102, x6104, x6105, x6106, x6108, x6109;
  wire x6110, x6112, x6113, x6114, x6116, x6117, x6118, x6120;
  wire x6121, x6122, x6124, x6125, x6126, x6128, x6129, x6130;
  wire x6132, x6133, x6134, x6136, x6137, x6138, x6140, x6141;
  wire x6142, x6144, x6145, x6146, x6148, x6149, x6150, x6152;
  wire x6153, x6154, x6156, x6157, x6158, x6160, x6161, x6162;
  wire x6164, x6165, x6166, x6168, x6169, x6170, x6172, x6173;
  wire x6174, x6176, x6177, x6178, x6180, x6181, x6182, x6184;
  wire x6185, x6186, x6188, x6189, x6190, x6192, x6193, x6194;
  wire x6196, x6197, x6198, x6200, x6201, x6202, x6204, x6205;
  wire x6206, x6208, x6209, x6210, x6212, x6213, x6214, x6216;
  wire x6217, x6218, x6220, x6222, x6223, x6224, x6226, x6227;
  wire x6228, x6230, x6231, x6232, x6234, x6235, x6236, x6238;
  wire x6239, x6240, x6242, x6243, x6244, x6246, x6247, x6248;
  wire x6250, x6251, x6252, x6254, x6255, x6256, x6258, x6259;
  wire x6260, x6262, x6263, x6264, x6266, x6267, x6268, x6270;
  wire x6271, x6272, x6274, x6275, x6276, x6278, x6279, x6280;
  wire x6282, x6283, x6284, x6286, x6287, x6288, x6290, x6291;
  wire x6292, x6294, x6295, x6296, x6298, x6299, x6300, x6302;
  wire x6303, x6304, x6306, x6307, x6308, x6310, x6311, x6312;
  wire x6314, x6315, x6316, x6318, x6319, x6320, x6322, x6323;
  wire x6324, x6326, x6327, x6328, x6330, x6331, x6332, x6334;
  wire x6335, x6336, x6338, x6339, x6340, x6342, x6343, x6344;
  wire x6346, x6347, x6348, x6350, x6352, x6353, x6354, x6356;
  wire x6357, x6358, x6360, x6361, x6362, x6364, x6365, x6366;
  wire x6368, x6369, x6370, x6372, x6373, x6374, x6376, x6377;
  wire x6378, x6380, x6381, x6382, x6384, x6385, x6386, x6388;
  wire x6389, x6390, x6392, x6393, x6394, x6396, x6397, x6398;
  wire x6400, x6401, x6402, x6404, x6405, x6406, x6408, x6409;
  wire x6410, x6412, x6413, x6414, x6416, x6417, x6418, x6420;
  wire x6421, x6422, x6424, x6425, x6426, x6428, x6429, x6430;
  wire x6432, x6433, x6434, x6436, x6437, x6438, x6440, x6441;
  wire x6442, x6444, x6445, x6446, x6448, x6449, x6450, x6452;
  wire x6453, x6454, x6456, x6457, x6458, x6460, x6461, x6462;
  wire x6464, x6465, x6466, x6468, x6469, x6470, x6472, x6473;
  wire x6474, x6476, x6477, x6478, x6480, x6482, x6483, x6484;
  wire x6485, x6486, x6487, x6488, x6489, x6490, x6491, x6492;
  wire x6493, x6495, x6496, x6497, x6498, x6499, x6500, x6502;
  wire x6503, x6504, x6505, x6506, x6507, x6508, x6509, x6510;
  wire x6511, x6512, x6513, x6514, x6515, x6516, x6517, x6518;
  wire x6519, x6520, x6521, x6522, x6523, x6524, x6525, x6526;
  wire x6527, x6528, x6529, x6530, x6531, x6532, x6533, x6534;
  wire x6535, x6536, x6537, x6538, x6539, x6540, x6541, x6542;
  wire x6543, x6544, x6545, x6546, x6547, x6548, x6549, x6550;
  wire x6551, x6552, x6553, x6554, x6555, x6556, x6557, x6558;
  wire x6559, x6560, x6561, x6562, x6563, x6564, x6565, x6566;
  wire x6567, x6568, x6569, x6570, x6571, x6572, x6573, x6574;
  wire x6575, x6576, x6577, x6578, x6579, x6580, x6581, x6582;
  wire x6583, x6584, x6585, x6586, x6587, x6588, x6589, x6590;
  wire x6591, x6592, x6593, x6594, x6595, x6596, x6597, x6598;
  wire x6599, x6600, x6601, x6602, x6603, x6604, x6605, x6606;
  wire x6607, x6608, x6609, x6610, x6611, x6612, x6613, x6614;
  wire x6615, x6616, x6617, x6618, x6619, x6620, x6621, x6622;
  wire x6623, x6624, x6625, x6626, x6627, x6628, x6629, x6630;
  wire x6631, x6632, x6633, x6634, x6635, x6636, x6637, x6638;
  wire x6639, x6640, x6641, x6642, x6643, x6644, x6645, x6646;
  wire x6647, x6648, x6649, x6650, x6651, x6652, x6653, x6654;
  wire x6655, x6656, x6657, x6658, x6659, x6660, x6661, x6662;
  wire x6663, x6664, x6665, x6666, x6667, x6668, x6669, x6670;
  wire x6671, x6672, x6673, x6674, x6675, x6676, x6677, x6678;
  wire x6679, x6680, x6681, x6682, x6683, x6684, x6685, x6686;
  wire x6687, x6688, x6689, x6690, x6691, x6692, x6693, x6694;
  wire x6695, x6696, x6697, x6698, x6699, x6700, x6701, x6702;
  wire x6703, x6704, x6705, x6706, x6707, x6708, x6709, x6710;
  wire x6711, x6712, x6713, x6714, x6715, x6716, x6717, x6718;
  wire x6719, x6720, x6721, x6722, x6723, x6724, x6725, x6726;
  wire x6727, x6728, x6729, x6730, x6731, x6732, x6733, x6734;
  wire x6735, x6736, x6737, x6738, x6739, x6740, x6741, x6742;
  wire x6743, x6744, x6745, x6746, x6747, x6748, x6749, x6750;
  wire x6751, x6752, x6753, x6754, x6755, x6756, x6757, x6758;
  wire x6759, x6760, x6761, x6762, x6763, x6764, x6765, x6766;
  wire x6767, x6768, x6769, x6770, x6771, x6772, x6773, x6774;
  wire x6775, x6776, x6777, x6778, x6779, x6780, x6781, x6782;
  wire x6783, x6784, x6785, x6786, x6787, x6788, x6789, x6790;
  wire x6791, x6792, x6793, x6794, x6795, x6796, x6797, x6798;
  wire x6799, x6800, x6801, x6802, x6803, x6804, x6805, x6806;
  wire x6807, x6808, x6809, x6810, x6811, x6812, x6813, x6814;
  wire x6815, x6816, x6817, x6818, x6819, x6820, x6821, x6822;
  wire x6823, x6824, x6825, x6826, x6827, x6828, x6829, x6830;
  wire x6831, x6832, x6833, x6834, x6835, x6836, x6837, x6838;
  wire x6839, x6840, x6841, x6842, x6843, x6844, x6845, x6846;
  wire x6847, x6848, x6849, x6850, x6851, x6852, x6853, x6854;
  wire x6855, x6856, x6857, x6858, x6859, x6860, x6861, x6862;
  wire x6863, x6864, x6865, x6866, x6867, x6868, x6869, x6870;
  wire x6871, x6872, x6873, x6874, x6875, x6876, x6877, x6878;
  wire x6879, x6880, x6881, x6882, x6883, x6884, x6885, x6886;
  wire x6887, x6888, x6889, x6890, x6891, x6892, x6893, x6894;
  wire x6895, x6896, x6897, x6898, x6899, x6900, x6901, x6902;
  wire x6903, x6904, x6905, x6906, x6907, x6908, x6909, x6910;
  wire x6911, x6912, x6913, x6914, x6915, x6916, x6917, x6918;
  wire x6919, x6920, x6921, x6922, x6923, x6924, x6925, x6926;
  wire x6927, x6928, x6929, x6930, x6931, x6932, x6933, x6934;
  wire x6935, x6936, x6937, x6938, x6939, x6940, x6941, x6942;
  wire x6943, x6944, x6945, x6946, x6947, x6948, x6949, x6950;
  wire x6951, x6952, x6953, x6954, x6955, x6956, x6957, x6958;
  wire x6959, x6960, x6961, x6962, x6963, x6964, x6965, x6966;
  wire x6967, x6968, x6969, x6970, x6971, x6972, x6973, x6974;
  wire x6975, x6976, x6977, x6978, x6979, x6980, x6981, x6982;
  wire x6983, x6984, x6985, x6986, x6987, x6988, x6989, x6990;
  wire x6991, x6992, x6993, x6994, x6995, x6996, x6997, x6998;
  wire x6999, x7000, x7001, x7002, x7003, x7004, x7005, x7006;
  wire x7007, x7008, x7009, x7010, x7011, x7012, x7013, x7014;
  wire x7015, x7016, x7017, x7018, x7019, x7020, x7021, x7022;
  wire x7023, x7024, x7025, x7026, x7027, x7028, x7029, x7030;
  wire x7031, x7032, x7033, x7034, x7035, x7036, x7037, x7038;
  wire x7039, x7040, x7041, x7042, x7043, x7044, x7045, x7046;
  wire x7047, x7048, x7049, x7050, x7051, x7052, x7053, x7054;
  wire x7055, x7056, x7057, x7058, x7059, x7060, x7061, x7062;
  wire x7063, x7064, x7065, x7066, x7067, x7068, x7069, x7070;
  wire x7071, x7072, x7073, x7074, x7075, x7076, x7077, x7078;
  wire x7079, x7080, x7081, x7082, x7083, x7084, x7085, x7086;
  wire x7087, x7088, x7089, x7090, x7091, x7092, x7093, x7094;
  wire x7095, x7096, x7097, x7098, x7099, x7100, x7101, x7102;
  wire x7103, x7104, x7105, x7106, x7107, x7108, x7109, x7110;
  wire x7111, x7112, x7113, x7114, x7115, x7116, x7117, x7118;
  wire x7119, x7120, x7121, x7122, x7123, x7124, x7125, x7126;
  wire x7127, x7128, x7129, x7130, x7131, x7132, x7133, x7134;
  wire x7135, x7136, x7137, x7138, x7139, x7140, x7141, x7142;
  wire x7143, x7144, x7145, x7146, x7147, x7148, x7149, x7150;
  wire x7151, x7152, x7153, x7154, x7155, x7157, x7158, x7159;
  wire x7160, x7161, x7162, x7163, x7164, x7165, x7166, x7167;
  wire x7168, x7170, x7171, x7172, x7173, x7174, x7175, x7177;
  wire x7178, x7179, x7180, x7181, x7182, x7183, x7184, x7185;
  wire x7186, x7187, x7188, x7189, x7190, x7191, x7192, x7193;
  wire x7194, x7195, x7196, x7197, x7198, x7199, x7200, x7201;
  wire x7202, x7203, x7204, x7205, x7206, x7207, x7208, x7209;
  wire x7210, x7211, x7212, x7213, x7214, x7215, x7216, x7217;
  wire x7218, x7219, x7220, x7221, x7222, x7223, x7224, x7225;
  wire x7226, x7227, x7228, x7229, x7230, x7231, x7232, x7233;
  wire x7234, x7235, x7236, x7237, x7238, x7239, x7240, x7241;
  wire x7242, x7243, x7244, x7245, x7246, x7247, x7248, x7249;
  wire x7250, x7251, x7252, x7253, x7254, x7255, x7256, x7257;
  wire x7258, x7259, x7260, x7261, x7262, x7263, x7264, x7265;
  wire x7266, x7267, x7268, x7269, x7270, x7271, x7272, x7273;
  wire x7274, x7275, x7276, x7277, x7278, x7279, x7280, x7281;
  wire x7282, x7283, x7284, x7285, x7286, x7287, x7288, x7289;
  wire x7290, x7291, x7292, x7293, x7294, x7295, x7296, x7297;
  wire x7298, x7299, x7300, x7301, x7302, x7303, x7304, x7305;
  wire x7306, x7307, x7308, x7309, x7310, x7311, x7312, x7313;
  wire x7314, x7315, x7316, x7317, x7318, x7319, x7320, x7321;
  wire x7322, x7323, x7324, x7325, x7326, x7327, x7328, x7329;
  wire x7330, x7331, x7332, x7333, x7334, x7335, x7336, x7337;
  wire x7338, x7339, x7340, x7341, x7342, x7343, x7344, x7345;
  wire x7346, x7347, x7348, x7349, x7350, x7351, x7352, x7353;
  wire x7354, x7355, x7356, x7357, x7358, x7359, x7360, x7361;
  wire x7362, x7363, x7364, x7365, x7366, x7367, x7368, x7369;
  wire x7370, x7371, x7372, x7373, x7374, x7375, x7376, x7377;
  wire x7378, x7379, x7380, x7381, x7382, x7383, x7384, x7385;
  wire x7386, x7387, x7388, x7389, x7390, x7391, x7392, x7393;
  wire x7394, x7395, x7396, x7397, x7398, x7399, x7400, x7401;
  wire x7402, x7403, x7404, x7405, x7406, x7407, x7408, x7409;
  wire x7410, x7411, x7412, x7413, x7414, x7415, x7416, x7417;
  wire x7418, x7419, x7420, x7421, x7422, x7423, x7424, x7425;
  wire x7426, x7427, x7428, x7429, x7430, x7431, x7432, x7433;
  wire x7434, x7435, x7436, x7437, x7438, x7439, x7440, x7441;
  wire x7442, x7443, x7444, x7445, x7446, x7447, x7448, x7449;
  wire x7450, x7451, x7452, x7453, x7454, x7455, x7456, x7457;
  wire x7458, x7459, x7460, x7461, x7462, x7463, x7464, x7465;
  wire x7466, x7467, x7468, x7469, x7470, x7471, x7472, x7473;
  wire x7474, x7475, x7476, x7477, x7478, x7479, x7480, x7481;
  wire x7482, x7483, x7484, x7485, x7486, x7487, x7488, x7489;
  wire x7490, x7491, x7492, x7493, x7494, x7495, x7496, x7497;
  wire x7498, x7499, x7500, x7501, x7502, x7503, x7504, x7505;
  wire x7506, x7507, x7508, x7509, x7510, x7511, x7512, x7513;
  wire x7514, x7515, x7516, x7517, x7518, x7519, x7520, x7521;
  wire x7522, x7523, x7524, x7525, x7526, x7527, x7528, x7529;
  wire x7530, x7531, x7532, x7533, x7534, x7535, x7536, x7537;
  wire x7538, x7539, x7540, x7541, x7542, x7543, x7544, x7545;
  wire x7546, x7547, x7548, x7549, x7550, x7551, x7552, x7553;
  wire x7554, x7555, x7556, x7557, x7558, x7559, x7560, x7561;
  wire x7562, x7563, x7564, x7565, x7566, x7567, x7568, x7569;
  wire x7570, x7571, x7572, x7573, x7574, x7575, x7576, x7577;
  wire x7578, x7579, x7580, x7581, x7582, x7583, x7584, x7585;
  wire x7586, x7587, x7588, x7589, x7590, x7591, x7592, x7593;
  wire x7594, x7595, x7596, x7597, x7598, x7599, x7600, x7601;
  wire x7602, x7603, x7604, x7605, x7606, x7607, x7608, x7609;
  wire x7610, x7611, x7612, x7613, x7614, x7615, x7616, x7617;
  wire x7618, x7619, x7620, x7621, x7622, x7623, x7624, x7625;
  wire x7626, x7627, x7628, x7629, x7630, x7631, x7632, x7633;
  wire x7634, x7635, x7636, x7637, x7638, x7639, x7640, x7641;
  wire x7642, x7643, x7644, x7645, x7646, x7647, x7648, x7649;
  wire x7650, x7651, x7652, x7653, x7654, x7655, x7656, x7657;
  wire x7658, x7659, x7660, x7661, x7662, x7663, x7664, x7665;
  wire x7666, x7667, x7668, x7669, x7670, x7671, x7672, x7673;
  wire x7674, x7675, x7676, x7677, x7678, x7679, x7680, x7681;
  wire x7682, x7683, x7684, x7685, x7686, x7687, x7688, x7689;
  wire x7690, x7691, x7692, x7693, x7694, x7695, x7696, x7697;
  wire x7698, x7699, x7700, x7701, x7702, x7703, x7704, x7705;
  wire x7706, x7707, x7708, x7709, x7710, x7711, x7712, x7713;
  wire x7714, x7715, x7716, x7717, x7718, x7719, x7720, x7721;
  wire x7722, x7723, x7724, x7725, x7726, x7727, x7728, x7729;
  wire x7730, x7731, x7732, x7733, x7734, x7735, x7736, x7737;
  wire x7738, x7739, x7740, x7741, x7742, x7743, x7744, x7745;
  wire x7746, x7747, x7748, x7749, x7750, x7751, x7752, x7753;
  wire x7754, x7755, x7756, x7757, x7758, x7759, x7760, x7761;
  wire x7762, x7763, x7764, x7765, x7766, x7767, x7768, x7769;
  wire x7770, x7771, x7772, x7773, x7774, x7775, x7776, x7777;
  wire x7778, x7779, x7780, x7781, x7782, x7783, x7784, x7785;
  wire x7786, x7787, x7788, x7789, x7790, x7791, x7792, x7793;
  wire x7794, x7795, x7796, x7797, x7798, x7799, x7800, x7801;
  wire x7802, x7803, x7804, x7805, x7806, x7807, x7808, x7809;
  wire x7810, x7811, x7812, x7813, x7814, x7815, x7816, x7817;
  wire x7818, x7819, x7820, x7821, x7822, x7823, x7824, x7825;
  wire x7826, x7827, x7828, x7829, x7830, x7831, x7832, x7833;
  wire x7834, x7835, x7836, x7837, x7838, x7839, x7840, x7841;
  wire x7842, x7843, x7844, x7845, x7846, x7847, x7848, x7849;
  wire x7850, x7851, x7852, x7853, x7854, x7855, x7856, x7857;
  wire x7858, x7859, x7860, x7861, x7862, x7863, x7864, x7865;
  wire x7866, x7867, x7868, x7869, x7870, x7871, x7872, x7873;
  wire x7874, x7875, x7876, x7877, x7878, x7879, x7880, x7881;
  wire x7882, x7883, x7884, x7885, x7886, x7887, x7888, x7889;
  wire x7890, x7891, x7892, x7893, x7894, x7895, x7896, x7897;
  wire x7898, x7899, x7900, x7901, x7902, x7903, x7904, x7905;
  wire x7906, x7907, x7908, x7909, x7910, x7911, x7912, x7913;
  wire x7914, x7915, x7916, x7917, x7918, x7919, x7920, x7921;
  wire x7922, x7923, x7924, x7925, x7926, x7927, x7928, x7929;
  wire x7930, x7931, x7932, x7933, x7934, x7935, x7936, x7937;
  wire x7938, x7939, x7940, x7941, x7942, x7943, x7944, x7945;
  wire x7946, x7947, x7948, x7949, x7950, x7951, x7952, x7953;
  wire x7954, x7955, x7956, x7957, x7958, x7959, x7960, x7961;
  wire x7962, x7963, x7964, x7965, x7966, x7967, x7968, x7969;
  wire x7970, x7971, x7972, x7973, x7974, x7975, x7976, x7977;
  wire x7978, x7979, x7980, x7981, x7982, x7983, x7984, x7985;
  wire x7986, x7987, x7988, x7989, x7990, x7991, x7992, x7993;
  wire x7994, x7995, x7996, x7997, x7998, x7999, x8000, x8001;
  wire x8002, x8003, x8004, x8005, x8006, x8007, x8008, x8009;
  wire x8010, x8011, x8012, x8013, x8014, x8015, x8016, x8017;
  wire x8018, x8019, x8020, x8021, x8022, x8023, x8024, x8025;
  wire x8026, x8027, x8028, x8029, x8030, x8031, x8032, x8033;
  wire x8034, x8035, x8036, x8037, x8038, x8039, x8040, x8041;
  wire x8042, x8043, x8044, x8045, x8046, x8047, x8048, x8049;
  wire x8050, x8051, x8052, x8053, x8054, x8055, x8056, x8057;
  wire x8058, x8059, x8060, x8061, x8062, x8063, x8064, x8065;
  wire x8066, x8067, x8068, x8069, x8070, x8071, x8072, x8073;
  wire x8074, x8075, x8076, x8077, x8078, x8079, x8080, x8081;
  wire x8082, x8083, x8084, x8085, x8086, x8087, x8088, x8089;
  wire x8090, x8091, x8092, x8093, x8094, x8095, x8096, x8097;
  wire x8098, x8099, x8100, x8101, x8102, x8103, x8104, x8105;
  wire x8106, x8107, x8108, x8109, x8110, x8111, x8112, x8113;
  wire x8114, x8115, x8116, x8117, x8118, x8119, x8120, x8121;
  wire x8122, x8123, x8124, x8125, x8126, x8127, x8128, x8129;
  wire x8130, x8131, x8132, x8133, x8134, x8135, x8136, x8137;
  wire x8138, x8139, x8140, x8141, x8142, x8143, x8144, x8145;
  wire x8146, x8147, x8148, x8149, x8150, x8151, x8152, x8153;
  wire x8154, x8155, x8156, x8157, x8158, x8159, x8160, x8161;
  wire x8162, x8163, x8164, x8165, x8166, x8167, x8168, x8169;
  wire x8170, x8171, x8172, x8173, x8174, x8175, x8176, x8177;
  wire x8178, x8179, x8180, x8181, x8182, x8183, x8184, x8185;
  wire x8186, x8187, x8188, x8189, x8190, x8191, x8192, x8193;
  wire x8194, x8195, x8196, x8197, x8198, x8199, x8200, x8201;
  wire x8202, x8203, x8204, x8205, x8206, x8207, x8208, x8209;
  wire x8210, x8211, x8212, x8213, x8214, x8215, x8216, x8217;
  wire x8218, x8219, x8220, x8221, x8222, x8223, x8224, x8225;
  wire x8226, x8227, x8228, x8229, x8230, x8231, x8232, x8233;
  wire x8234, x8235, x8236, x8237, x8238, x8239, x8240, x8241;
  wire x8242, x8243, x8244, x8245, x8246, x8247, x8248, x8249;
  wire x8250, x8251, x8252, x8253, x8254, x8255, x8256, x8257;
  wire x8258, x8259, x8260, x8261, x8262, x8263, x8264, x8265;
  wire x8266, x8267, x8268, x8269, x8270, x8271, x8272, x8273;
  wire x8274, x8275, x8276, x8277, x8278, x8279, x8280, x8281;
  wire x8282, x8283, x8284, x8285, x8286, x8287, x8288, x8289;
  wire x8290, x8291, x8292, x8293, x8294, x8295, x8296, x8297;
  wire x8298, x8299, x8300, x8301, x8302, x8303, x8304, x8305;
  wire x8306, x8307, x8308, x8309, x8310, x8311, x8312, x8313;
  wire x8314, x8315, x8316, x8317, x8318, x8319, x8320, x8321;
  wire x8322, x8323, x8324, x8325, x8326, x8327, x8328, x8329;
  wire x8330, x8331, x8332, x8333, x8334, x8335, x8336, x8337;
  wire x8338, x8339, x8340, x8341, x8342, x8343, x8344, x8345;
  wire x8346, x8347, x8348, x8349, x8350, x8351, x8352, x8353;
  wire x8354, x8355, x8356, x8357, x8358, x8359, x8360, x8361;
  wire x8362, x8363, x8364, x8365, x8366, x8367, x8368, x8369;
  wire x8370, x8371, x8372, x8373, x8374, x8375, x8376, x8377;
  wire x8378, x8379, x8380, x8381, x8382, x8383, x8384, x8385;
  wire x8386, x8387, x8388, x8389, x8390, x8391, x8392, x8393;
  wire x8394, x8395, x8396, x8397, x8398, x8399, x8400, x8401;
  wire x8402, x8403, x8404, x8405, x8406, x8407, x8408, x8409;
  wire x8410, x8411, x8412, x8413, x8414, x8415, x8416, x8417;
  wire x8418, x8419, x8420, x8421, x8422, x8423, x8424, x8425;
  wire x8426, x8427, x8428, x8429, x8430, x8431, x8432, x8433;
  wire x8434, x8435, x8436, x8437, x8438, x8439, x8440, x8441;
  wire x8442, x8443, x8444, x8445, x8446, x8447, x8448, x8449;
  wire x8450, x8451, x8452, x8453, x8454, x8455, x8456, x8457;
  wire x8458, x8459, x8460, x8461, x8462, x8463, x8464, x8465;
  wire x8466, x8467, x8468, x8469, x8470, x8471, x8472, x8473;
  wire x8474, x8475, x8476, x8477, x8478, x8479, x8480, x8481;
  wire x8482, x8483, x8484, x8485, x8486, x8487, x8488, x8489;
  wire x8490, x8491, x8492, x8493, x8494, x8495, x8496, x8497;
  wire x8498, x8499, x8500, x8501, x8502, x8503, x8504, x8505;
  wire x8506, x8507, x8508, x8509, x8510, x8511, x8512, x8513;
  wire x8514, x8515, x8516, x8517, x8518, x8519, x8520, x8521;
  wire x8522, x8523, x8524, x8525, x8526, x8527, x8528, x8529;
  wire x8530, x8531, x8532, x8533, x8534, x8535, x8536, x8537;
  wire x8538, x8539, x8540, x8541, x8542, x8543, x8544, x8545;
  wire x8546, x8547, x8548, x8549, x8550, x8551, x8552, x8553;
  wire x8554, x8555, x8556, x8557, x8558, x8559, x8560, x8561;
  wire x8562, x8563, x8564, x8565, x8566, x8567, x8568, x8569;
  wire x8570, x8571, x8572, x8573, x8574, x8575, x8576, x8577;
  wire x8578, x8579, x8580, x8581, x8582, x8583, x8584, x8585;
  wire x8586, x8587, x8588, x8589, x8590, x8591, x8592, x8593;
  wire x8594, x8595, x8596, x8597, x8598, x8599, x8600, x8601;
  wire x8602, x8603, x8604, x8605, x8606, x8607, x8608, x8609;
  wire x8610, x8611, x8612, x8613, x8614, x8615, x8616, x8617;
  wire x8618, x8619, x8620, x8621, x8622, x8623, x8624, x8625;
  wire x8626, x8627, x8628, x8629, x8630, x8631, x8632, x8633;
  wire x8634, x8635, x8636, x8637, x8638, x8639, x8640, x8641;
  wire x8642, x8643, x8644, x8645, x8646, x8647, x8648, x8649;
  wire x8650, x8651, x8652, x8653, x8654, x8655, x8656, x8657;
  wire x8658, x8659, x8660, x8661, x8662, x8663, x8664, x8665;
  wire x8666, x8667, x8668, x8669, x8670, x8671, x8672, x8673;
  wire x8674, x8675, x8676, x8677, x8678, x8679, x8680, x8681;
  wire x8682, x8683, x8684, x8685, x8686, x8687, x8688, x8689;
  wire x8690, x8691, x8692, x8693, x8694, x8695, x8696, x8697;
  wire x8698, x8699, x8700, x8701, x8702, x8703, x8704, x8705;
  wire x8706, x8707, x8708, x8709, x8710, x8711, x8712, x8713;
  wire x8714, x8715, x8716, x8717, x8718, x8719, x8720, x8721;
  wire x8722, x8723, x8724, x8725, x8726, x8727, x8728, x8729;
  wire x8730, x8731, x8732, x8733, x8734, x8735, x8736, x8737;
  wire x8738, x8739, x8740, x8741, x8742, x8743, x8744, x8745;
  wire x8746, x8747, x8748, x8749, x8750, x8751, x8752, x8753;
  wire x8754, x8755, x8756, x8757, x8758, x8759, x8760, x8761;
  wire x8762, x8763, x8764, x8765, x8766, x8767, x8768, x8769;
  wire x8770, x8771, x8772, x8773, x8774, x8775, x8776, x8777;
  wire x8778, x8779, x8780, x8781, x8782, x8783, x8784, x8785;
  wire x8786, x8787, x8788, x8789, x8790, x8791, x8792, x8793;
  wire x8794, x8795, x8796, x8797, x8798, x8799, x8800, x8801;
  wire x8802, x8803, x8804, x8805, x8806, x8807, x8808, x8809;
  wire x8810, x8811, x8812, x8813, x8814, x8815, x8816, x8817;
  wire x8818, x8819, x8820, x8821, x8822, x8823, x8824, x8825;
  wire x8826, x8827, x8828, x8829, x8830, x8831, x8832, x8833;
  wire x8834, x8835, x8836, x8837, x8838, x8839, x8840, x8841;
  wire x8842, x8843, x8844, x8845, x8846, x8847, x8848, x8849;
  wire x8850, x8851, x8852, x8853, x8854, x8855, x8856, x8857;
  wire x8858, x8859, x8860, x8861, x8862, x8863, x8864, x8865;
  wire x8866, x8867, x8868, x8869, x8870, x8871, x8872, x8873;
  wire x8874, x8875, x8876, x8877, x8878, x8879, x8880, x8881;
  wire x8882, x8883, x8884, x8885, x8886, x8887, x8888, x8889;
  wire x8890, x8891, x8892, x8893, x8894, x8895, x8896, x8897;
  wire x8898, x8899, x8900, x8901, x8902, x8903, x8904, x8905;
  wire x8906, x8907, x8908, x8909, x8910, x8911, x8912, x8913;
  wire x8914, x8915, x8916, x8917, x8918, x8919, x8920, x8921;
  wire x8922, x8923, x8924, x8925, x8926, x8927, x8928, x8929;
  wire x8930, x8931, x8932, x8933, x8934, x8935, x8936, x8937;
  wire x8938, x8939, x8940, x8941, x8942, x8943, x8944, x8945;
  wire x8946, x8947, x8948, x8949, x8950, x8951, x8952, x8953;
  wire x8954, x8955, x8956, x8957, x8958, x8959, x8960, x8961;
  wire x8962, x8963, x8964, x8965, x8966, x8967, x8968, x8969;
  wire x8970, x8971, x8972, x8973, x8974, x8975, x8976, x8977;
  wire x8978, x8979, x8980, x8981, x8982, x8983, x8984, x8985;
  wire x8986, x8987, x8988, x8989, x8990, x8991, x8992, x8993;
  wire x8994, x8995, x8996, x8997, x8998, x8999, x9000, x9001;
  wire x9002, x9003, x9004, x9005, x9006, x9007, x9008, x9009;
  wire x9010, x9011, x9012, x9013, x9014, x9015, x9016, x9017;
  wire x9018, x9019, x9020, x9021, x9022, x9023, x9024, x9025;
  wire x9026, x9027, x9028, x9029, x9030, x9031, x9032, x9033;
  wire x9034, x9035, x9036, x9037, x9038, x9039, x9040, x9041;
  wire x9042, x9043, x9044, x9045, x9046, x9047, x9048, x9049;
  wire x9050, x9051, x9052, x9053, x9054, x9055, x9056, x9057;
  wire x9058, x9059, x9060, x9061, x9062, x9063, x9064, x9065;
  wire x9066, x9067, x9068, x9069, x9070, x9071, x9072, x9073;
  wire x9074, x9075, x9076, x9077, x9078, x9079, x9080, x9081;
  wire x9082, x9083, x9084, x9085, x9086, x9087, x9088, x9089;
  wire x9090, x9091, x9092, x9093, x9094, x9095, x9096, x9097;
  wire x9098, x9099, x9100, x9101, x9102, x9103, x9104, x9105;
  wire x9106, x9107, x9108, x9109, x9110, x9111, x9112, x9113;
  wire x9114, x9115, x9116, x9117, x9118, x9119, x9120, x9121;
  wire x9122, x9123, x9124, x9125, x9126, x9127, x9128, x9129;
  wire x9130, x9131, x9132, x9133, x9134, x9135, x9136, x9137;
  wire x9138, x9139, x9140, x9141, x9142, x9143, x9144, x9145;
  wire x9146, x9147, x9148, x9149, x9150, x9151, x9152, x9153;
  wire x9154, x9155, x9156, x9157, x9158, x9159, x9160, x9161;
  wire x9162, x9163, x9164, x9165, x9166, x9167, x9168, x9169;
  wire x9170, x9171, x9172, x9173, x9174, x9175, x9176, x9177;
  wire x9178, x9179, x9180, x9181, x9182, x9183, x9184, x9185;
  wire x9186, x9187, x9188, x9189, x9190, x9191, x9192, x9193;
  wire x9194, x9195, x9196, x9197, x9198, x9199, x9200, x9201;
  wire x9202, x9203, x9204, x9205, x9206, x9207, x9208, x9209;
  wire x9210, x9211, x9212, x9213, x9214, x9215, x9216, x9217;
  wire x9218, x9219, x9220, x9221, x9222, x9223, x9224, x9225;
  wire x9226, x9227, x9228, x9229, x9230, x9231, x9232, x9233;
  wire x9234, x9235, x9236, x9237, x9238, x9239, x9240, x9241;
  wire x9242, x9243, x9244, x9245, x9246, x9247, x9248, x9249;
  wire x9250, x9251, x9252, x9253, x9254, x9255, x9256, x9257;
  wire x9258, x9259, x9260, x9261, x9262, x9263, x9264, x9265;
  wire x9266, x9267, x9268, x9269, x9270, x9271, x9272, x9273;
  wire x9274, x9275, x9276, x9277, x9278, x9279, x9280, x9281;
  wire x9282, x9283, x9284, x9285, x9286, x9287, x9288, x9289;
  wire x9290, x9291, x9292, x9293, x9294, x9295, x9296, x9297;
  wire x9298, x9299, x9300, x9301, x9302, x9303, x9304, x9305;
  wire x9306, x9307, x9308, x9309, x9310, x9311, x9312, x9313;
  wire x9314, x9315, x9316, x9317, x9318, x9319, x9320, x9321;
  wire x9322, x9323, x9324, x9325, x9326, x9327, x9328, x9329;
  wire x9330, x9331, x9332, x9333, x9334, x9335, x9336, x9337;
  wire x9338, x9339, x9340, x9341, x9342, x9343, x9344, x9345;
  wire x9346, x9347, x9348, x9349, x9350, x9351, x9352, x9353;
  wire x9354, x9355, x9356, x9357, x9358, x9359, x9360, x9361;
  wire x9362, x9363, x9364, x9365, x9366, x9367, x9368, x9369;
  wire x9370, x9371, x9372, x9373, x9374, x9375, x9376, x9377;
  wire x9378, x9379, x9380, x9381, x9382, x9383, x9384, x9385;
  wire x9386, x9387, x9388, x9389, x9390, x9391, x9392, x9393;
  wire x9394, x9395, x9396, x9397, x9398, x9399, x9400, x9401;
  wire x9402, x9403, x9404, x9405, x9406, x9407, x9408, x9409;
  wire x9410, x9411, x9412, x9413, x9414, x9415, x9416, x9417;
  wire x9418, x9419, x9420, x9421, x9422, x9423, x9424, x9425;
  wire x9426, x9427, x9428, x9429, x9430, x9431, x9432, x9433;
  wire x9434, x9435, x9436, x9437, x9438, x9439, x9440, x9441;
  wire x9442, x9443, x9444, x9445, x9446, x9447, x9448, x9449;
  wire x9450, x9451, x9452, x9453, x9454, x9455, x9456, x9457;
  wire x9458, x9459, x9460, x9461, x9462, x9463, x9464, x9465;
  wire x9466, x9467, x9468, x9469, x9470, x9471, x9472, x9473;
  wire x9474, x9475, x9476, x9477, x9478, x9479, x9480, x9481;
  wire x9482, x9483, x9484, x9485, x9486, x9487, x9488, x9489;
  wire x9490, x9491, x9492, x9493, x9494, x9495, x9496, x9497;
  wire x9498, x9499, x9500, x9501, x9502, x9503, x9504, x9505;
  wire x9506, x9507, x9508, x9509, x9510, x9511, x9512, x9513;
  wire x9514, x9515, x9516, x9517, x9518, x9519, x9520, x9521;
  wire x9522, x9523, x9524, x9525, x9526, x9527, x9528, x9529;
  wire x9530, x9531, x9532, x9533, x9534, x9535, x9536, x9537;
  wire x9538, x9539, x9540, x9541, x9542, x9543, x9544, x9545;
  wire x9546, x9547, x9548, x9549, x9550, x9551, x9552, x9553;
  wire x9554, x9555, x9556, x9557, x9558, x9559, x9560, x9561;
  wire x9562, x9563, x9564, x9565, x9566, x9567, x9568, x9569;
  wire x9570, x9571, x9572, x9573, x9574, x9575, x9576, x9577;
  wire x9578, x9579, x9580, x9581, x9582, x9583, x9584, x9585;
  wire x9586, x9587, x9588, x9589, x9590, x9591, x9592, x9593;
  wire x9594, x9595, x9596, x9597, x9598, x9599, x9600, x9601;
  wire x9602, x9603, x9604, x9605, x9606, x9607, x9608, x9609;
  wire x9610, x9611, x9612, x9613, x9614, x9615, x9616, x9617;
  wire x9618, x9619, x9620, x9621, x9622, x9623, x9624, x9625;
  wire x9626, x9627, x9628, x9629, x9630, x9631, x9632, x9633;
  wire x9634, x9635, x9636, x9637, x9638, x9639, x9640, x9641;
  wire x9642, x9643, x9644, x9645, x9646, x9647, x9648, x9649;
  wire x9650, x9651, x9652, x9653, x9654, x9655, x9656, x9657;
  wire x9658, x9659, x9660, x9661, x9662, x9663, x9664, x9665;
  wire x9666, x9667, x9668, x9669, x9670, x9671, x9672, x9673;
  wire x9674, x9675, x9676, x9677, x9678, x9679, x9680, x9681;
  wire x9682, x9683, x9684, x9685, x9686, x9687, x9688, x9689;
  wire x9690, x9691, x9692, x9693, x9694, x9695, x9696, x9697;
  wire x9698, x9699, x9700, x9701, x9702, x9703, x9704, x9705;
  wire x9706, x9707, x9708, x9709, x9710, x9711, x9712, x9713;
  wire x9714, x9715, x9716, x9717, x9718, x9719, x9720, x9721;
  wire x9722, x9723, x9724, x9725, x9726, x9727, x9728, x9729;
  wire x9730, x9731, x9732, x9733, x9734, x9735, x9736, x9737;
  wire x9738, x9739, x9740, x9741, x9742, x9743, x9744, x9745;
  wire x9746, x9747, x9748, x9749, x9750, x9751, x9752, x9753;
  wire x9754, x9755, x9756, x9757, x9758, x9759, x9760, x9761;
  wire x9762, x9763, x9764, x9765, x9766, x9767, x9768, x9769;
  wire x9770, x9771, x9772, x9773, x9774, x9775, x9776, x9777;
  wire x9778, x9779, x9780, x9781, x9782, x9783, x9784, x9785;
  wire x9786, x9787, x9788, x9789, x9790, x9791, x9792, x9793;
  wire x9794, x9795, x9796, x9797, x9798, x9799, x9800, x9801;
  wire x9802, x9803, x9804, x9805, x9806, x9807, x9808, x9809;
  wire x9810, x9811, x9812, x9813, x9814, x9815, x9816, x9817;
  wire x9818, x9819, x9820, x9821, x9822, x9823, x9824, x9825;
  wire x9826, x9827, x9828, x9829, x9830, x9831, x9832, x9833;
  wire x9834, x9835, x9836, x9837, x9838, x9839, x9840, x9841;
  wire x9842, x9843, x9844, x9845, x9846, x9847, x9848, x9849;
  wire x9850, x9851, x9852, x9853, x9854, x9855, x9856, x9857;
  wire x9858, x9859, x9860, x9861, x9862, x9863, x9864, x9865;
  wire x9866, x9867, x9868, x9869, x9870, x9871, x9872, x9873;
  wire x9874, x9875, x9876, x9877, x9878, x9879, x9880, x9881;
  wire x9882, x9883, x9884, x9885, x9886, x9887, x9888, x9889;
  wire x9890, x9891, x9892, x9893, x9894, x9895, x9896, x9897;
  wire x9898, x9899, x9900, x9901, x9902, x9903, x9904, x9905;
  wire x9906, x9907, x9908, x9909, x9910, x9911, x9912, x9913;
  wire x9914, x9915, x9916, x9917, x9918, x9919, x9920, x9921;
  wire x9922, x9923, x9924, x9925, x9926, x9927, x9928, x9929;
  wire x9930, x9931, x9932, x9933, x9934, x9935, x9936, x9937;
  wire x9938, x9939, x9940, x9941, x9942, x9943, x9944, x9945;
  wire x9946, x9947, x9948, x9949, x9950, x9951, x9952, x9953;
  wire x9954, x9955, x9956, x9957, x9958, x9959, x9960, x9961;
  wire x9962, x9963, x9964, x9965, x9966, x9967, x9968, x9969;
  wire x9970, x9971, x9972, x9973, x9974, x9975, x9976, x9977;
  wire x9978, x9979, x9980, x9981, x9982, x9983, x9984, x9985;
  wire x9986, x9987, x9988, x9989, x9990, x9991, x9992, x9993;
  wire x9994, x9995, x9996, x9997, x9998, x9999, x10000, x10001;
  wire x10002, x10003, x10004, x10005, x10006, x10007, x10008, x10009;
  wire x10010, x10011, x10012, x10013, x10014, x10015, x10016, x10017;
  wire x10018, x10019, x10020, x10021, x10022, x10023, x10024, x10025;
  wire x10026, x10027, x10028, x10029, x10030, x10031, x10032, x10033;
  wire x10034, x10035, x10036, x10037, x10038, x10039, x10040, x10041;
  wire x10042, x10043, x10044, x10045, x10046, x10047, x10048, x10049;
  wire x10050, x10051, x10052, x10053, x10054, x10055, x10056, x10057;
  wire x10058, x10059, x10060, x10061, x10062, x10063, x10064, x10065;
  wire x10066, x10067, x10068, x10069, x10070, x10071, x10072, x10073;
  wire x10074, x10075, x10076, x10077, x10078, x10079, x10080, x10081;
  wire x10082, x10083, x10084, x10085, x10086, x10087, x10088, x10089;
  wire x10090, x10091, x10092, x10093, x10094, x10095, x10096, x10097;
  wire x10098, x10099, x10100, x10101, x10102, x10103, x10104, x10105;
  wire x10106, x10107, x10108, x10109, x10110, x10111, x10112, x10113;
  wire x10114, x10115, x10116, x10117, x10118, x10119, x10120, x10121;
  wire x10122, x10123, x10124, x10125, x10126, x10127, x10128, x10129;
  wire x10130, x10131, x10132, x10133, x10134, x10135, x10136, x10137;
  wire x10138, x10139, x10140, x10141, x10142, x10143, x10144, x10145;
  wire x10146, x10147, x10148, x10149, x10150, x10151, x10152, x10153;
  wire x10154, x10155, x10156, x10157, x10158, x10159, x10160, x10161;
  wire x10162, x10163, x10164, x10165, x10166, x10167, x10168, x10169;
  wire x10170, x10171, x10172, x10173, x10174, x10175, x10176, x10177;
  wire x10178, x10179, x10180, x10181, x10182, x10183, x10184, x10185;
  wire x10186, x10187, x10188, x10189, x10190, x10191, x10192, x10193;
  wire x10194, x10195, x10196, x10197, x10198, x10199, x10200, x10201;
  wire x10202, x10203, x10204, x10205, x10206, x10207, x10208, x10209;
  wire x10210, x10211, x10212, x10213, x10214, x10215, x10216, x10217;
  wire x10218, x10219, x10220, x10221, x10222, x10223, x10224, x10225;
  wire x10226, x10227, x10228, x10229, x10230, x10231, x10232, x10233;
  wire x10234, x10235, x10236, x10237, x10238, x10239, x10240, x10241;
  wire x10242, x10243, x10244, x10245, x10246, x10247, x10248, x10249;
  wire x10250, x10251, x10252, x10253, x10254, x10255, x10256, x10257;
  wire x10258, x10259, x10260, x10261, x10262, x10263, x10264, x10265;
  wire x10266, x10267, x10268, x10269, x10270, x10271, x10272, x10273;
  wire x10274, x10275, x10276, x10277, x10278, x10279, x10280, x10281;
  wire x10282, x10283, x10284, x10285, x10286, x10287, x10288, x10289;
  wire x10290, x10291, x10292, x10293, x10294, x10295, x10296, x10297;
  wire x10298, x10299, x10300, x10301, x10302, x10303, x10304, x10305;
  wire x10306, x10307, x10308, x10309, x10310, x10311, x10312, x10313;
  wire x10314, x10315, x10316, x10317, x10318, x10319, x10320, x10321;
  wire x10322, x10323, x10324, x10325, x10326, x10327, x10328, x10329;
  wire x10330, x10331, x10332, x10333, x10334, x10335, x10336, x10337;
  wire x10338, x10339, x10340, x10341, x10342, x10343, x10344, x10345;
  wire x10346, x10347, x10348, x10349, x10350, x10351, x10352, x10353;
  wire x10354, x10355, x10356, x10357, x10358, x10359, x10360, x10361;
  wire x10362, x10363, x10364, x10365, x10366, x10367, x10368, x10369;
  wire x10370, x10371, x10372, x10373, x10374, x10375, x10376, x10377;
  wire x10378, x10379, x10380, x10381, x10382, x10383, x10384, x10385;
  wire x10386, x10387, x10388, x10389, x10390, x10391, x10392, x10393;
  wire x10394, x10395, x10396, x10397, x10398, x10399, x10400, x10401;
  wire x10402, x10403, x10404, x10405, x10406, x10407, x10408, x10409;
  wire x10410, x10411, x10412, x10413, x10414, x10415, x10416, x10417;
  wire x10418, x10419, x10420, x10421, x10422, x10423, x10424, x10425;
  wire x10426, x10427, x10428, x10429, x10430, x10431, x10432, x10433;
  wire x10434, x10435, x10436, x10437, x10438, x10439, x10440, x10441;
  wire x10442, x10443, x10444, x10445, x10446, x10447, x10448, x10449;
  wire x10450, x10451, x10452, x10453, x10454, x10455, x10456, x10457;
  wire x10458, x10459, x10460, x10461, x10462, x10463, x10464, x10465;
  wire x10466, x10467, x10468, x10469, x10470, x10471, x10472, x10473;
  wire x10474, x10475, x10476, x10477, x10478, x10479, x10480, x10481;
  wire x10482, x10483, x10484, x10485, x10486, x10487, x10488, x10489;
  wire x10490, x10491, x10492, x10493, x10494, x10495, x10496, x10497;
  wire x10498, x10499, x10500, x10501, x10502, x10503, x10504, x10505;
  wire x10506, x10507, x10508, x10509, x10510, x10511, x10512, x10513;
  wire x10514, x10515, x10516, x10517, x10518, x10519, x10520, x10521;
  wire x10522, x10523, x10524, x10525, x10526, x10527, x10528, x10529;
  wire x10530, x10531, x10532, x10533, x10534, x10535, x10536, x10537;
  wire x10538, x10539, x10540, x10541, x10542, x10543, x10544, x10545;
  wire x10546, x10547, x10548, x10549, x10550, x10551, x10552, x10553;
  wire x10554, x10555, x10556, x10557, x10558, x10559, x10560, x10561;
  wire x10562, x10563, x10564, x10565, x10566, x10567, x10568, x10569;
  wire x10570, x10571, x10572, x10573, x10574, x10575, x10576, x10577;
  wire x10578, x10579, x10580, x10581, x10582, x10583, x10584, x10585;
  wire x10586, x10587, x10588, x10589, x10590, x10591, x10592, x10593;
  wire x10594, x10595, x10596, x10597, x10598, x10599, x10600, x10601;
  wire x10602, x10603, x10604, x10605, x10606, x10607, x10608, x10609;
  wire x10610, x10611, x10612, x10613, x10614, x10615, x10616, x10617;
  wire x10618, x10619, x10620, x10621, x10622, x10623, x10624, x10625;
  wire x10626, x10627, x10628, x10629, x10630, x10631, x10632, x10633;
  wire x10634, x10635, x10636, x10637, x10638, x10639, x10640, x10641;
  wire x10642, x10643, x10644, x10645, x10646, x10647, x10648, x10649;
  wire x10650, x10651, x10652, x10653, x10654, x10655, x10656, x10657;
  wire x10658, x10659, x10660, x10661, x10662, x10663, x10664, x10665;
  wire x10666, x10667, x10668, x10669, x10670, x10671, x10672, x10673;
  wire x10674, x10675, x10676, x10677, x10678, x10679, x10680, x10681;
  wire x10682, x10683, x10684, x10685, x10686, x10687, x10688, x10689;
  wire x10690, x10691, x10692, x10693, x10694, x10695, x10696, x10697;
  wire x10698, x10699, x10700, x10701, x10702, x10703, x10704, x10705;
  wire x10706, x10707, x10708, x10709, x10710, x10711, x10712, x10713;
  wire x10714, x10715, x10716, x10717, x10718, x10719, x10720, x10721;
  wire x10722, x10723, x10724, x10725, x10726, x10727, x10728, x10729;
  wire x10730, x10731, x10732, x10733, x10734, x10735, x10736, x10737;
  wire x10738, x10739, x10740, x10741, x10742, x10743, x10744, x10745;
  wire x10746, x10747, x10748, x10749, x10750, x10751, x10752, x10753;
  wire x10754, x10755, x10756, x10757, x10758, x10759, x10760, x10761;
  wire x10762, x10763, x10764, x10765, x10766, x10767, x10768, x10769;
  wire x10770, x10771, x10772, x10773, x10774, x10775, x10776, x10777;
  wire x10778, x10779, x10780, x10781, x10782, x10783, x10784, x10785;
  wire x10786, x10787, x10788, x10789, x10790, x10791, x10792, x10793;
  wire x10794, x10795, x10796, x10797, x10798, x10799, x10800, x10801;
  wire x10802, x10803, x10804, x10805, x10806, x10807, x10808, x10809;
  wire x10810, x10811, x10812, x10813, x10814, x10815, x10816, x10817;
  wire x10818, x10819, x10820, x10821, x10822, x10823, x10824, x10825;
  wire x10826, x10827, x10828, x10829, x10830, x10831, x10832, x10833;
  wire x10834, x10835, x10836, x10837, x10838, x10839, x10840, x10841;
  wire x10842, x10843, x10844, x10845, x10846, x10847, x10848, x10849;
  wire x10850, x10851, x10852, x10853, x10854, x10855, x10856, x10857;
  wire x10858, x10859, x10860, x10861, x10862, x10863, x10864, x10865;
  wire x10866, x10867, x10868, x10869, x10870, x10871, x10872, x10873;
  wire x10874, x10875, x10876, x10877, x10878, x10879, x10880, x10881;
  wire x10882, x10883, x10884, x10885, x10886, x10887, x10888, x10889;
  wire x10890, x10891, x10892, x10893, x10894, x10895, x10896, x10897;
  wire x10898, x10899, x10900, x10901, x10902, x10903, x10904, x10905;
  wire x10906, x10907, x10908, x10909, x10910, x10911, x10912, x10913;
  wire x10914, x10915, x10916, x10917, x10918, x10919, x10920, x10921;
  wire x10922, x10923, x10924, x10925, x10926, x10927, x10928, x10929;
  wire x10930, x10931, x10932, x10933, x10934, x10935, x10936, x10937;
  wire x10938, x10939, x10940, x10941, x10942, x10943, x10944, x10945;
  wire x10946, x10947, x10948, x10949, x10950, x10951, x10952, x10953;
  wire x10954, x10955, x10956, x10957, x10958, x10959, x10960, x10961;
  wire x10962, x10963, x10964, x10965, x10966, x10967, x10968, x10969;
  wire x10970, x10971, x10972, x10973, x10974, x10975, x10976, x10977;
  wire x10978, x10979, x10980, x10981, x10982, x10983, x10984, x10985;
  wire x10986, x10987, x10988, x10989, x10990, x10991, x10992, x10993;
  wire x10994, x10995, x10996, x10997, x10998, x10999, x11000, x11001;
  wire x11002, x11003, x11004, x11005, x11006, x11007, x11008, x11009;
  wire x11010, x11011, x11012, x11013, x11014, x11015, x11016, x11017;
  wire x11018, x11019, x11020, x11021, x11022, x11023, x11024, x11025;
  wire x11026, x11027, x11028, x11029, x11030, x11031, x11032, x11033;
  wire x11034, x11035, x11036, x11037, x11038, x11039, x11040, x11041;
  wire x11042, x11043, x11044, x11045, x11046, x11047, x11048, x11049;
  wire x11050, x11051, x11052, x11053, x11054, x11055, x11056, x11057;
  wire x11058, x11059, x11060, x11061, x11062, x11063, x11064, x11065;
  wire x11066, x11067, x11068, x11069, x11070, x11071, x11072, x11073;
  wire x11074, x11075, x11076, x11077, x11078, x11079, x11080, x11081;
  wire x11082, x11083, x11084, x11085, x11086, x11087, x11088, x11089;
  wire x11090, x11091, x11092, x11093, x11094, x11095, x11096, x11097;
  wire x11098, x11099, x11100, x11101, x11102, x11103, x11104, x11105;
  wire x11106, x11107, x11108, x11109, x11110, x11111, x11112, x11113;
  wire x11114, x11115, x11116, x11117, x11118, x11119, x11120, x11121;
  wire x11122, x11123, x11124, x11125, x11126, x11127, x11128, x11129;
  wire x11130, x11131, x11132, x11133, x11134, x11135, x11136, x11137;
  wire x11138, x11139, x11140, x11141, x11142, x11143, x11144, x11145;
  wire x11146, x11147, x11148, x11149, x11150, x11151, x11152, x11153;
  wire x11154, x11155, x11156, x11157, x11158, x11159, x11160, x11161;
  wire x11162, x11163, x11164, x11165, x11166, x11167, x11168, x11169;
  wire x11170, x11171, x11172, x11173, x11174, x11175, x11176, x11177;
  wire x11178, x11179, x11180, x11181, x11182, x11183, x11184, x11185;
  wire x11186, x11187, x11188, x11189, x11190, x11191, x11192, x11193;
  wire x11194, x11195, x11196, x11197, x11198, x11199, x11200, x11201;
  wire x11202, x11203, x11204, x11205, x11206, x11207, x11208, x11209;
  wire x11210, x11211, x11212, x11213, x11214, x11215, x11216, x11217;
  wire x11218, x11219, x11220, x11221, x11222, x11223, x11224, x11225;
  wire x11226, x11227, x11228, x11229, x11230, x11231, x11232, x11233;
  wire x11234, x11235, x11236, x11237, x11238, x11239, x11240, x11241;
  wire x11242, x11243, x11244, x11245, x11246, x11247, x11248, x11249;
  wire x11250, x11251, x11252, x11253, x11254, x11255, x11256, x11257;
  wire x11258, x11259, x11260, x11261, x11262, x11263, x11264, x11265;
  wire x11266, x11267, x11268, x11269, x11270, x11271, x11272, x11273;
  wire x11274, x11275, x11276, x11277, x11278, x11279, x11280, x11281;
  wire x11282, x11283, x11284, x11285, x11286, x11287, x11288, x11289;
  wire x11290, x11291, x11292, x11293, x11294, x11295, x11296, x11297;
  wire x11298, x11299, x11300, x11301, x11302, x11303, x11304, x11305;
  wire x11306, x11307, x11308, x11309, x11310, x11311, x11312, x11313;
  wire x11314, x11315, x11316, x11317, x11318, x11319, x11320, x11321;
  wire x11322, x11323, x11324, x11325, x11326, x11327, x11328, x11329;
  wire x11330, x11331, x11332, x11333, x11334, x11335, x11336, x11337;
  wire x11338, x11339, x11340, x11341, x11342, x11343, x11344, x11345;
  wire x11346, x11347, x11348, x11349, x11350, x11351, x11352, x11353;
  wire x11354, x11355, x11356, x11357, x11358, x11359, x11360, x11361;
  wire x11362, x11363, x11364, x11365, x11366, x11367, x11368, x11369;
  wire x11370, x11371, x11372, x11373, x11374, x11375, x11376, x11377;
  wire x11378, x11379, x11380, x11381, x11382, x11383, x11384, x11385;
  wire x11386, x11387, x11388, x11389, x11390, x11391, x11392, x11393;
  wire x11394, x11395, x11396, x11397, x11398, x11399, x11400, x11401;
  wire x11402, x11403, x11404, x11405, x11406, x11407, x11408, x11409;
  wire x11410, x11411, x11412, x11413, x11414, x11415, x11416, x11417;
  wire x11418, x11419, x11420, x11421, x11422, x11423, x11424, x11425;
  wire x11426, x11427, x11428, x11429, x11430, x11431, x11432, x11433;
  wire x11434, x11435, x11436, x11437, x11438, x11439, x11440, x11441;
  wire x11442, x11443, x11444, x11445, x11446, x11447, x11448, x11449;
  wire x11450, x11451, x11452, x11453, x11454, x11455, x11456, x11457;
  wire x11458, x11459, x11460, x11461, x11462, x11463, x11464, x11465;
  wire x11466, x11467, x11468, x11469, x11470, x11471, x11472, x11473;
  wire x11474, x11475, x11476, x11477, x11478, x11479, x11480, x11481;
  wire x11482, x11483, x11484, x11485, x11486, x11487, x11488, x11489;
  wire x11490, x11491, x11492, x11493, x11494, x11495, x11496, x11497;
  wire x11498, x11499, x11500, x11501, x11502, x11503, x11504, x11505;
  wire x11506, x11507, x11508, x11509, x11510, x11511, x11512, x11513;
  wire x11514, x11515, x11516, x11517, x11518, x11519, x11520, x11521;
  wire x11522, x11523, x11524, x11525, x11526, x11527, x11528, x11529;
  wire x11530, x11531, x11532, x11533, x11534, x11535, x11536, x11537;
  wire x11538, x11539, x11540, x11541, x11542, x11543, x11544, x11545;
  wire x11546, x11547, x11548, x11549, x11550, x11551, x11552, x11553;
  wire x11554, x11555, x11556, x11557, x11558, x11559, x11560, x11561;
  wire x11562, x11563, x11564, x11565, x11566, x11567, x11568, x11569;
  wire x11570, x11571, x11572, x11573, x11574, x11575, x11576, x11577;
  wire x11578, x11579, x11580, x11581, x11582, x11583, x11584, x11585;
  wire x11586, x11587, x11588, x11589, x11590, x11591, x11592, x11593;
  wire x11594, x11595, x11596, x11597, x11598, x11599, x11600, x11601;
  wire x11602, x11603, x11604, x11605, x11606, x11607, x11608, x11609;
  wire x11610, x11611, x11612, x11613, x11614, x11615, x11616, x11617;
  wire x11618, x11619, x11620, x11621, x11622, x11623, x11624, x11625;
  wire x11626, x11627, x11628, x11629, x11630, x11631, x11632, x11633;
  wire x11634, x11635, x11636, x11637, x11638, x11639, x11640, x11641;
  wire x11642, x11643, x11644, x11645, x11646, x11647, x11648, x11649;
  wire x11650, x11651, x11652, x11653, x11654, x11655, x11656, x11657;
  wire x11658, x11659, x11660, x11661, x11662, x11663, x11664, x11665;
  wire x11666, x11667, x11668, x11669, x11670, x11671, x11672, x11673;
  wire x11674, x11675, x11676, x11677, x11678, x11679, x11680, x11681;
  wire x11682, x11683, x11684, x11685, x11686, x11687, x11688, x11689;
  wire x11690, x11691, x11692, x11693, x11694, x11695, x11696, x11697;
  wire x11698, x11699, x11700, x11701, x11702, x11703, x11704, x11705;
  wire x11706, x11707, x11708, x11709, x11710, x11711, x11712, x11713;
  wire x11714, x11715, x11716, x11717, x11718, x11719, x11720, x11721;
  wire x11722, x11723, x11724, x11725, x11726, x11727, x11728, x11729;
  wire x11730, x11731, x11732, x11733, x11734, x11735, x11736, x11737;
  wire x11738, x11739, x11740, x11741, x11742, x11743, x11744, x11745;
  wire x11746, x11747, x11748, x11749, x11750, x11751, x11752, x11753;
  wire x11754, x11755, x11756, x11757, x11758, x11759, x11760, x11761;
  wire x11762, x11763, x11764, x11765, x11766, x11767, x11768, x11769;
  wire x11770, x11771, x11772, x11773, x11774, x11775, x11776, x11777;
  wire x11778, x11779, x11780, x11781, x11782, x11783, x11784, x11785;
  wire x11786, x11787, x11788, x11789, x11790, x11791, x11792, x11793;
  wire x11794, x11795, x11796, x11797, x11798, x11799, x11800, x11801;
  wire x11802, x11803, x11804, x11805, x11806, x11807, x11808, x11809;
  wire x11810, x11811, x11812, x11813, x11814, x11815, x11816, x11817;
  wire x11818, x11819, x11820, x11821, x11822, x11823, x11824, x11825;
  wire x11826, x11827, x11828, x11829, x11830, x11831, x11832, x11833;
  wire x11834, x11835, x11836, x11837, x11838, x11839, x11840, x11841;
  wire x11842, x11843, x11844, x11845, x11846, x11847, x11848, x11849;
  wire x11850, x11851, x11852, x11853, x11854, x11855, x11856, x11857;
  wire x11858, x11859, x11860, x11861, x11862, x11863, x11864, x11865;
  wire x11866, x11867, x11868, x11869, x11870, x11871, x11872, x11873;
  wire x11874, x11875, x11876, x11877, x11878, x11879, x11880, x11881;
  wire x11882, x11883, x11884, x11885, x11886, x11887, x11888, x11889;
  wire x11890, x11891, x11892, x11893, x11894, x11895, x11896, x11897;
  wire x11898, x11899, x11900, x11901, x11902, x11903, x11904, x11905;
  wire x11906, x11907, x11908, x11909, x11910, x11911, x11912, x11913;
  wire x11914, x11915, x11916, x11917, x11918, x11919, x11920, x11921;
  wire x11922, x11923, x11924, x11925, x11926, x11927, x11928, x11929;
  wire x11930, x11931, x11932, x11933, x11934, x11935, x11936, x11937;
  wire x11938, x11939, x11940, x11941, x11942, x11943, x11944, x11945;
  wire x11946, x11947, x11948, x11949, x11950, x11951, x11952, x11953;
  wire x11954, x11955, x11956, x11957, x11958, x11959, x11960, x11961;
  wire x11962, x11963, x11964, x11965, x11966, x11967, x11968, x11969;
  wire x11970, x11971, x11972, x11973, x11974, x11975, x11976, x11977;
  wire x11978, x11979, x11980, x11981, x11982, x11983, x11984, x11985;
  wire x11986, x11987, x11988, x11989, x11990, x11991, x11992, x11993;
  wire x11994, x11995, x11996, x11997, x11998, x11999, x12000, x12001;
  wire x12002, x12003, x12004, x12005, x12006, x12007, x12008, x12009;
  wire x12010, x12011, x12012, x12013, x12014, x12015, x12016, x12017;
  wire x12018, x12019, x12020, x12021, x12022, x12023, x12024, x12025;
  wire x12026, x12027, x12028, x12029, x12030, x12031, x12032, x12033;
  wire x12034, x12035, x12036, x12037, x12038, x12039, x12040, x12041;
  wire x12042, x12043, x12044, x12045, x12046, x12047, x12048, x12049;
  wire x12050, x12051, x12052, x12053, x12054, x12055, x12056, x12057;
  wire x12058, x12059, x12060, x12061, x12062, x12063, x12064, x12065;
  wire x12066, x12067, x12068, x12069, x12070, x12071, x12072, x12073;
  wire x12074, x12075, x12076, x12077, x12078, x12079, x12080, x12081;
  wire x12082, x12083, x12084, x12085, x12086, x12087, x12088, x12089;
  wire x12090, x12091, x12092, x12093, x12094, x12095, x12096, x12097;
  wire x12098, x12099, x12100, x12101, x12102, x12103, x12104, x12105;
  wire x12106, x12107, x12108, x12109, x12110, x12111, x12112, x12113;
  wire x12114, x12115, x12116, x12117, x12118, x12119, x12120, x12121;
  wire x12122, x12123, x12124, x12125, x12126, x12127, x12128, x12129;
  wire x12130, x12131, x12132, x12133, x12134, x12135, x12136, x12137;
  wire x12138, x12139, x12140, x12141, x12142, x12143, x12144, x12145;
  wire x12146, x12147, x12148, x12149, x12150, x12151, x12152, x12153;
  wire x12154, x12155, x12156, x12157, x12158, x12159, x12160, x12161;
  wire x12162, x12163, x12164, x12165, x12166, x12167, x12168, x12169;
  wire x12170, x12171, x12172, x12173, x12174, x12175, x12176, x12177;
  wire x12178, x12179, x12180, x12181, x12182, x12183, x12184, x12185;
  wire x12186, x12187, x12188, x12189, x12190, x12191, x12192, x12193;
  wire x12194, x12195, x12196, x12197, x12198, x12199, x12200, x12201;
  wire x12202, x12203, x12204, x12205, x12206, x12207, x12208, x12209;
  wire x12210, x12211, x12212, x12213, x12214, x12215, x12216, x12217;
  wire x12218, x12219, x12220, x12221, x12222, x12223, x12224, x12225;
  wire x12226, x12227, x12228, x12229, x12230, x12231, x12232, x12233;
  wire x12234, x12235, x12236, x12237, x12238, x12239, x12240, x12241;
  wire x12242, x12243, x12244, x12245, x12246, x12247, x12248, x12249;
  wire x12250, x12251, x12252, x12253, x12254, x12255, x12256, x12257;
  wire x12258, x12259, x12260, x12261, x12262, x12263, x12264, x12265;
  wire x12266, x12267, x12268, x12269, x12270, x12271, x12272, x12273;
  wire x12274, x12275, x12276, x12277, x12278, x12279, x12280, x12281;
  wire x12282, x12283, x12284, x12285, x12286, x12287, x12288, x12289;
  wire x12290, x12291, x12292, x12293, x12294, x12295, x12296, x12297;
  wire x12298, x12299, x12300, x12301, x12302, x12303, x12304, x12305;
  wire x12306, x12307, x12308, x12309, x12310, x12311, x12312, x12313;
  wire x12314, x12315, x12316, x12317, x12318, x12319, x12320, x12321;
  wire x12322, x12323, x12324, x12325, x12326, x12327, x12328, x12329;
  wire x12330, x12331, x12332, x12333, x12334, x12335, x12336, x12337;
  wire x12338, x12339, x12340, x12341, x12342, x12343, x12344, x12345;
  wire x12346, x12347, x12348, x12349, x12350, x12351, x12352, x12353;
  wire x12354, x12355, x12356, x12357, x12358, x12359, x12360, x12361;
  wire x12362, x12363, x12364, x12365, x12366, x12367, x12368, x12369;
  wire x12370, x12371, x12372, x12373, x12374, x12375, x12376, x12377;
  wire x12378, x12379, x12380, x12381, x12382, x12383, x12384, x12385;
  wire x12386, x12387, x12388, x12389, x12390, x12391, x12392, x12393;
  wire x12394, x12395, x12396, x12397, x12398, x12399, x12400, x12401;
  wire x12402, x12403, x12404, x12405, x12406, x12407, x12408, x12409;
  wire x12410, x12411, x12412, x12413, x12414, x12415, x12416, x12417;
  wire x12418, x12419, x12420, x12421, x12422, x12423, x12424, x12425;
  wire x12426, x12427, x12428, x12429, x12430, x12431, x12432, x12433;
  wire x12434, x12435, x12436, x12437, x12438, x12439, x12440, x12441;
  wire x12442, x12443, x12444, x12445, x12446, x12447, x12448, x12449;
  wire x12450, x12451, x12452, x12453, x12454, x12455, x12456, x12457;
  wire x12458, x12459, x12460, x12461, x12462, x12463, x12464, x12465;
  wire x12466, x12467, x12468, x12469, x12470, x12471, x12472, x12473;
  wire x12474, x12475, x12476, x12477, x12478, x12479, x12480, x12481;
  wire x12482, x12483, x12484, x12485, x12486, x12487, x12488, x12489;
  wire x12490, x12491, x12492, x12493, x12494, x12495, x12496, x12497;
  wire x12498, x12499, x12500, x12501, x12502, x12503, x12504, x12505;
  wire x12506, x12507, x12508, x12509, x12510, x12511, x12512, x12513;
  wire x12514, x12515, x12516, x12517, x12518, x12519, x12520, x12521;
  wire x12522, x12523, x12524, x12525, x12526, x12527, x12528, x12529;
  wire x12530, x12531, x12532, x12533, x12534, x12535, x12536, x12537;
  wire x12538, x12539, x12540, x12541, x12542, x12543, x12544, x12545;
  wire x12546, x12547, x12548, x12549, x12550, x12551, x12552, x12553;
  wire x12554, x12555, x12556, x12557, x12558, x12559, x12560, x12561;
  wire x12562, x12563, x12564, x12565, x12566, x12567, x12568, x12569;
  wire x12570, x12571, x12572, x12573, x12574, x12575, x12576, x12577;
  wire x12578, x12579, x12580, x12581, x12582, x12583, x12584, x12585;
  wire x12586, x12587, x12588, x12589, x12590, x12591, x12592, x12593;
  wire x12594, x12595, x12596, x12597, x12598, x12599, x12600, x12601;
  wire x12602, x12603, x12604, x12605, x12606, x12607, x12608, x12609;
  wire x12610, x12611, x12612, x12613, x12614, x12615, x12616, x12617;
  wire x12618, x12619, x12620, x12621, x12622, x12623, x12624, x12625;
  wire x12626, x12627, x12628, x12629, x12630, x12631, x12632, x12633;
  wire x12634, x12635, x12636, x12637, x12638, x12639, x12640, x12641;
  wire x12642, x12643, x12644, x12645, x12646, x12647, x12648, x12649;
  wire x12650, x12651, x12652, x12653, x12654, x12655, x12656, x12657;
  wire x12658, x12659, x12660, x12661, x12662, x12663, x12664, x12665;
  wire x12666, x12667, x12668, x12669, x12670, x12671, x12672, x12673;
  wire x12674, x12675, x12676, x12677, x12678, x12679, x12680, x12681;
  wire x12682, x12683, x12684, x12685, x12686, x12687, x12688, x12689;
  wire x12690, x12691, x12692, x12693, x12694, x12695, x12696, x12697;
  wire x12698, x12699, x12700, x12701, x12702, x12703, x12704, x12705;
  wire x12706, x12707, x12708, x12709, x12710, x12711, x12712, x12713;
  wire x12714, x12715, x12716, x12717, x12718, x12719, x12720, x12721;
  wire x12722, x12723, x12724, x12725, x12726, x12727, x12728, x12729;
  wire x12730, x12731, x12732, x12733, x12734, x12735, x12736, x12737;
  wire x12738, x12739, x12740, x12741, x12742, x12743, x12744, x12745;
  wire x12746, x12747, x12748, x12749, x12750, x12751, x12752, x12753;
  wire x12754, x12755, x12756, x12757, x12758, x12759, x12760, x12761;
  wire x12762, x12763, x12764, x12765, x12766, x12767, x12768, x12769;
  wire x12770, x12771, x12772, x12773, x12774, x12775, x12776, x12777;
  wire x12778, x12779, x12780, x12781, x12782, x12783, x12784, x12785;
  wire x12786, x12787, x12788, x12789, x12790, x12791, x12792, x12793;
  wire x12794, x12795, x12796, x12797, x12798, x12799, x12800, x12801;
  wire x12802, x12803, x12804, x12805, x12806, x12807, x12808, x12809;
  wire x12810, x12811, x12812, x12813, x12814, x12815, x12816, x12817;
  wire x12818, x12819, x12820, x12821, x12822, x12823, x12824, x12825;
  wire x12826, x12827, x12828, x12829, x12830, x12831, x12832, x12833;
  wire x12834, x12835, x12836, x12837, x12838, x12839, x12840, x12841;
  wire x12842, x12843, x12844, x12845, x12846, x12847, x12848, x12849;
  wire x12850, x12851, x12852, x12853, x12854, x12855, x12856, x12857;
  wire x12858, x12859, x12860, x12861, x12862, x12863, x12864, x12865;
  wire x12866, x12867, x12868, x12869, x12870, x12871, x12872, x12873;
  wire x12874, x12875, x12876, x12877, x12878, x12879, x12880, x12881;
  wire x12882, x12883, x12884, x12885, x12886, x12887, x12888, x12889;
  wire x12890, x12891, x12892, x12893, x12894, x12895, x12896, x12897;
  wire x12898, x12899, x12900, x12901, x12902, x12903, x12904, x12905;
  wire x12906, x12907, x12908, x12909, x12910, x12911, x12912, x12913;
  wire x12914, x12915, x12916, x12917, x12918, x12919, x12920, x12921;
  wire x12922, x12923, x12924, x12925, x12926, x12927, x12928, x12929;
  wire x12930, x12931, x12932, x12933, x12934, x12935, x12936, x12937;
  wire x12938, x12939, x12940, x12941, x12942, x12943, x12944, x12945;
  wire x12946, x12947, x12948, x12949, x12950, x12951, x12952, x12953;
  wire x12954, x12955, x12956, x12957, x12958, x12959, x12960, x12961;
  wire x12962, x12963, x12964, x12965, x12966, x12967, x12968, x12969;
  wire x12970, x12971, x12972, x12973, x12974, x12975, x12976, x12977;
  wire x12978, x12979, x12980, x12981, x12982, x12983, x12984, x12985;
  wire x12986, x12987, x12988, x12989, x12990, x12991, x12992, x12993;
  wire x12994, x12995, x12996, x12997, x12998, x12999, x13000, x13001;
  wire x13002, x13003, x13004, x13005, x13006, x13007, x13008, x13009;
  wire x13010, x13011, x13012, x13013, x13014, x13015, x13016, x13017;
  wire x13018, x13019, x13020, x13021, x13022, x13023, x13024, x13025;
  wire x13026, x13027, x13028, x13029, x13030, x13031, x13032, x13033;
  wire x13034, x13035, x13036, x13037, x13038, x13039, x13040, x13041;
  wire x13042, x13043, x13044, x13045, x13046, x13047, x13048, x13049;
  wire x13050, x13051, x13052, x13053, x13054, x13055, x13056, x13057;
  wire x13058, x13059, x13060, x13061, x13062, x13063, x13064, x13065;
  wire x13066, x13067, x13068, x13069, x13070, x13071, x13072, x13073;
  wire x13074, x13075, x13076, x13077, x13078, x13079, x13080, x13081;
  wire x13082, x13083, x13084, x13085, x13086, x13087, x13088, x13089;
  wire x13090, x13091, x13092, x13093, x13094, x13095, x13096, x13097;
  wire x13098, x13099, x13100, x13101, x13102, x13103, x13104, x13105;
  wire x13106, x13107, x13108, x13109, x13110, x13111, x13112, x13113;
  wire x13114, x13115, x13116, x13117, x13118, x13119, x13120, x13121;
  wire x13122, x13123, x13124, x13125, x13126, x13127, x13128, x13129;
  wire x13130, x13131, x13132, x13133, x13134, x13135, x13136, x13137;
  wire x13138, x13139, x13140, x13141, x13142, x13143, x13144, x13145;
  wire x13146, x13147, x13148, x13149, x13150, x13151, x13152, x13153;
  wire x13154, x13155, x13156, x13157, x13158, x13159, x13160, x13161;
  wire x13162, x13163, x13164, x13165, x13166, x13167, x13168, x13169;
  wire x13170, x13171, x13172, x13173, x13174, x13175, x13176, x13177;
  wire x13178, x13179, x13180, x13181, x13182, x13183, x13184, x13185;
  wire x13186, x13187, x13188, x13189, x13190, x13191, x13192, x13193;
  wire x13194, x13195, x13196, x13197, x13198, x13199, x13200, x13201;
  wire x13202, x13203, x13204, x13205, x13206, x13207, x13208, x13209;
  wire x13210, x13211, x13212, x13213, x13214, x13215, x13216, x13217;
  wire x13218, x13219, x13220, x13221, x13222, x13223, x13224, x13225;
  wire x13226, x13227, x13228, x13229, x13230, x13231, x13232, x13233;
  wire x13234, x13235, x13236, x13237, x13238, x13239, x13240, x13241;
  wire x13242, x13243, x13244, x13245, x13246, x13247, x13248, x13249;
  wire x13250, x13251, x13252, x13253, x13254, x13255, x13256, x13257;
  wire x13258, x13259, x13260, x13261, x13262, x13263, x13264, x13265;
  wire x13266, x13267, x13268, x13269, x13270, x13271, x13272, x13273;
  wire x13274, x13275, x13276, x13277, x13278, x13279, x13280, x13281;
  wire x13282, x13283, x13284, x13285, x13286, x13287, x13288, x13289;
  wire x13290, x13291, x13292, x13293, x13294, x13295, x13296, x13297;
  wire x13298, x13299, x13300, x13301, x13302, x13303, x13304, x13305;
  wire x13306, x13307, x13308, x13309, x13310, x13311, x13312, x13313;
  wire x13314, x13315, x13316, x13317, x13318, x13319, x13320, x13321;
  wire x13322, x13323, x13324, x13325, x13326, x13327, x13328, x13329;
  wire x13330, x13331, x13332, x13333, x13334, x13335, x13336, x13337;
  wire x13338, x13339, x13340, x13341, x13342, x13343, x13344, x13345;
  wire x13346, x13347, x13348, x13349, x13350, x13351, x13352, x13353;
  wire x13354, x13355, x13356, x13357, x13358, x13359, x13360, x13361;
  wire x13362, x13363, x13364, x13365, x13366, x13367, x13368, x13369;
  wire x13370, x13371, x13372, x13373, x13374, x13375, x13376, x13377;
  wire x13378, x13379, x13380, x13381, x13382, x13383, x13384, x13385;
  wire x13386, x13387, x13388, x13389, x13390, x13391, x13392, x13393;
  wire x13394, x13395, x13396, x13397, x13398, x13399, x13400, x13401;
  wire x13402, x13403, x13404, x13405, x13406, x13407, x13408, x13409;
  wire x13410, x13411, x13412, x13413, x13414, x13415, x13416, x13417;
  wire x13418, x13419, x13420, x13421, x13422, x13423, x13424, x13425;
  wire x13426, x13427, x13428, x13429, x13430, x13431, x13432, x13433;
  wire x13434, x13435, x13436, x13437, x13438, x13439, x13440, x13441;
  wire x13442, x13443, x13444, x13445, x13446, x13447, x13448, x13449;
  wire x13450, x13451, x13452, x13453, x13454, x13455, x13456, x13457;
  wire x13458, x13459, x13460, x13461, x13462, x13463, x13464, x13465;
  wire x13466, x13467, x13468, x13469, x13470, x13471, x13472, x13473;
  wire x13474, x13475, x13476, x13477, x13478, x13479, x13480, x13481;
  wire x13482, x13483, x13484, x13485, x13486, x13487, x13488, x13489;
  wire x13490, x13491, x13492, x13493, x13494, x13495, x13496, x13497;
  wire x13498, x13499, x13500, x13501, x13502, x13503, x13504, x13505;
  wire x13506, x13507, x13508, x13509, x13510, x13511, x13512, x13513;
  wire x13514, x13515, x13516, x13517, x13518, x13519, x13520, x13521;
  wire x13522, x13523, x13524, x13525, x13526, x13527, x13528, x13529;
  wire x13530, x13531, x13532, x13533, x13534, x13535, x13536, x13537;
  wire x13538, x13539, x13540, x13541, x13542, x13543, x13544, x13545;
  wire x13546, x13547, x13548, x13549, x13550, x13551, x13552, x13553;
  wire x13554, x13555, x13556, x13557, x13558, x13559, x13560, x13561;
  wire x13562, x13563, x13564, x13565, x13566, x13567, x13568, x13569;
  wire x13570, x13571, x13572, x13573, x13574, x13575, x13576, x13577;
  wire x13578, x13579, x13580, x13581, x13582, x13583, x13584, x13585;
  wire x13586, x13587, x13588, x13589, x13590, x13591, x13592, x13593;
  wire x13594, x13595, x13596, x13597, x13598, x13599, x13600, x13601;
  wire x13602, x13603, x13604, x13605, x13606, x13607, x13608, x13609;
  wire x13610, x13611, x13612, x13613, x13614, x13615, x13616, x13617;
  wire x13618, x13619, x13620, x13621, x13622, x13623, x13624, x13625;
  wire x13626, x13627, x13628, x13629, x13630, x13631, x13632, x13633;
  wire x13634, x13635, x13636, x13637, x13638, x13639, x13640, x13641;
  wire x13642, x13643, x13644, x13645, x13646, x13647, x13648, x13649;
  wire x13650, x13651, x13652, x13653, x13654, x13655, x13656, x13657;
  wire x13658, x13659, x13660, x13661, x13662, x13663, x13664, x13665;
  wire x13666, x13667, x13668, x13669, x13670, x13671, x13672, x13673;
  wire x13674, x13675, x13676, x13677, x13678, x13679, x13680, x13681;
  wire x13682, x13683, x13684, x13685, x13686, x13687, x13688, x13689;
  wire x13690, x13691, x13692, x13693, x13694, x13695, x13696, x13697;
  wire x13698, x13699, x13700, x13701, x13702, x13703, x13704, x13705;
  wire x13706, x13707, x13708, x13709, x13710, x13711, x13712, x13713;
  wire x13714, x13715, x13716, x13717, x13718, x13719, x13720, x13721;
  wire x13722, x13723, x13724, x13725, x13726, x13727, x13728, x13729;
  wire x13730, x13731, x13732, x13733, x13734, x13735, x13736, x13737;
  wire x13738, x13739, x13740, x13741, x13742, x13743, x13744, x13745;
  wire x13746, x13747, x13748, x13749, x13750, x13751, x13752, x13753;
  wire x13754, x13755, x13756, x13757, x13758, x13759, x13760, x13761;
  wire x13762, x13763, x13764, x13765, x13766, x13767, x13768, x13769;
  wire x13770, x13771, x13772, x13773, x13774, x13775, x13776, x13777;
  wire x13778, x13779, x13780, x13781, x13782, x13783, x13784, x13785;
  wire x13786, x13787, x13788, x13789, x13790, x13791, x13792, x13793;
  wire x13794, x13795, x13796, x13797, x13798, x13799, x13800, x13801;
  wire x13802, x13803, x13804, x13805, x13806, x13807, x13808, x13809;
  wire x13810, x13811, x13812, x13813, x13814, x13815, x13816, x13817;
  wire x13818, x13819, x13820, x13821, x13822, x13823, x13824, x13825;
  wire x13826, x13827, x13828, x13829, x13830, x13831, x13832, x13833;
  wire x13834, x13835, x13836, x13837, x13838, x13839, x13840, x13841;
  wire x13842, x13843, x13844, x13845, x13846, x13847, x13848, x13849;
  wire x13850, x13851, x13852, x13853, x13854, x13855, x13856, x13857;
  wire x13858, x13859, x13860, x13861, x13862, x13863, x13864, x13865;
  wire x13866, x13867, x13868, x13869, x13870, x13871, x13872, x13873;
  wire x13874, x13875, x13876, x13877, x13878, x13879, x13880, x13881;
  wire x13882, x13883, x13884, x13885, x13886, x13887, x13888, x13889;
  wire x13890, x13891, x13892, x13893, x13894, x13895, x13896, x13897;
  wire x13898, x13899, x13900, x13901, x13902, x13903, x13904, x13905;
  wire x13906, x13907, x13908, x13909, x13910, x13911, x13912, x13913;
  wire x13914, x13915, x13916, x13917, x13918, x13919, x13920, x13921;
  wire x13922, x13923, x13924, x13925, x13926, x13927, x13928, x13929;
  wire x13930, x13931, x13932, x13933, x13934, x13935, x13936, x13937;
  wire x13938, x13939, x13940, x13941, x13942, x13943, x13944, x13945;
  wire x13946, x13947, x13948, x13949, x13950, x13951, x13952, x13953;
  wire x13954, x13955, x13956, x13957, x13958, x13959, x13960, x13961;
  wire x13962, x13963, x13964, x13965, x13966, x13967, x13968, x13969;
  wire x13970, x13971, x13972, x13973, x13974, x13975, x13976, x13977;
  wire x13978, x13979, x13980, x13981, x13982, x13983, x13984, x13985;
  wire x13986, x13987, x13988, x13989, x13990, x13991, x13992, x13993;
  wire x13994, x13995, x13996, x13997, x13998, x13999, x14000, x14001;
  wire x14002, x14003, x14004, x14005, x14006, x14007, x14008, x14009;
  wire x14010, x14011, x14012, x14013, x14014, x14015, x14016, x14017;
  wire x14018, x14019, x14020, x14021, x14022, x14023, x14024, x14025;
  wire x14026, x14027, x14028, x14029, x14030, x14031, x14032, x14033;
  wire x14034, x14035, x14036, x14037, x14038, x14039, x14040, x14041;
  wire x14042, x14043, x14044, x14045, x14046, x14047, x14048, x14049;
  wire x14050, x14051, x14052, x14053, x14054, x14055, x14056, x14057;
  wire x14058, x14059, x14060, x14061, x14062, x14063, x14064, x14065;
  wire x14066, x14067, x14068, x14069, x14070, x14071, x14072, x14073;
  wire x14074, x14075, x14076, x14077, x14078, x14079, x14080, x14081;
  wire x14082, x14083, x14084, x14085, x14086, x14087, x14088, x14089;
  wire x14090, x14091, x14092, x14093, x14094, x14095, x14096, x14097;
  wire x14098, x14099, x14100, x14101, x14102, x14103, x14104, x14105;
  wire x14106, x14107, x14108, x14109, x14110, x14111, x14112, x14113;
  wire x14114, x14115, x14116, x14117, x14118, x14119, x14120, x14121;
  wire x14122, x14123, x14124, x14125, x14126, x14127, x14128, x14129;
  wire x14130, x14131, x14132, x14133, x14134, x14135, x14136, x14137;
  wire x14138, x14139, x14140, x14141, x14142, x14143, x14144, x14145;
  wire x14146, x14147, x14148, x14149, x14150, x14151, x14152, x14153;
  wire x14154, x14155, x14156, x14157, x14158, x14159, x14160, x14161;
  wire x14162, x14163, x14164, x14165, x14166, x14167, x14168, x14169;
  wire x14170, x14171, x14172, x14173, x14174, x14175, x14176, x14177;
  wire x14178, x14179, x14180, x14181, x14182, x14183, x14184, x14185;
  wire x14186, x14187, x14188, x14189, x14190, x14191, x14192, x14193;
  wire x14194, x14195, x14196, x14197, x14198, x14199, x14200, x14201;
  wire x14202, x14203, x14204, x14205, x14206, x14207, x14208, x14209;
  wire x14210, x14211, x14212, x14213, x14214, x14215, x14216, x14217;
  wire x14218, x14219, x14220, x14221, x14222, x14223, x14224, x14225;
  wire x14226, x14227, x14228, x14229, x14230, x14231, x14232, x14233;
  wire x14234, x14235, x14236, x14237, x14238, x14239, x14240, x14241;
  wire x14242, x14243, x14244, x14245, x14246, x14247, x14248, x14249;
  wire x14250, x14251, x14252, x14253, x14254, x14255, x14256, x14257;
  wire x14258, x14259, x14260, x14261, x14262, x14263, x14264, x14265;
  wire x14266, x14267, x14268, x14269, x14270, x14271, x14272, x14273;
  wire x14274, x14275, x14276, x14277, x14278, x14279, x14280, x14281;
  wire x14282, x14283, x14284, x14285, x14286, x14287, x14288, x14289;
  wire x14290, x14291, x14292, x14293, x14294, x14295, x14296, x14297;
  wire x14298, x14299, x14300, x14301, x14302, x14303, x14304, x14305;
  wire x14306, x14307, x14308, x14309, x14310, x14311, x14312, x14313;
  wire x14314, x14315, x14316, x14317, x14318, x14319, x14320, x14321;
  wire x14322, x14323, x14324, x14325, x14326, x14327, x14328, x14329;
  wire x14330, x14331, x14332, x14333, x14334, x14335, x14336, x14337;
  wire x14338, x14339, x14340, x14341, x14342, x14343, x14344, x14345;
  wire x14346, x14347, x14348, x14349, x14350, x14351, x14352, x14353;
  wire x14354, x14355, x14356, x14357, x14358, x14359, x14360, x14361;
  wire x14362, x14363, x14364, x14365, x14366, x14367, x14368, x14369;
  wire x14370, x14371, x14372, x14373, x14374, x14375, x14376, x14377;
  wire x14378, x14379, x14380, x14381, x14382, x14383, x14384, x14385;
  wire x14386, x14387, x14388, x14389, x14390, x14391, x14392, x14393;
  wire x14394, x14395, x14396, x14397, x14398, x14399, x14400, x14401;
  wire x14402, x14403, x14404, x14405, x14406, x14407, x14408, x14409;
  wire x14410, x14411, x14412, x14413, x14414, x14415, x14416, x14417;
  wire x14418, x14419, x14420, x14421, x14422, x14423, x14424, x14425;
  wire x14426, x14427, x14428, x14429, x14430, x14431, x14432, x14433;
  wire x14434, x14435, x14436, x14437, x14438, x14439, x14440, x14441;
  wire x14442, x14443, x14444, x14445, x14446, x14447, x14448, x14449;
  wire x14450, x14451, x14452, x14453, x14454, x14455, x14456, x14457;
  wire x14458, x14459, x14460, x14461, x14462, x14463, x14464, x14465;
  wire x14466, x14467, x14468, x14469, x14470, x14471, x14472, x14473;
  wire x14474, x14475, x14476, x14477, x14478, x14479, x14480, x14481;
  wire x14482, x14483, x14484, x14485, x14486, x14487, x14488, x14489;
  wire x14490, x14491, x14492, x14493, x14494, x14495, x14496, x14497;
  wire x14498, x14499, x14500, x14501, x14502, x14503, x14504, x14505;
  wire x14506, x14507, x14508, x14509, x14510, x14511, x14512, x14513;
  wire x14514, x14515, x14516, x14517, x14518, x14519, x14520, x14521;
  wire x14522, x14523, x14524, x14525, x14526, x14527, x14528, x14529;
  wire x14530, x14531, x14532, x14533, x14534, x14535, x14536, x14537;
  wire x14538, x14539, x14540, x14541, x14542, x14543, x14544, x14545;
  wire x14546, x14547, x14548, x14549, x14550, x14551, x14552, x14553;
  wire x14554, x14556, x14558, x14559, x14561, x14562, x14563, x14564;
  wire x14565, x14566, x14569, x14570, x14572, x14574, x14576, x14578;
  wire x14580, x14582, x14583, x14584, x14585, x14586, x14587, x14588;
  wire x14589, x14590, x14592, x14593, x14595, x14596, x14600, x14602;
  wire x14603, x14605, x14606, x14610, x14612, x14613, x14615, x14616;
  wire x14620, x14622, x14623, x14625, x14626, x14630, x14632, x14633;
  wire x14635, x14636, x14640, x14642, x14643, x14645, x14646, x14650;
  wire x14652, x14653, x14655, x14656, x14660, x14662, x14663, x14665;
  wire x14666, x14670, x14671, x14672, x14673, x14674, x14675, x14676;
  wire x14677, x14678, x14679, x14680, x14681, x14682, x14683, x14684;
  wire x14685, x14686, x14687, x14688, x14689, x14690, x14691, x14692;
  wire x14693, x14694, x14695, x14696, x14697, x14698, x14699, x14700;
  wire x14701, x14702, x14703, x14704, x14705, x14706, x14707, x14708;
  wire x14709, x14710, x14711, x14712, x14713, x14714, x14715, x14716;
  wire x14717, x14718, x14719, x14720, x14721, x14722, x14723, x14724;
  wire x14725, x14726, x14727, x14728, x14729, x14730, x14731, x14732;
  wire x14734, x14736, x14738, x14740, x14742, x14744, x14745, x14747;
  wire x14749, x14750, x14753, x14762, x14764, x14765, x14766, x14768;
  wire x14769, x14770, x14772, x14773, x14774, x14776, x14777, x14778;
  wire x14780, x14781, x14782, x14784, x14785, x14786, x14788, x14790;
  wire x14791, x14792, x14794, x14795, x14796, x14798, x14799, x14800;
  wire x14802, x14803, x14804, x14806, x14807, x14808, x14810, x14811;
  wire x14812, x14814, x14816, x14817, x14818, x14820, x14821, x14822;
  wire x14824, x14825, x14826, x14828, x14829, x14830, x14832, x14833;
  wire x14834, x14836, x14837, x14838, x14840, x14842, x14843, x14844;
  wire x14846, x14847, x14848, x14850, x14851, x14852, x14854, x14855;
  wire x14856, x14858, x14859, x14860, x14862, x14863, x14864, x14866;
  wire x14868, x14869, x14870, x14872, x14873, x14874, x14876, x14877;
  wire x14878, x14880, x14881, x14882, x14884, x14885, x14886, x14888;
  wire x14889, x14890, x14892, x14894, x14895, x14896, x14898, x14899;
  wire x14900, x14902, x14903, x14904, x14906, x14907, x14908, x14910;
  wire x14911, x14912, x14914, x14915, x14916, x14918, x14920, x14921;
  wire x14922, x14924, x14925, x14926, x14928, x14929, x14930, x14932;
  wire x14933, x14934, x14936, x14937, x14938, x14940, x14941, x14942;
  wire x14944, x14946, x14947, x14948, x14950, x14951, x14952, x14954;
  wire x14955, x14956, x14958, x14959, x14960, x14962, x14963, x14964;
  wire x14966, x14967, x14968, x14970, x14971, x14972, x14973, x14974;
  wire x14975, x14976, x14977, x14978, x14979, x14980, x14981, x14982;
  wire x14983, x14984, x14985, x14986, x14987, x14988, x14989, x14990;
  wire x14991, x14992, x14993, x14994, x14995, x14996, x14997, x14998;
  wire x14999, x15000, x15001, x15002, x15003, x15004, x15005, x15006;
  wire x15007, x15008, x15009, x15010, x15011, x15012, x15013, x15014;
  wire x15015, x15016, x15017, x15018, x15019, x15020, x15021, x15022;
  wire x15023, x15024, x15025, x15026, x15027, x15028, x15029, x15030;
  wire x15031, x15032, x15033, x15034, x15035, x15036, x15037, x15038;
  wire x15039, x15040, x15041, x15042, x15043, x15044, x15045, x15046;
  wire x15047, x15048, x15049, x15050, x15051, x15052, x15053, x15054;
  wire x15055, x15056, x15057, x15058, x15059, x15060, x15061, x15062;
  wire x15063, x15064, x15065, x15066, x15067, x15068, x15069, x15070;
  wire x15071, x15072, x15073, x15074, x15075, x15076, x15077, x15078;
  wire x15079, x15080, x15081, x15082, x15083, x15084, x15085, x15086;
  wire x15087, x15088, x15089, x15090, x15091, x15092, x15093, x15094;
  wire x15095, x15097, x15098, x15099, x15100, x15101, x15102, x15103;
  wire x15104, x15105, x15106, x15107, x15108, x15109, x15110, x15111;
  wire x15112, x15113, x15114, x15115, x15116, x15117, x15118, x15119;
  wire x15120, x15121, x15122, x15123, x15124, x15125, x15126, x15127;
  wire x15128, x15129, x15130, x15131, x15132, x15133, x15134, x15135;
  wire x15136, x15137, x15138, x15139, x15140, x15141, x15142, x15143;
  wire x15144, x15145, x15146, x15147, x15148, x15149, x15150, x15151;
  wire x15153, x15154, x15155, x15156, x15157, x15158, x15159, x15160;
  wire x15161, x15162, x15163, x15164, x15165, x15166, x15167, x15168;
  wire x15169, x15170, x15171, x15172, x15173, x15174, x15175, x15176;
  wire x15177, x15178, x15179, x15180, x15181, x15182, x15183, x15184;
  wire x15185, x15186, x15187, x15188, x15189, x15190, x15191, x15192;
  wire x15193, x15194, x15195, x15196, x15197, x15198, x15199, x15200;
  wire x15201, x15202, x15203, x15204, x15205, x15206, x15207, x15208;
  wire x15209, x15210, x15211, x15212, x15213, x15214, x15215, x15216;
  wire x15218, x15220, x15221, x15223, x15225, x15226, x15228, x15230;
  wire x15233, x15234, x15235, x15238, x15239, x15241, x15244, x15245;
  wire x15247, x15250, x15251, x15253, x15256, x15257, x15259, x15262;
  wire x15263, x15265, x15268, x15269, x15271, x15274, x15275, x15277;
  wire x15280, x15281, x15283, x15286, x15287, x15289, x15292, x15293;
  wire x15295, x15298, x15299, x15301, x15304, x15305, x15307, x15310;
  wire x15311, x15313, x15316, x15317, x15319, x15322, x15323, x15325;
  wire x15328, x15329, x15331, x15334, x15335, x15337, x15340, x15341;
  wire x15343, x15346, x15347, x15349, x15352, x15353, x15355, x15358;
  wire x15359, x15361, x15363, x15364, x15366, x15368, x15369, x15371;
  wire x15373, x15374, x15376, x15378, x15379, x15381, x15383, x15384;
  wire x15386, x15388, x15389, x15391, x15393, x15394, x15396, x15398;
  wire x15399, x15401, x15403, x15404, x15406, x15408, x15409, x15441;
  wire x15442, x15443, x15444, x15445, x15447, x15448, x15449, x15451;
  wire x15452, x15453, x15455, x15456, x15457, x15459, x15460, x15461;
  wire x15463, x15464, x15465, x15467, x15468, x15469, x15471, x15472;
  wire x15473, x15475, x15476, x15477, x15479, x15480, x15481, x15483;
  wire x15484, x15485, x15487, x15488, x15489, x15491, x15492, x15493;
  wire x15495, x15496, x15497, x15499, x15500, x15501, x15503, x15504;
  wire x15505, x15507, x15508, x15509, x15511, x15512, x15513, x15515;
  wire x15516, x15517, x15519, x15520, x15521, x15523, x15524, x15525;
  wire x15527, x15528, x15529, x15531, x15532, x15533, x15535, x15536;
  wire x15537, x15539, x15540, x15541, x15543, x15544, x15545, x15547;
  wire x15548, x15549, x15551, x15552, x15553, x15555, x15556, x15557;
  wire x15560, x15562, x15563, x15565, x15566, x15568, x15569, x15571;
  wire x15573, x15574, x15576, x15578, x15579, x15581, x15583, x15584;
  wire x15586, x15588, x15589, x15591, x15593, x15594, x15596, x15598;
  wire x15599, x15601, x15603, x15604, x15606, x15608, x15609, x15611;
  wire x15613, x15614, x15616, x15618, x15619, x15621, x15623, x15624;
  wire x15626, x15628, x15629, x15631, x15633, x15634, x15636, x15638;
  wire x15639, x15641, x15643, x15644, x15646, x15648, x15649, x15651;
  wire x15653, x15654, x15656, x15658, x15659, x15661, x15663, x15664;
  wire x15666, x15668, x15669, x15671, x15673, x15674, x15676, x15678;
  wire x15679, x15681, x15683, x15684, x15686, x15688, x15689, x15691;
  wire x15693, x15694, x15696, x15698, x15699, x15702, x15704, x15705;
  wire x15707, x15708, x15710, x15711, x15713, x15714, x15716, x15717;
  wire x15719, x15721, x15722, x15724, x15726, x15727, x15729, x15731;
  wire x15732, x15734, x15736, x15737, x15739, x15741, x15742, x15744;
  wire x15746, x15747, x15749, x15751, x15752, x15754, x15756, x15757;
  wire x15759, x15761, x15762, x15764, x15766, x15767, x15769, x15771;
  wire x15772, x15774, x15776, x15777, x15779, x15781, x15782, x15784;
  wire x15786, x15787, x15789, x15791, x15792, x15794, x15796, x15797;
  wire x15799, x15801, x15802, x15804, x15806, x15807, x15809, x15811;
  wire x15812, x15814, x15816, x15817, x15819, x15821, x15822, x15824;
  wire x15826, x15827, x15830, x15832, x15833, x15835, x15836, x15838;
  wire x15839, x15841, x15842, x15844, x15845, x15847, x15848, x15850;
  wire x15851, x15853, x15854, x15856, x15857, x15859, x15861, x15862;
  wire x15864, x15866, x15867, x15869, x15871, x15872, x15874, x15876;
  wire x15877, x15879, x15881, x15882, x15884, x15886, x15887, x15889;
  wire x15891, x15892, x15894, x15896, x15897, x15899, x15901, x15902;
  wire x15904, x15906, x15907, x15909, x15911, x15912, x15914, x15916;
  wire x15917, x15919, x15921, x15922, x15924, x15926, x15927, x15930;
  wire x15932, x15933, x15935, x15936, x15938, x15939, x15941, x15942;
  wire x15944, x15945, x15947, x15948, x15950, x15951, x15953, x15954;
  wire x15956, x15957, x15959, x15960, x15962, x15963, x15965, x15966;
  wire x15968, x15969, x15971, x15972, x15974, x15975, x15976, x15977;
  wire x15978, x15979, x15981, x15983, x15984, x15985, x15986, x15987;
  wire x15988, x15990, x15991, x15992, x15994, x15995, x15996, x15998;
  wire x15999, x16000, x16001, x16002, x16003, x16005, x16006, x16007;
  wire x16009, x16010, x16011, x16013, x16014, x16015, x16017, x16018;
  wire x16019, x16021, x16022, x16023, x16025, x16026, x16027, x16029;
  wire x16030, x16031, x16032, x16033, x16034, x16036, x16037, x16038;
  wire x16040, x16041, x16042, x16044, x16045, x16046, x16048, x16049;
  wire x16050, x16052, x16053, x16054, x16056, x16057, x16058, x16060;
  wire x16061, x16062, x16064, x16065, x16066, x16068, x16069, x16070;
  wire x16072, x16073, x16074, x16076, x16077, x16078, x16080, x16081;
  wire x16082, x16084, x16085, x16086, x16088, x16089, x16090, x16092;
  wire x16093, x16094, x16095, x16097, x16099, x16101, x16103, x16105;
  wire x16107, x16109, x16111, x16113, x16115, x16117, x16119, x16121;
  wire x16123, x16125, x16127, x16129, x16131, x16133, x16135, x16137;
  wire x16139, x16141, x16143, x16145, x16147, x16149, x16150, x16151;
  wire x16153, x16155, x16157, x16159, x16161, x16163, x16165, x16167;
  wire x16169, x16171, x16173, x16175, x16177, x16179, x16181, x16183;
  wire x16185, x16187, x16189, x16191, x16193, x16195, x16197, x16199;
  wire x16201, x16202, x16203, x16204, x16205, x16207, x16209, x16211;
  wire x16213, x16215, x16217, x16219, x16221, x16223, x16225, x16227;
  wire x16229, x16231, x16233, x16235, x16237, x16239, x16241, x16243;
  wire x16245, x16247, x16248, x16249, x16250, x16251, x16252, x16253;
  wire x16254, x16255, x16257, x16259, x16261, x16263, x16265, x16267;
  wire x16269, x16271, x16273, x16275, x16277, x16279, x16281, x16282;
  wire x16283, x16284, x16285, x16286, x16287, x16288, x16289, x16290;
  wire x16291, x16292, x16293, x16294, x16295, x16297, x16298, x16299;
  wire x16301, x16302, x16303, x16305, x16306, x16307, x16309, x16310;
  wire x16311, x16313, x16314, x16315, x16317, x16318, x16319, x16321;
  wire x16322, x16323, x16325, x16326, x16327, x16329, x16330, x16331;
  wire x16333, x16334, x16335, x16337, x16338, x16339, x16341, x16342;
  wire x16343, x16345, x16346, x16347, x16349, x16350, x16351, x16353;
  wire x16354, x16355, x16357, x16358, x16359, x16361, x16362, x16363;
  wire x16365, x16366, x16367, x16369, x16370, x16371, x16373, x16374;
  wire x16375, x16377, x16378, x16379, x16381, x16382, x16383, x16385;
  wire x16386, x16387, x16389, x16390, x16391, x16393, x16394, x16395;
  wire x16397, x16398, x16399, x16401, x16402, x16403, x16405, x16406;
  wire x16407, x16409, x16411, x16412, x16413, x16414, x16415, x16416;
  wire x16417, x16418, x16419, x16420, x16421, x16422, x16423, x16424;
  wire x16425, x16426, x16427, x16428, x16429, x16430, x16431, x16432;
  wire x16433, x16434, x16435, x16436, x16437, x16438, x16439, x16440;
  wire x16441, x16442, x16443, x16444, x16445, x16446, x16447, x16448;
  wire x16449, x16450, x16451, x16452, x16453, x16454, x16455, x16456;
  wire x16457, x16458, x16459, x16460, x16461, x16462, x16463, x16464;
  wire x16465, x16466, x16467, x16468, x16469, x16470, x16471, x16472;
  wire x16473, x16474, x16475, x16476, x16477, x16478, x16479, x16480;
  wire x16481, x16482, x16483, x16484, x16485, x16486, x16487, x16488;
  wire x16489, x16490, x16491, x16492, x16493, x16494, x16495, x16496;
  wire x16497, x16498, x16499, x16500, x16501, x16502, x16503, x16504;
  wire x16505, x16506, x16507, x16510, x16511, x16513, x16515, x16517;
  wire x16519, x16521, x16523, x16525, x16527, x16529, x16531, x16533;
  wire x16535, x16537, x16539, x16541, x16543, x16545, x16547, x16549;
  wire x16551, x16553, x16555, x16557, x16559, x16561, x16563, x16565;
  wire x16567, x16569, x16571, x16573, x16575, x16577, x16579, x16581;
  wire x16583, x16585, x16587, x16589, x16591, x16593, x16595, x16597;
  wire x16599, x16601, x16603, x16605, x16607, x16609, x16611, x16613;
  wire x16614, x16615, x16616, x16617, x16618, x16619, x16620, x16621;
  wire x16622, x16623, x16624, x16625, x16626, x16627, x16628, x16629;
  wire x16630, x16631, x16632, x16633, x16634, x16635, x16636, x16637;
  wire x16638, x16639, x16640, x16641, x16642, x16643, x16644, x16645;
  wire x16646, x16647, x16648, x16649, x16650, x16651, x16652, x16653;
  wire x16654, x16655, x16656, x16657, x16660, x16663, x16666, x16668;
  wire x16669, x16670, x16671, x16672, x16673, x16674, x16675, x16676;
  wire x16677, x16678, x16681, x16684, x16687, x16690, x16693, x16696;
  wire x16699, x16701, x16704, x16707, x16708, x16710, x16711, x16712;
  wire x16715, x16717, x16720, x16721, x16723, x16724, x16727, x16728;
  wire x16730, x16731, x16733, x16734, x16737, x16739, x16740, x16742;
  wire x16743, x16746, x16748, x16749, x16750, x16751, x16752, x16753;
  wire x16754, x16755, x16756, x16757, x16758, x16759, x16760, x16761;
  wire x16762, x16763, x16764, x16765, x16766, x16767, x16768, x16769;
  wire x16770, x16771, x16772, x16773, x16774, x16775, x16776, x16777;
  wire x16778, x16779, x16780, x16781, x16782, x16783, x16784, x16785;
  wire x16786, x16787, x16788, x16789, x16790, x16791, x16792, x16793;
  wire x16794, x16795, x16796, x16797, x16798, x16799, x16800, x16801;
  wire x16802, x16803, x16804, x16805, x16806, x16807, x16808, x16809;
  wire x16810, x16811, x16812, x16813, x16814, x16815, x16816, x16817;
  wire x16818, x16819, x16820, x16821, x16822, x16823, x16824, x16825;
  wire x16826, x16827, x16828, x16829, x16830, x16831, x16832, x16833;
  wire x16834, x16835, x16836, x16837, x16838, x16839, x16840, x16841;
  wire x16842, x16875, x16877, x16878, x16879, x16880, x16881, x16882;
  wire x16883, x16884, x16885, x16886, x16887, x16888, x16889, x16890;
  wire x16891, x16892, x16893, x16894, x16895, x16896, x16897, x16898;
  wire x16899, x16900, x16901, x16902, x16903, x16904, x16905, x16906;
  wire x16907, x16908, x16909, x16910, x16911, x16912, x16913, x16914;
  wire x16915, x16916, x16917, x16918, x16919, x16920, x16921, x16922;
  wire x16923, x16924, x16925, x16926, x16927, x16928, x16929, x16930;
  wire x16931, x16932, x16933, x16934, x16935, x16936, x16937, x16938;
  wire x16939, x16940, x16941, x16942, x16943, x16944, x16945, x16946;
  wire x16947, x16948, x16949, x16950, x16951, x16952, x16953, x16954;
  wire x16955, x16956, x16957, x16958, x16959, x16960, x16961, x16962;
  wire x16963, x16964, x16965, x16966, x16967, x16968, x16969, x16970;
  wire x16971, x16972, x16975, x16976, x16978, x16981, x16982, x16984;
  wire x16987, x16988, x16990, x16993, x16994, x16996, x16999, x17000;
  wire x17002, x17005, x17006, x17008, x17011, x17012, x17014, x17017;
  wire x17018, x17020, x17023, x17024, x17026, x17029, x17030, x17032;
  wire x17035, x17036, x17038, x17041, x17042, x17044, x17047, x17048;
  wire x17050, x17053, x17054, x17056, x17059, x17060, x17062, x17065;
  wire x17066, x17068, x17071, x17072, x17074, x17077, x17078, x17080;
  wire x17083, x17084, x17086, x17089, x17090, x17092, x17095, x17096;
  wire x17098, x17101, x17102, x17104, x17107, x17108, x17110, x17113;
  wire x17114, x17116, x17119, x17120, x17122, x17125, x17126, x17128;
  wire x17131, x17132, x17134, x17137, x17138, x17140, x17143, x17144;
  wire x17146, x17149, x17150, x17152, x17155, x17156, x17158, x17161;
  wire x17162, x17194, x17195, x17196, x17197, x17198, x17200, x17201;
  wire x17202, x17204, x17205, x17206, x17208, x17209, x17210, x17212;
  wire x17213, x17214, x17216, x17217, x17218, x17220, x17221, x17222;
  wire x17224, x17225, x17226, x17228, x17229, x17230, x17232, x17233;
  wire x17234, x17236, x17237, x17238, x17240, x17241, x17242, x17244;
  wire x17245, x17246, x17248, x17249, x17250, x17252, x17253, x17254;
  wire x17256, x17257, x17258, x17260, x17261, x17262, x17264, x17265;
  wire x17266, x17268, x17269, x17270, x17272, x17273, x17274, x17276;
  wire x17277, x17278, x17280, x17281, x17282, x17284, x17285, x17286;
  wire x17288, x17289, x17290, x17292, x17293, x17294, x17296, x17297;
  wire x17298, x17300, x17301, x17302, x17304, x17305, x17306, x17308;
  wire x17309, x17310, x17312, x17313, x17314, x17316, x17318, x17319;
  wire x17321, x17322, x17324, x17325, x17327, x17329, x17330, x17332;
  wire x17334, x17335, x17337, x17339, x17340, x17342, x17344, x17345;
  wire x17347, x17349, x17350, x17352, x17354, x17355, x17357, x17359;
  wire x17360, x17362, x17364, x17365, x17367, x17369, x17370, x17372;
  wire x17374, x17375, x17377, x17379, x17380, x17382, x17384, x17385;
  wire x17387, x17389, x17390, x17392, x17394, x17395, x17397, x17399;
  wire x17400, x17402, x17404, x17405, x17407, x17409, x17410, x17412;
  wire x17414, x17415, x17417, x17419, x17420, x17422, x17424, x17425;
  wire x17427, x17429, x17430, x17432, x17434, x17435, x17437, x17439;
  wire x17440, x17442, x17444, x17445, x17447, x17449, x17450, x17452;
  wire x17454, x17455, x17457, x17459, x17460, x17462, x17464, x17465;
  wire x17467, x17468, x17470, x17471, x17473, x17474, x17476, x17477;
  wire x17479, x17481, x17482, x17484, x17486, x17487, x17489, x17491;
  wire x17492, x17494, x17496, x17497, x17499, x17501, x17502, x17504;
  wire x17506, x17507, x17509, x17511, x17512, x17514, x17516, x17517;
  wire x17519, x17521, x17522, x17524, x17526, x17527, x17529, x17531;
  wire x17532, x17534, x17536, x17537, x17539, x17541, x17542, x17544;
  wire x17546, x17547, x17549, x17551, x17552, x17554, x17556, x17557;
  wire x17559, x17561, x17562, x17564, x17566, x17567, x17569, x17571;
  wire x17572, x17574, x17576, x17577, x17579, x17581, x17582, x17584;
  wire x17586, x17587, x17589, x17591, x17592, x17594, x17596, x17597;
  wire x17599, x17600, x17602, x17603, x17605, x17606, x17608, x17609;
  wire x17611, x17612, x17614, x17615, x17617, x17618, x17620, x17621;
  wire x17623, x17625, x17626, x17628, x17630, x17631, x17633, x17635;
  wire x17636, x17638, x17640, x17641, x17643, x17645, x17646, x17648;
  wire x17650, x17651, x17653, x17655, x17656, x17658, x17660, x17661;
  wire x17663, x17665, x17666, x17668, x17670, x17671, x17673, x17675;
  wire x17676, x17678, x17680, x17681, x17683, x17685, x17686, x17688;
  wire x17690, x17691, x17693, x17695, x17696, x17698, x17700, x17701;
  wire x17703, x17704, x17706, x17707, x17709, x17710, x17712, x17713;
  wire x17715, x17716, x17718, x17719, x17721, x17722, x17724, x17725;
  wire x17727, x17728, x17730, x17731, x17733, x17734, x17736, x17737;
  wire x17739, x17740, x17742, x17743, x17745, x17746, x17747, x17749;
  wire x17751, x17752, x17754, x17756, x17757, x17759, x17761, x17762;
  wire x17764, x17766, x17767, x17769, x17771, x17772, x17774, x17776;
  wire x17777, x17779, x17781, x17782, x17784, x17786, x17787, x17789;
  wire x17791, x17792, x17794, x17796, x17797, x17799, x17801, x17802;
  wire x17804, x17806, x17807, x17809, x17811, x17812, x17814, x17816;
  wire x17817, x17819, x17821, x17822, x17824, x17826, x17827, x17829;
  wire x17831, x17832, x17834, x17836, x17837, x17839, x17841, x17842;
  wire x17844, x17846, x17847, x17849, x17851, x17852, x17854, x17856;
  wire x17857, x17859, x17861, x17862, x17864, x17866, x17867, x17869;
  wire x17871, x17872, x17874, x17876, x17877, x17879, x17881, x17882;
  wire x17884, x17886, x17887, x17889, x17891, x17892, x17894, x17896;
  wire x17897, x17899, x17901, x17902, x17904, x17905, x17907, x17909;
  wire x17911, x17913, x17915, x17917, x17919, x17921, x17922, x17924;
  wire x17926, x17928, x17930, x17932, x17934, x17936, x17938, x17940;
  wire x17942, x17944, x17946, x17948, x17950, x17952, x17954, x17956;
  wire x17957, x17959, x17961, x17963, x17965, x17967, x17969, x17971;
  wire x17973, x17975, x17977, x17979, x17981, x17983, x17985, x17987;
  wire x17989, x17991, x17993, x17995, x17997, x17999, x18001, x18003;
  wire x18005, x18007, x18009, x18010, x18012, x18014, x18016, x18018;
  wire x18020, x18022, x18024, x18026, x18028, x18030, x18032, x18034;
  wire x18036, x18038, x18040, x18042, x18044, x18046, x18048, x18050;
  wire x18052, x18054, x18056, x18058, x18060, x18062, x18064, x18066;
  wire x18068, x18070, x18072, x18074, x18076, x18078, x18080, x18081;
  wire x18083, x18085, x18087, x18089, x18091, x18093, x18095, x18097;
  wire x18099, x18101, x18103, x18105, x18107, x18109, x18111, x18113;
  wire x18115, x18117, x18119, x18121, x18123, x18125, x18127, x18129;
  wire x18131, x18133, x18135, x18137, x18139, x18141, x18143, x18145;
  wire x18147, x18149, x18151, x18153, x18155, x18157, x18159, x18161;
  wire x18163, x18165, x18167, x18169, x18170, x18172, x18174, x18176;
  wire x18178, x18180, x18182, x18184, x18186, x18188, x18190, x18192;
  wire x18194, x18196, x18198, x18200, x18202, x18204, x18206, x18208;
  wire x18210, x18212, x18214, x18216, x18218, x18220, x18222, x18224;
  wire x18226, x18228, x18230, x18232, x18234, x18236, x18238, x18240;
  wire x18242, x18244, x18246, x18248, x18250, x18252, x18254, x18256;
  wire x18258, x18260, x18262, x18264, x18266, x18268, x18270, x18272;
  wire x18274, x18276, x18277, x18279, x18281, x18283, x18285, x18287;
  wire x18289, x18291, x18293, x18295, x18297, x18299, x18301, x18303;
  wire x18305, x18307, x18309, x18311, x18313, x18315, x18317, x18319;
  wire x18321, x18323, x18325, x18327, x18329, x18331, x18333, x18335;
  wire x18337, x18339, x18341, x18343, x18345, x18347, x18349, x18351;
  wire x18353, x18355, x18357, x18359, x18361, x18363, x18365, x18367;
  wire x18369, x18371, x18373, x18375, x18377, x18379, x18381, x18383;
  wire x18385, x18387, x18389, x18391, x18393, x18395, x18397, x18399;
  wire x18401, x18402, x18404, x18406, x18408, x18410, x18412, x18414;
  wire x18416, x18418, x18420, x18422, x18424, x18426, x18428, x18430;
  wire x18432, x18434, x18436, x18438, x18440, x18442, x18444, x18446;
  wire x18448, x18450, x18452, x18454, x18456, x18458, x18460, x18462;
  wire x18464, x18466, x18468, x18470, x18472, x18474, x18476, x18478;
  wire x18480, x18482, x18484, x18486, x18488, x18490, x18492, x18494;
  wire x18496, x18498, x18500, x18502, x18504, x18506, x18508, x18510;
  wire x18512, x18514, x18516, x18518, x18520, x18522, x18524, x18526;
  wire x18528, x18530, x18532, x18534, x18536, x18538, x18540, x18542;
  wire x18544, x18545, x18547, x18549, x18551, x18553, x18555, x18557;
  wire x18559, x18561, x18563, x18565, x18567, x18569, x18571, x18573;
  wire x18575, x18577, x18579, x18581, x18583, x18585, x18587, x18589;
  wire x18591, x18593, x18595, x18597, x18599, x18601, x18603, x18605;
  wire x18607, x18609, x18611, x18613, x18615, x18617, x18619, x18621;
  wire x18623, x18625, x18627, x18629, x18631, x18633, x18635, x18637;
  wire x18639, x18641, x18643, x18645, x18647, x18649, x18651, x18653;
  wire x18655, x18657, x18659, x18661, x18663, x18665, x18667, x18669;
  wire x18671, x18673, x18675, x18677, x18679, x18681, x18683, x18685;
  wire x18687, x18689, x18691, x18693, x18695, x18697, x18699, x18701;
  wire x18703, x18705, x18706, x18708, x18710, x18712, x18714, x18716;
  wire x18718, x18720, x18722, x18724, x18726, x18728, x18730, x18732;
  wire x18734, x18736, x18738, x18740, x18742, x18744, x18746, x18748;
  wire x18750, x18752, x18754, x18756, x18758, x18760, x18762, x18764;
  wire x18766, x18768, x18770, x18772, x18774, x18776, x18778, x18780;
  wire x18782, x18784, x18786, x18788, x18790, x18792, x18794, x18796;
  wire x18798, x18800, x18802, x18804, x18806, x18808, x18810, x18812;
  wire x18814, x18816, x18818, x18820, x18822, x18824, x18826, x18828;
  wire x18830, x18832, x18834, x18836, x18838, x18840, x18842, x18844;
  wire x18846, x18848, x18850, x18852, x18854, x18856, x18858, x18860;
  wire x18862, x18864, x18866, x18868, x18870, x18872, x18874, x18876;
  wire x18878, x18880, x18882, x18884, x18885, x18887, x18889, x18891;
  wire x18893, x18895, x18897, x18899, x18901, x18903, x18905, x18907;
  wire x18909, x18911, x18913, x18915, x18917, x18919, x18921, x18923;
  wire x18925, x18927, x18929, x18931, x18933, x18935, x18937, x18939;
  wire x18941, x18943, x18945, x18947, x18949, x18950, x18951, x18952;
  wire x18953, x18954, x18956, x18957, x18958, x18959, x18960, x18961;
  wire x18962, x18964, x18965, x18966, x18967, x18968, x18969, x18970;
  wire x18972, x18973, x18974, x18975, x18976, x18977, x18978, x18979;
  wire x18980, x18981, x18983, x18984, x18985, x18986, x18987, x18988;
  wire x18989, x18991, x18992, x18993, x18994, x18995, x18996, x18997;
  wire x18999, x19000, x19001, x19002, x19003, x19004, x19005, x19007;
  wire x19008, x19009, x19011, x19012, x19013, x19014, x19016, x19017;
  wire x19018, x19019, x19020, x19021, x19022, x19024, x19025, x19026;
  wire x19028, x19029, x19030, x19031, x19032, x19033, x19034, x19036;
  wire x19037, x19038, x19039, x19040, x19041, x19042, x19044, x19045;
  wire x19046, x19048, x19049, x19050, x19051, x19053, x19054, x19055;
  wire x19057, x19058, x19059, x19060, x19062, x19063, x19064, x19065;
  wire x19066, x19067, x19068, x19070, x19071, x19072, x19074, x19075;
  wire x19076, x19077, x19079, x19080, x19081, x19083, x19084, x19085;
  wire x19086, x19088, x19089, x19090, x19091, x19092, x19093, x19094;
  wire x19096, x19097, x19098, x19100, x19101, x19102, x19103, x19105;
  wire x19106, x19107, x19109, x19110, x19111, x19112, x19113, x19114;
  wire x19115, x19117, x19118, x19119, x19120, x19121, x19122, x19123;
  wire x19125, x19126, x19127, x19129, x19130, x19131, x19132, x19134;
  wire x19135, x19136, x19138, x19139, x19140, x19141, x19143, x19144;
  wire x19145, x19147, x19148, x19149, x19150, x19152, x19153, x19154;
  wire x19155, x19156, x19157, x19158, x19160, x19161, x19162, x19164;
  wire x19165, x19166, x19167, x19169, x19170, x19171, x19173, x19174;
  wire x19175, x19176, x19178, x19179, x19180, x19182, x19183, x19184;
  wire x19185, x19187, x19188, x19189, x19190, x19191, x19192, x19193;
  wire x19195, x19196, x19197, x19199, x19200, x19201, x19202, x19204;
  wire x19205, x19206, x19208, x19209, x19210, x19211, x19213, x19214;
  wire x19215, x19217, x19218, x19219, x19220, x19221, x19222, x19223;
  wire x19225, x19226, x19227, x19228, x19229, x19230, x19231, x19233;
  wire x19234, x19235, x19237, x19238, x19239, x19240, x19242, x19243;
  wire x19244, x19246, x19247, x19248, x19249, x19251, x19252, x19253;
  wire x19255, x19256, x19257, x19258, x19260, x19261, x19262, x19263;
  wire x19264, x19265, x19266, x19268, x19269, x19270, x19271, x19272;
  wire x19273, x19274, x19276, x19277, x19278, x19280, x19281, x19282;
  wire x19283, x19285, x19286, x19287, x19289, x19290, x19291, x19292;
  wire x19294, x19295, x19296, x19298, x19299, x19300, x19301, x19303;
  wire x19304, x19305, x19307, x19308, x19309, x19310, x19312, x19313;
  wire x19314, x19315, x19316, x19317, x19318, x19320, x19321, x19322;
  wire x19324, x19325, x19326, x19327, x19329, x19330, x19331, x19333;
  wire x19334, x19335, x19336, x19338, x19339, x19340, x19342, x19343;
  wire x19344, x19345, x19347, x19348, x19349, x19351, x19352, x19353;
  wire x19354, x19355, x19356, x19357, x19359, x19360, x19361, x19362;
  wire x19363, x19364, x19365, x19367, x19368, x19369, x19371, x19372;
  wire x19373, x19374, x19376, x19377, x19378, x19380, x19381, x19382;
  wire x19383, x19385, x19386, x19387, x19389, x19390, x19391, x19392;
  wire x19394, x19395, x19396, x19398, x19399, x19400, x19401, x19403;
  wire x19404, x19405, x19407, x19408, x19409, x19410, x19412, x19413;
  wire x19414, x19415, x19416, x19417, x19418, x19420, x19421, x19422;
  wire x19424, x19425, x19426, x19427, x19429, x19430, x19431, x19433;
  wire x19434, x19435, x19436, x19438, x19439, x19440, x19442, x19443;
  wire x19444, x19445, x19447, x19448, x19449, x19451, x19452, x19453;
  wire x19454, x19456, x19457, x19458, x19460, x19461, x19462, x19463;
  wire x19465, x19466, x19467, x19468, x19469, x19470, x19471, x19473;
  wire x19474, x19475, x19477, x19478, x19479, x19480, x19482, x19483;
  wire x19484, x19486, x19487, x19488, x19489, x19491, x19492, x19493;
  wire x19495, x19496, x19497, x19498, x19500, x19501, x19502, x19504;
  wire x19505, x19506, x19507, x19509, x19510, x19511, x19513, x19514;
  wire x19515, x19516, x19517, x19518, x19519, x19521, x19522, x19523;
  wire x19524, x19525, x19526, x19527, x19529, x19530, x19531, x19533;
  wire x19534, x19535, x19536, x19538, x19539, x19540, x19542, x19543;
  wire x19544, x19545, x19547, x19548, x19549, x19551, x19552, x19553;
  wire x19554, x19556, x19557, x19558, x19560, x19561, x19562, x19563;
  wire x19565, x19566, x19567, x19569, x19570, x19571, x19572, x19574;
  wire x19575, x19576, x19578, x19579, x19580, x19581, x19583, x19584;
  wire x19585, x19586, x19587, x19588, x19589, x19591, x19592, x19593;
  wire x19595, x19596, x19597, x19598, x19600, x19601, x19602, x19604;
  wire x19605, x19606, x19607, x19609, x19610, x19611, x19613, x19614;
  wire x19615, x19616, x19618, x19619, x19620, x19622, x19623, x19624;
  wire x19625, x19627, x19628, x19629, x19631, x19632, x19633, x19634;
  wire x19636, x19637, x19638, x19640, x19641, x19642, x19643, x19645;
  wire x19646, x19647, x19648, x19649, x19650, x19651, x19653, x19654;
  wire x19655, x19657, x19658, x19659, x19660, x19662, x19663, x19664;
  wire x19666, x19667, x19668, x19669, x19671, x19672, x19673, x19675;
  wire x19676, x19677, x19678, x19680, x19681, x19682, x19684, x19685;
  wire x19686, x19687, x19689, x19690, x19691, x19693, x19694, x19695;
  wire x19696, x19698, x19699, x19700, x19702, x19703, x19704, x19705;
  wire x19706, x19707, x19708, x19710, x19711, x19712, x19713, x19714;
  wire x19715, x19716, x19718, x19719, x19720, x19722, x19723, x19724;
  wire x19725, x19727, x19728, x19729, x19731, x19732, x19733, x19734;
  wire x19736, x19737, x19738, x19740, x19741, x19742, x19743, x19745;
  wire x19746, x19747, x19749, x19750, x19751, x19752, x19754, x19755;
  wire x19756, x19758, x19759, x19760, x19761, x19763, x19764, x19765;
  wire x19767, x19768, x19769, x19770, x19772, x19773, x19774, x19775;
  wire x19776, x19777, x19778, x19780, x19781, x19782, x19783, x19784;
  wire x19785, x19786, x19788, x19789, x19790, x19792, x19793, x19794;
  wire x19795, x19797, x19798, x19799, x19801, x19802, x19803, x19804;
  wire x19806, x19807, x19808, x19810, x19811, x19812, x19813, x19815;
  wire x19816, x19817, x19819, x19820, x19821, x19822, x19824, x19825;
  wire x19826, x19828, x19829, x19830, x19831, x19833, x19834, x19835;
  wire x19837, x19838, x19839, x19840, x19842, x19843, x19844, x19846;
  wire x19847, x19848, x19849, x19851, x19852, x19853, x19854, x19855;
  wire x19856, x19857, x19859, x19860, x19861, x19863, x19864, x19865;
  wire x19866, x19868, x19869, x19870, x19872, x19873, x19874, x19875;
  wire x19877, x19878, x19879, x19881, x19882, x19883, x19884, x19886;
  wire x19887, x19888, x19890, x19891, x19892, x19893, x19895, x19896;
  wire x19897, x19899, x19900, x19901, x19902, x19904, x19905, x19906;
  wire x19908, x19909, x19910, x19911, x19913, x19914, x19915, x19917;
  wire x19918, x19919, x19920, x19921, x19922, x19923, x19925, x19926;
  wire x19927, x19928, x19929, x19930, x19931, x19933, x19934, x19935;
  wire x19937, x19938, x19939, x19940, x19942, x19943, x19944, x19946;
  wire x19947, x19948, x19949, x19951, x19952, x19953, x19955, x19956;
  wire x19957, x19958, x19960, x19961, x19962, x19964, x19965, x19966;
  wire x19967, x19969, x19970, x19971, x19973, x19974, x19975, x19976;
  wire x19978, x19979, x19980, x19982, x19983, x19984, x19985, x19987;
  wire x19988, x19989, x19991, x19992, x19993, x19994, x19996, x19997;
  wire x19998, x20000, x20001, x20002, x20003, x20005, x20006, x20007;
  wire x20008, x20009, x20010, x20011, x20013, x20014, x20015, x20017;
  wire x20018, x20019, x20020, x20022, x20023, x20024, x20026, x20027;
  wire x20028, x20029, x20031, x20032, x20033, x20035, x20036, x20037;
  wire x20038, x20040, x20041, x20042, x20044, x20045, x20046, x20047;
  wire x20049, x20050, x20051, x20053, x20054, x20055, x20056, x20058;
  wire x20059, x20060, x20062, x20063, x20064, x20065, x20067, x20068;
  wire x20069, x20071, x20072, x20073, x20074, x20076, x20077, x20078;
  wire x20080, x20081, x20082, x20083, x20085, x20086, x20087, x20088;
  wire x20089, x20090, x20091, x20093, x20094, x20095, x20097, x20098;
  wire x20099, x20100, x20102, x20103, x20104, x20106, x20107, x20108;
  wire x20109, x20111, x20112, x20113, x20115, x20116, x20117, x20118;
  wire x20120, x20121, x20122, x20124, x20125, x20126, x20127, x20129;
  wire x20130, x20131, x20133, x20134, x20135, x20136, x20138, x20139;
  wire x20140, x20142, x20143, x20144, x20145, x20147, x20148, x20149;
  wire x20151, x20152, x20153, x20154, x20156, x20157, x20158, x20160;
  wire x20161, x20162, x20163, x20164, x20165, x20166, x20168, x20169;
  wire x20170, x20172, x20173, x20174, x20175, x20177, x20178, x20179;
  wire x20181, x20182, x20183, x20184, x20186, x20187, x20188, x20190;
  wire x20191, x20192, x20193, x20195, x20196, x20197, x20199, x20200;
  wire x20201, x20202, x20204, x20205, x20206, x20208, x20209, x20210;
  wire x20211, x20213, x20214, x20215, x20217, x20218, x20219, x20220;
  wire x20222, x20223, x20224, x20226, x20227, x20228, x20229, x20231;
  wire x20232, x20233, x20235, x20236, x20237, x20238, x20240, x20241;
  wire x20242, x20244, x20245, x20246, x20247, x20249, x20250, x20251;
  wire x20253, x20254, x20255, x20256, x20258, x20259, x20260, x20262;
  wire x20263, x20264, x20265, x20267, x20268, x20269, x20271, x20272;
  wire x20273, x20274, x20276, x20277, x20278, x20280, x20281, x20282;
  wire x20283, x20285, x20286, x20287, x20289, x20290, x20291, x20292;
  wire x20294, x20295, x20296, x20298, x20299, x20300, x20301, x20303;
  wire x20304, x20305, x20307, x20308, x20309, x20310, x20312, x20313;
  wire x20314, x20316, x20317, x20318, x20319, x20321, x20322, x20323;
  wire x20325, x20326, x20327, x20328, x20330, x20331, x20332, x20334;
  wire x20335, x20336, x20337, x20339, x20340, x20341, x20343, x20344;
  wire x20345, x20346, x20348, x20349, x20350, x20352, x20353, x20354;
  wire x20356, x20357, x20358, x20360, x20361, x20362, x20364, x20365;
  wire x20366, x20368, x20369, x20370, x20372, x20373, x20374, x20376;
  wire x20377, x20378, x20380, x20381, x20382, x20384, x20385, x20386;
  wire x20388, x20389, x20390, x20392, x20393, x20394, x20396, x20397;
  wire x20398, x20400, x20401, x20402, x20404, x20405, x20406, x20408;
  wire x20409, x20410, x20412, x20413, x20414, x20416, x20417, x20418;
  wire x20420, x20421, x20422, x20424, x20425, x20426, x20430, x20432;
  wire x20433, x20434, x20437, x20438, x20439, x20440, x20441, x20442;
  wire x20445, x20446, x20447, x20448, x20449, x20450, x20453, x20454;
  wire x20456, x20457, x20458, x20459, x20460, x20461, x20462, x20463;
  wire x20466, x20467, x20469, x20471, x20472, x20473, x20474, x20475;
  wire x20476, x20478, x20479, x20480, x20482, x20483, x20486, x20487;
  wire x20489, x20491, x20492, x20493, x20494, x20495, x20496, x20498;
  wire x20499, x20500, x20502, x20503, x20506, x20507, x20509, x20511;
  wire x20512, x20513, x20514, x20515, x20516, x20518, x20519, x20520;
  wire x20522, x20523, x20526, x20527, x20529, x20531, x20532, x20533;
  wire x20535, x20536, x20537, x20539, x20540, x20541, x20543, x20544;
  wire x20547, x20548, x20550, x20552, x20553, x20554, x20556, x20557;
  wire x20558, x20560, x20561, x20562, x20564, x20565, x20568, x20569;
  wire x20571, x20573, x20574, x20575, x20576, x20578, x20579, x20580;
  wire x20581, x20582, x20584, x20585, x20586, x20588, x20589, x20592;
  wire x20593, x20595, x20597, x20598, x20599, x20600, x20603, x20604;
  wire x20605, x20606, x20607, x20609, x20610, x20611, x20613, x20614;
  wire x20615, x20616, x20617, x20620, x20621, x20623, x20625, x20626;
  wire x20627, x20628, x20631, x20632, x20633, x20634, x20635, x20637;
  wire x20638, x20639, x20641, x20642, x20643, x20644, x20645, x20648;
  wire x20649, x20651, x20653, x20654, x20655, x20656, x20659, x20660;
  wire x20662, x20663, x20664, x20666, x20667, x20668, x20669, x20671;
  wire x20672, x20673, x20675, x20676, x20677, x20678, x20679, x20682;
  wire x20683, x20685, x20687, x20688, x20689, x20690, x20693, x20694;
  wire x20696, x20698, x20699, x20701, x20702, x20703, x20704, x20706;
  wire x20707, x20708, x20710, x20711, x20712, x20713, x20715, x20716;
  wire x20717, x20718, x20719, x20722, x20723, x20725, x20727, x20728;
  wire x20729, x20730, x20733, x20734, x20736, x20738, x20739, x20741;
  wire x20742, x20743, x20744, x20746, x20747, x20748, x20750, x20751;
  wire x20752, x20753, x20755, x20756, x20757, x20758, x20759, x20762;
  wire x20763, x20765, x20767, x20768, x20769, x20770, x20773, x20774;
  wire x20776, x20778, x20779, x20781, x20782, x20783, x20784, x20786;
  wire x20787, x20788, x20790, x20791, x20792, x20793, x20795, x20796;
  wire x20797, x20798, x20799, x20802, x20803, x20805, x20807, x20808;
  wire x20809, x20810, x20813, x20814, x20816, x20818, x20819, x20821;
  wire x20823, x20824, x20825, x20827, x20828, x20829, x20831, x20832;
  wire x20833, x20834, x20836, x20837, x20838, x20840, x20841, x20844;
  wire x20845, x20847, x20849, x20850, x20851, x20852, x20855, x20856;
  wire x20858, x20860, x20861, x20863, x20865, x20866, x20867, x20869;
  wire x20870, x20871, x20873, x20874, x20875, x20876, x20878, x20879;
  wire x20880, x20882, x20883, x20886, x20887, x20889, x20891, x20892;
  wire x20893, x20894, x20897, x20898, x20900, x20902, x20903, x20905;
  wire x20906, x20908, x20909, x20910, x20911, x20912, x20914, x20915;
  wire x20916, x20918, x20919, x20920, x20921, x20923, x20924, x20925;
  wire x20927, x20928, x20931, x20932, x20934, x20936, x20937, x20938;
  wire x20939, x20942, x20943, x20945, x20947, x20948, x20950, x20951;
  wire x20954, x20955, x20956, x20957, x20958, x20960, x20961, x20962;
  wire x20964, x20965, x20966, x20967, x20969, x20970, x20971, x20973;
  wire x20974, x20975, x20976, x20977, x20980, x20981, x20983, x20985;
  wire x20986, x20988, x20989, x20992, x20993, x20995, x20997, x20998;
  wire x21000, x21001, x21004, x21005, x21006, x21007, x21008, x21010;
  wire x21011, x21012, x21014, x21015, x21016, x21017, x21019, x21020;
  wire x21021, x21023, x21024, x21025, x21026, x21027, x21030, x21031;
  wire x21033, x21035, x21036, x21038, x21039, x21042, x21043, x21045;
  wire x21047, x21048, x21050, x21051, x21054, x21055, x21057, x21058;
  wire x21059, x21061, x21062, x21063, x21064, x21066, x21067, x21068;
  wire x21070, x21071, x21072, x21073, x21075, x21076, x21077, x21079;
  wire x21080, x21081, x21082, x21083, x21086, x21087, x21089, x21091;
  wire x21092, x21094, x21095, x21098, x21099, x21101, x21103, x21104;
  wire x21106, x21107, x21110, x21111, x21113, x21115, x21116, x21118;
  wire x21119, x21120, x21121, x21123, x21124, x21125, x21127, x21128;
  wire x21129, x21130, x21132, x21133, x21134, x21136, x21137, x21138;
  wire x21139, x21141, x21142, x21143, x21145, x21146, x21149, x21150;
  wire x21152, x21154, x21155, x21157, x21158, x21161, x21162, x21164;
  wire x21166, x21167, x21169, x21170, x21173, x21174, x21176, x21178;
  wire x21179, x21181, x21182, x21183, x21184, x21186, x21187, x21188;
  wire x21190, x21191, x21192, x21193, x21195, x21196, x21197, x21199;
  wire x21200, x21201, x21202, x21204, x21205, x21206, x21208, x21209;
  wire x21212, x21213, x21215, x21217, x21218, x21220, x21221, x21224;
  wire x21225, x21227, x21229, x21230, x21232, x21233, x21236, x21237;
  wire x21239, x21241, x21242, x21244, x21245, x21246, x21247, x21249;
  wire x21250, x21251, x21253, x21254, x21255, x21257, x21258, x21259;
  wire x21260, x21262, x21263, x21264, x21266, x21267, x21268, x21269;
  wire x21271, x21272, x21273, x21275, x21276, x21279, x21280, x21282;
  wire x21284, x21285, x21287, x21288, x21291, x21292, x21294, x21296;
  wire x21297, x21299, x21300, x21303, x21304, x21306, x21308, x21309;
  wire x21311, x21313, x21314, x21315, x21317, x21318, x21319, x21321;
  wire x21322, x21323, x21325, x21326, x21327, x21328, x21330, x21331;
  wire x21332, x21334, x21335, x21336, x21337, x21339, x21340, x21341;
  wire x21343, x21344, x21347, x21348, x21350, x21352, x21353, x21355;
  wire x21358, x21359, x21361, x21363, x21364, x21366, x21369, x21370;
  wire x21372, x21374, x21375, x21378, x21379, x21380, x21382, x21383;
  wire x21384, x21386, x21387, x21388, x21390, x21391, x21392, x21394;
  wire x21395, x21396, x21398, x21399, x21400, x21402, x21403, x21404;
  wire x21406, x21407, x21408, x21410, x21411, x21412, x21414, x21415;
  wire x21416, x21418, x21419, x21420, x21422, x21423, x21424, x21426;
  wire x21427, x21428, x21431, x21432, x21433, x21437, x21438, x21439;
  wire x21443, x21444, x21445, x21447, x21448, x21449, x21453, x21454;
  wire x21455, x21457, x21458, x21459, x21463, x21464, x21465, x21467;
  wire x21468, x21469, x21473, x21474, x21475, x21477, x21478, x21479;
  wire x21481, x21483, x21484, x21486, x21487, x21488, x21490, x21491;
  wire x21492, x21494, x21496, x21497, x21499, x21500, x21501, x21503;
  wire x21504, x21505, x21507, x21508, x21509, x21511, x21513, x21514;
  wire x21516, x21517, x21518, x21520, x21521, x21522, x21524, x21525;
  wire x21526, x21528, x21531, x21532, x21534, x21535, x21536, x21538;
  wire x21539, x21540, x21542, x21543, x21544, x21546, x21549, x21550;
  wire x21552, x21554, x21555, x21557, x21558, x21559, x21561, x21562;
  wire x21563, x21565, x21568, x21569, x21571, x21573, x21574, x21576;
  wire x21577, x21578, x21580, x21581, x21582, x21584, x21585, x21586;
  wire x21588, x21589, x21592, x21593, x21595, x21597, x21598, x21600;
  wire x21601, x21602, x21604, x21605, x21606, x21608, x21609, x21610;
  wire x21612, x21613, x21614, x21615, x21616, x21619, x21620, x21622;
  wire x21624, x21625, x21627, x21628, x21629, x21631, x21632, x21633;
  wire x21635, x21636, x21637, x21639, x21640, x21641, x21642, x21643;
  wire x21646, x21647, x21649, x21651, x21652, x21654, x21655, x21656;
  wire x21658, x21659, x21660, x21662, x21663, x21664, x21666, x21667;
  wire x21668, x21669, x21670, x21673, x21674, x21676, x21677, x21678;
  wire x21680, x21682, x21684, x21685, x21687, x21688, x21689, x21691;
  wire x21692, x21693, x21695, x21696, x21697, x21699, x21700, x21701;
  wire x21702, x21703, x21706, x21707, x21709, x21710, x21711, x21713;
  wire x21715, x21717, x21718, x21720, x21721, x21722, x21724, x21725;
  wire x21726, x21728, x21729, x21730, x21731, x21733, x21734, x21735;
  wire x21737, x21738, x21739, x21740, x21741, x21744, x21745, x21747;
  wire x21748, x21749, x21751, x21753, x21755, x21756, x21758, x21759;
  wire x21760, x21762, x21763, x21764, x21766, x21767, x21768, x21769;
  wire x21771, x21772, x21773, x21775, x21776, x21777, x21778, x21779;
  wire x21782, x21783, x21785, x21787, x21788, x21790, x21792, x21794;
  wire x21795, x21797, x21798, x21799, x21801, x21802, x21803, x21805;
  wire x21806, x21807, x21808, x21810, x21811, x21812, x21814, x21815;
  wire x21816, x21817, x21818, x21821, x21822, x21824, x21826, x21827;
  wire x21829, x21831, x21833, x21834, x21836, x21838, x21839, x21841;
  wire x21842, x21843, x21845, x21846, x21847, x21848, x21850, x21851;
  wire x21852, x21854, x21855, x21856, x21857, x21858, x21861, x21862;
  wire x21864, x21866, x21867, x21869, x21871, x21873, x21874, x21876;
  wire x21878, x21879, x21881, x21882, x21883, x21885, x21886, x21887;
  wire x21888, x21890, x21891, x21892, x21894, x21895, x21896, x21897;
  wire x21898, x21901, x21902, x21904, x21906, x21907, x21909, x21910;
  wire x21912, x21913, x21915, x21917, x21918, x21920, x21921, x21923;
  wire x21924, x21926, x21927, x21928, x21930, x21931, x21932, x21933;
  wire x21935, x21936, x21937, x21939, x21940, x21941, x21942, x21944;
  wire x21945, x21946, x21948, x21949, x21952, x21953, x21955, x21957;
  wire x21958, x21960, x21962, x21963, x21965, x21967, x21968, x21970;
  wire x21972, x21973, x21975, x21976, x21977, x21979, x21980, x21981;
  wire x21983, x21984, x21985, x21987, x21988, x21989, x21991, x21992;
  wire x21993, x21995, x21996, x21997, x21998, x21999, x22000, x22001;
  wire x22002, x22003, x22005, x22006, x22007, x22009, x22010, x22011;
  wire x22012, x22013, x22014, x22016, x22017, x22018, x22019, x22020;
  wire x22021, x22023, x22024, x22025, x22027, x22028, x22029, x22030;
  wire x22031, x22032, x22033, x22035, x22036, x22037, x22039, x22040;
  wire x22041, x22042, x22043, x22044, x22045, x22047, x22048, x22049;
  wire x22051, x22052, x22053, x22054, x22055, x22056, x22057, x22059;
  wire x22060, x22061, x22063, x22064, x22065, x22066, x22067, x22068;
  wire x22069, x22071, x22072, x22073, x22075, x22076, x22077, x22078;
  wire x22080, x22081, x22082, x22084, x22085, x22086, x22088, x22089;
  wire x22090, x22091, x22093, x22094, x22095, x22097, x22098, x22099;
  wire x22101, x22102, x22103, x22104, x22106, x22107, x22108, x22110;
  wire x22111, x22112, x22114, x22115, x22116, x22117, x22119, x22120;
  wire x22121, x22123, x22124, x22125, x22127, x22128, x22129, x22130;
  wire x22132, x22133, x22134, x22136, x22137, x22138, x22140, x22141;
  wire x22142, x22144, x22145, x22146, x22147, x22149, x22150, x22151;
  wire x22153, x22154, x22155, x22156, x22158, x22159, x22160, x22162;
  wire x22163, x22164, x22166, x22167, x22168, x22169, x22171, x22172;
  wire x22173, x22175, x22176, x22177, x22178, x22180, x22181, x22182;
  wire x22184, x22185, x22186, x22188, x22189, x22190, x22191, x22193;
  wire x22194, x22195, x22197, x22198, x22199, x22200, x22202, x22203;
  wire x22204, x22206, x22207, x22208, x22210, x22211, x22212, x22213;
  wire x22215, x22216, x22217, x22219, x22220, x22221, x22222, x22224;
  wire x22225, x22226, x22228, x22229, x22230, x22232, x22233, x22234;
  wire x22235, x22237, x22238, x22239, x22241, x22243, x22244, x22245;
  wire x22247, x22248, x22249, x22251, x22252, x22253, x22255, x22256;
  wire x22257, x22258, x22260, x22261, x22262, x22264, x22265, x22267;
  wire x22268, x22270, x22271, x22272, x22274, x22275, x22276, x22277;
  wire x22279, x22280, x22281, x22283, x22284, x22285, x22286, x22288;
  wire x22289, x22290, x22292, x22293, x22295, x22296, x22298, x22299;
  wire x22300, x22302, x22303, x22304, x22305, x22307, x22308, x22309;
  wire x22311, x22312, x22313, x22314, x22316, x22317, x22318, x22320;
  wire x22321, x22323, x22324, x22326, x22327, x22328, x22330, x22331;
  wire x22332, x22333, x22335, x22336, x22337, x22339, x22340, x22342;
  wire x22343, x22345, x22346, x22347, x22349, x22350, x22352, x22353;
  wire x22355, x22356, x22357, x22359, x22360, x22361, x22362, x22364;
  wire x22365, x22366, x22368, x22369, x22371, x22372, x22374, x22376;
  wire x22377, x22379, x22380, x22382, x22383, x22385, x22386, x22387;
  wire x22389, x22390, x22391, x22392, x22394, x22395, x22396, x22398;
  wire x22399, x22401, x22402, x22404, x22406, x22407, x22409, x22410;
  wire x22412, x22413, x22415, x22416, x22417, x22419, x22420, x22421;
  wire x22422, x22424, x22425, x22426, x22428, x22429, x22431, x22432;
  wire x22434, x22436, x22437, x22439, x22440, x22442, x22443, x22445;
  wire x22446, x22447, x22449, x22450, x22451, x22452, x22454, x22455;
  wire x22456, x22458, x22459, x22461, x22462, x22464, x22466, x22467;
  wire x22469, x22470, x22472, x22473, x22475, x22476, x22477, x22479;
  wire x22480, x22481, x22482, x22484, x22485, x22486, x22488, x22489;
  wire x22491, x22492, x22494, x22496, x22497, x22499, x22500, x22502;
  wire x22503, x22505, x22506, x22507, x22509, x22510, x22511, x22512;
  wire x22514, x22515, x22516, x22518, x22519, x22522, x22523, x22525;
  wire x22527, x22528, x22530, x22533, x22534, x22536, x22537, x22538;
  wire x22540, x22541, x22542, x22544, x22545, x22546, x22548, x22549;
  wire x22550, x22551, x22552, x22553, x22554, x22555, x22556, x22557;
  wire x22558, x22559, x22561, x22562, x22563, x22564, x22566, x22567;
  wire x22569, x22570, x22571, x22572, x22574, x22575, x22577, x22578;
  wire x22579, x22580, x22582, x22583, x22585, x22586, x22587, x22588;
  wire x22590, x22591, x22593, x22594, x22595, x22596, x22598, x22599;
  wire x22601, x22602, x22603, x22605, x22606, x22607, x22609, x22610;
  wire x22612, x22613, x22615, x22616, x22617, x22619, x22620, x22621;
  wire x22623, x22624, x22626, x22627, x22629, x22630, x22631, x22633;
  wire x22634, x22635, x22637, x22638, x22640, x22641, x22643, x22644;
  wire x22645, x22647, x22648, x22649, x22651, x22652, x22654, x22655;
  wire x22657, x22658, x22659, x22661, x22662, x22663, x22665, x22666;
  wire x22667, x22668, x22670, x22672, x22673, x22675, x22676, x22677;
  wire x22678, x22680, x22681, x22682, x22684, x22685, x22687, x22688;
  wire x22690, x22692, x22693, x22695, x22696, x22697, x22698, x22700;
  wire x22701, x22702, x22704, x22705, x22707, x22708, x22710, x22712;
  wire x22713, x22715, x22716, x22717, x22718, x22720, x22721, x22722;
  wire x22724, x22725, x22727, x22728, x22730, x22732, x22733, x22735;
  wire x22736, x22737, x22738, x22740, x22741, x22742, x22744, x22745;
  wire x22747, x22748, x22750, x22752, x22753, x22755, x22756, x22757;
  wire x22758, x22760, x22761, x22762, x22764, x22765, x22767, x22768;
  wire x22770, x22772, x22773, x22775, x22776, x22777, x22778, x22780;
  wire x22781, x22782, x22784, x22785, x22788, x22789, x22791, x22793;
  wire x22794, x22796, x22797, x22798, x22799, x22801, x22802, x22803;
  wire x22805, x22806, x22809, x22810, x22812, x22814, x22815, x22817;
  wire x22818, x22819, x22820, x22822, x22823, x22824, x22826, x22827;
  wire x22830, x22831, x22833, x22835, x22836, x22838, x22839, x22840;
  wire x22841, x22843, x22844, x22845, x22847, x22848, x22851, x22852;
  wire x22854, x22856, x22857, x22859, x22860, x22861, x22862, x22864;
  wire x22865, x22866, x22868, x22869, x22872, x22873, x22875, x22877;
  wire x22878, x22880, x22881, x22882, x22883, x22885, x22886, x22887;
  wire x22889, x22890, x22893, x22894, x22896, x22898, x22899, x22901;
  wire x22902, x22903, x22904, x22906, x22907, x22908, x22910, x22911;
  wire x22914, x22915, x22917, x22919, x22920, x22922, x22923, x22924;
  wire x22925, x22927, x22928, x22929, x22931, x22932, x22935, x22936;
  wire x22938, x22940, x22941, x22943, x22944, x22945, x22946, x22948;
  wire x22949, x22950, x22952, x22953, x22956, x22957, x22959, x22961;
  wire x22962, x22964, x22965, x22966, x22968, x22969, x22970, x22972;
  wire x22973, x22974, x22975, x22976, x22977, x22979, x22980, x22981;
  wire x22983, x22984, x22985, x22987, x22988, x22989, x22991, x22992;
  wire x22993, x22994, x22996, x22997, x22998, x23000, x23001, x23002;
  wire x23003, x23005, x23006, x23007, x23009, x23010, x23011, x23012;
  wire x23014, x23015, x23016, x23018, x23019, x23020, x23021, x23023;
  wire x23024, x23025, x23027, x23028, x23029, x23030, x23033, x23035;
  wire x23036, x23038, x23039, x23040, x23042, x23043, x23044, x23045;
  wire x23048, x23050, x23051, x23053, x23054, x23055, x23057, x23058;
  wire x23059, x23060, x23063, x23065, x23066, x23068, x23069, x23070;
  wire x23072, x23073, x23074, x23075, x23078, x23080, x23081, x23083;
  wire x23084, x23085, x23087, x23088, x23089, x23090, x23093, x23095;
  wire x23096, x23098, x23099, x23100, x23102, x23103, x23104, x23105;
  wire x23108, x23111, x23112, x23114, x23115, x23116, x23118, x23119;
  wire x23120, x23121, x23124, x23127, x23128, x23130, x23131, x23132;
  wire x23134, x23135, x23136, x23137, x23140, x23143, x23144, x23146;
  wire x23147, x23148, x23150, x23151, x23152, x23153, x23156, x23159;
  wire x23160, x23162, x23163, x23164, x23166, x23167, x23168, x23169;
  wire x23172, x23175, x23176, x23178, x23179, x23180, x23182, x23183;
  wire x23184, x23185, x23188, x23191, x23192, x23194, x23195, x23196;
  wire x23198, x23199, x23200, x23201, x23204, x23207, x23208, x23210;
  wire x23211, x23212, x23214, x23215, x23216, x23217, x23220, x23223;
  wire x23224, x23226, x23227, x23228, x23230, x23231, x23232, x23233;
  wire x23236, x23239, x23240, x23242, x23243, x23244, x23246, x23247;
  wire x23248, x23249, x23252, x23255, x23256, x23258, x23259, x23260;
  wire x23262, x23263, x23264, x23265, x23268, x23271, x23272, x23274;
  wire x23275, x23276, x23278, x23279, x23280, x23281, x23284, x23287;
  wire x23288, x23290, x23291, x23292, x23294, x23295, x23296, x23297;
  wire x23300, x23303, x23304, x23306, x23307, x23308, x23310, x23311;
  wire x23312, x23313, x23316, x23319, x23320, x23322, x23323, x23324;
  wire x23326, x23327, x23328, x23330, x23331, x23332, x23333, x23334;
  wire x23335, x23336, x23337, x23338, x23340, x23341, x23342, x23345;
  wire x23346, x23347, x23350, x23351, x23352, x23355, x23356, x23357;
  wire x23360, x23361, x23362, x23364, x23366, x23367, x23369, x23370;
  wire x23371, x23373, x23374, x23376, x23377, x23379, x23380, x23381;
  wire x23383, x23384, x23386, x23387, x23389, x23390, x23391, x23393;
  wire x23394, x23396, x23397, x23399, x23400, x23401, x23403, x23404;
  wire x23406, x23407, x23409, x23410, x23411, x23413, x23414, x23416;
  wire x23417, x23419, x23420, x23421, x23423, x23424, x23426, x23427;
  wire x23429, x23430, x23431, x23433, x23434, x23436, x23437, x23439;
  wire x23440, x23441, x23443, x23444, x23446, x23447, x23449, x23450;
  wire x23451, x23453, x23454, x23456, x23457, x23459, x23460, x23461;
  wire x23463, x23464, x23466, x23467, x23469, x23470, x23471, x23473;
  wire x23474, x23476, x23477, x23479, x23480, x23481, x23483, x23484;
  wire x23486, x23487, x23489, x23490, x23491, x23493, x23494, x23496;
  wire x23497, x23499, x23500, x23501, x23503, x23504, x23506, x23507;
  wire x23509, x23510, x23511, x23513, x23514, x23516, x23517, x23519;
  wire x23520, x23521, x23523, x23524, x23526, x23527, x23529, x23530;
  wire x23531, x23533, x23534, x23536, x23537, x23539, x23540, x23541;
  wire x23543, x23544, x23546, x23547, x23549, x23550, x23551, x23553;
  wire x23554, x23555, x23557, x23558, x23559, x23560, x23561, x23562;
  wire x23563, x23565, x23566, x23567, x23569, x23570, x23571, x23573;
  wire x23574, x23575, x23577, x23578, x23579, x23580, x23582, x23583;
  wire x23584, x23586, x23587, x23588, x23589, x23591, x23592, x23593;
  wire x23595, x23596, x23597, x23598, x23600, x23601, x23602, x23604;
  wire x23605, x23606, x23607, x23609, x23610, x23611, x23613, x23614;
  wire x23615, x23616, x23618, x23619, x23620, x23622, x23623, x23624;
  wire x23625, x23627, x23628, x23629, x23631, x23632, x23634, x23635;
  wire x23637, x23638, x23639, x23641, x23642, x23644, x23645, x23647;
  wire x23648, x23649, x23651, x23652, x23654, x23655, x23657, x23658;
  wire x23659, x23661, x23662, x23664, x23665, x23667, x23668, x23669;
  wire x23671, x23672, x23674, x23675, x23677, x23678, x23679, x23681;
  wire x23682, x23684, x23685, x23687, x23688, x23689, x23691, x23692;
  wire x23694, x23695, x23697, x23698, x23699, x23701, x23702, x23704;
  wire x23705, x23707, x23708, x23709, x23711, x23712, x23714, x23715;
  wire x23717, x23718, x23719, x23721, x23722, x23724, x23725, x23727;
  wire x23728, x23729, x23731, x23732, x23734, x23735, x23737, x23738;
  wire x23739, x23741, x23742, x23744, x23745, x23747, x23748, x23749;
  wire x23751, x23752, x23754, x23755, x23757, x23758, x23759, x23761;
  wire x23762, x23764, x23765, x23767, x23768, x23769, x23771, x23772;
  wire x23774, x23775, x23777, x23778, x23779, x23781, x23782, x23784;
  wire x23785, x23787, x23788, x23789, x23791, x23792, x23794, x23795;
  wire x23797, x23798, x23799, x23801, x23802, x23804, x23805, x23807;
  wire x23808, x23809, x23811, x23813, x23814, x23815, x23816, x23817;
  wire x23819, x23820, x23821, x23823, x23825, x23826, x23828, x23830;
  wire x23831, x23833, x23835, x23836, x23838, x23840, x23841, x23843;
  wire x23845, x23846, x23848, x23850, x23851, x23853, x23855, x23856;
  wire x23858, x23860, x23861, x23863, x23865, x23866, x23868, x23870;
  wire x23871, x23873, x23875, x23876, x23878, x23880, x23881, x23883;
  wire x23885, x23886, x23888, x23890, x23891, x23893, x23895, x23896;
  wire x23898, x23900, x23901, x23903, x23905, x23906, x23908, x23910;
  wire x23911, x23913, x23915, x23916, x23918, x23920, x23921, x23923;
  wire x23925, x23926, x23928, x23930, x23931, x23933, x23935, x23936;
  wire x23938, x23940, x23941, x23968, x23969, x23970, x23971, x23972;
  wire x23974, x23975, x23976, x23978, x23979, x23980, x23982, x23983;
  wire x23984, x23986, x23987, x23988, x23990, x23991, x23992, x23994;
  wire x23995, x23996, x23998, x23999, x24000, x24002, x24003, x24004;
  wire x24006, x24007, x24008, x24010, x24011, x24012, x24014, x24015;
  wire x24016, x24018, x24019, x24020, x24022, x24023, x24024, x24026;
  wire x24027, x24028, x24030, x24031, x24032, x24034, x24035, x24036;
  wire x24038, x24039, x24040, x24042, x24043, x24044, x24046, x24047;
  wire x24048, x24050, x24051, x24052, x24054, x24055, x24056, x24058;
  wire x24059, x24060, x24062, x24063, x24064, x24067, x24069, x24070;
  wire x24072, x24073, x24075, x24076, x24078, x24080, x24081, x24083;
  wire x24085, x24086, x24088, x24090, x24091, x24093, x24095, x24096;
  wire x24098, x24100, x24101, x24103, x24105, x24106, x24108, x24110;
  wire x24111, x24113, x24115, x24116, x24118, x24120, x24121, x24123;
  wire x24125, x24126, x24128, x24130, x24131, x24133, x24135, x24136;
  wire x24138, x24140, x24141, x24143, x24145, x24146, x24148, x24150;
  wire x24151, x24153, x24155, x24156, x24158, x24160, x24161, x24163;
  wire x24165, x24166, x24168, x24170, x24171, x24173, x24175, x24176;
  wire x24178, x24180, x24181, x24185, x24187, x24188, x24190, x24191;
  wire x24193, x24194, x24196, x24197, x24199, x24200, x24202, x24204;
  wire x24205, x24207, x24209, x24210, x24212, x24214, x24215, x24217;
  wire x24219, x24220, x24222, x24224, x24225, x24227, x24229, x24230;
  wire x24232, x24234, x24235, x24237, x24239, x24240, x24242, x24244;
  wire x24245, x24247, x24249, x24250, x24252, x24254, x24255, x24257;
  wire x24259, x24260, x24262, x24264, x24265, x24267, x24269, x24270;
  wire x24272, x24274, x24275, x24277, x24279, x24280, x24282, x24284;
  wire x24285, x24291, x24293, x24294, x24296, x24297, x24299, x24300;
  wire x24302, x24303, x24305, x24306, x24308, x24309, x24311, x24312;
  wire x24314, x24315, x24317, x24318, x24320, x24322, x24323, x24325;
  wire x24327, x24328, x24330, x24332, x24333, x24335, x24337, x24338;
  wire x24340, x24342, x24343, x24345, x24347, x24348, x24350, x24352;
  wire x24353, x24355, x24357, x24358, x24360, x24362, x24363, x24371;
  wire x24373, x24374, x24376, x24377, x24379, x24380, x24382, x24383;
  wire x24385, x24386, x24388, x24389, x24391, x24392, x24394, x24395;
  wire x24397, x24398, x24400, x24401, x24402, x24404, x24405, x24406;
  wire x24408, x24409, x24410, x24412, x24413, x24414, x24416, x24417;
  wire x24418, x24420, x24421, x24422, x24424, x24425, x24426, x24428;
  wire x24429, x24430, x24432, x24434, x24435, x24437, x24439, x24440;
  wire x24442, x24443, x24444, x24446, x24447, x24448, x24450, x24451;
  wire x24452, x24454, x24455, x24456, x24458, x24459, x24460, x24462;
  wire x24463, x24464, x24466, x24468, x24469, x24471, x24473, x24474;
  wire x24476, x24478, x24479, x24481, x24483, x24484, x24486, x24488;
  wire x24489, x24491, x24493, x24494, x24496, x24498, x24499, x24501;
  wire x24503, x24504, x24506, x24508, x24509, x24511, x24513, x24514;
  wire x24516, x24518, x24520, x24522, x24524, x24526, x24528, x24530;
  wire x24532, x24534, x24536, x24538, x24540, x24542, x24544, x24546;
  wire x24548, x24550, x24552, x24554, x24556, x24558, x24560, x24562;
  wire x24564, x24566, x24568, x24570, x24572, x24574, x24576, x24577;
  wire x24579, x24581, x24583, x24585, x24587, x24589, x24591, x24593;
  wire x24595, x24597, x24599, x24601, x24603, x24605, x24607, x24609;
  wire x24611, x24613, x24615, x24617, x24619, x24621, x24623, x24625;
  wire x24627, x24629, x24631, x24633, x24634, x24635, x24636, x24638;
  wire x24640, x24642, x24644, x24646, x24648, x24650, x24652, x24654;
  wire x24656, x24658, x24660, x24662, x24664, x24666, x24668, x24670;
  wire x24672, x24674, x24676, x24678, x24680, x24682, x24684, x24685;
  wire x24686, x24687, x24688, x24689, x24690, x24691, x24692, x24694;
  wire x24696, x24698, x24700, x24702, x24704, x24706, x24708, x24710;
  wire x24712, x24714, x24716, x24718, x24720, x24722, x24723, x24724;
  wire x24725, x24726, x24727, x24728, x24729, x24730, x24731, x24732;
  wire x24733, x24734, x24735, x24736, x24737, x24738, x24740, x24741;
  wire x24742, x24744, x24745, x24746, x24748, x24749, x24750, x24752;
  wire x24753, x24754, x24756, x24757, x24758, x24760, x24761, x24762;
  wire x24764, x24765, x24766, x24768, x24769, x24770, x24772, x24773;
  wire x24774, x24776, x24777, x24778, x24780, x24781, x24782, x24784;
  wire x24785, x24786, x24788, x24789, x24790, x24792, x24793, x24794;
  wire x24796, x24797, x24798, x24800, x24801, x24802, x24804, x24805;
  wire x24806, x24808, x24809, x24810, x24812, x24813, x24814, x24816;
  wire x24817, x24818, x24820, x24821, x24822, x24824, x24825, x24826;
  wire x24828, x24829, x24830, x24832, x24833, x24834, x24836, x24837;
  wire x24838, x24840, x24841, x24842, x24844, x24845, x24846, x24848;
  wire x24849, x24850, x24852, x24853, x24854, x24856, x24857, x24858;
  wire x24861, x24863, x24865, x24867, x24869, x24871, x24873, x24875;
  wire x24877, x24879, x24881, x24883, x24885, x24887, x24889, x24891;
  wire x24893, x24894, x24895, x24896, x24897, x24898, x24899, x24900;
  wire x24901, x24902, x24903, x24904, x24905, x24906, x24907, x24908;
  wire x24909, x24910, x24911, x24912, x24913, x24914, x24915, x24916;
  wire x24917, x24918, x24919, x24920, x24921, x24922, x24923, x24924;
  wire x24925, x24927, x24929, x24931, x24933, x24935, x24937, x24939;
  wire x24941, x24943, x24945, x24947, x24949, x24951, x24953, x24955;
  wire x24957, x24959, x24961, x24963, x24965, x24967, x24969, x24971;
  wire x24973, x24975, x24977, x24979, x24981, x24983, x24985, x24987;
  wire x24989, x24990, x24991, x24992, x24993, x24994, x24995, x24996;
  wire x24997, x24998, x24999, x25000, x25001, x25002, x25003, x25004;
  wire x25005, x25006, x25007, x25008, x25009, x25010, x25011, x25012;
  wire x25013, x25014, x25015, x25016, x25017, x25018, x25019, x25020;
  wire x25021, x25022, x25023, x25024, x25025, x25026, x25027, x25028;
  wire x25029, x25030, x25031, x25032, x25033, x25034, x25035, x25036;
  wire x25037, x25038, x25039, x25040, x25041, x25042, x25043, x25044;
  wire x25045, x25046, x25047, x25048, x25049, x25050, x25051, x25052;
  wire x25053, x25054, x25055, x25056, x25057, x25058, x25059, x25060;
  wire x25061, x25062, x25063, x25064, x25065, x25066, x25067, x25068;
  wire x25069, x25070, x25071, x25072, x25073, x25074, x25075, x25076;
  wire x25077, x25078, x25079, x25080, x25081, x25082, x25083, x25084;
  wire x25085, x25086, x25087, x25088, x25089, x25090, x25091, x25092;
  wire x25093, x25094, x25095, x25096, x25097, x25098, x25099, x25100;
  wire x25101, x25102, x25103, x25104, x25105, x25106, x25107, x25108;
  wire x25109, x25110, x25111, x25112, x25113, x25114, x25115, x25116;
  wire x25117, x25118, x25119, x25120, x25121, x25122, x25123, x25124;
  wire x25125, x25126, x25127, x25128, x25129, x25130, x25131, x25132;
  wire x25133, x25134, x25135, x25136, x25137, x25138, x25139, x25140;
  wire x25141, x25142, x25143, x25144, x25145, x25146, x25147, x25148;
  wire x25149, x25150, x25151, x25152, x25153, x25154, x25155, x25156;
  wire x25157, x25158, x25159, x25160, x25161, x25162, x25163, x25164;
  wire x25165, x25166, x25167, x25168, x25169, x25170, x25171, x25172;
  wire x25173, x25174, x25175, x25176, x25177, x25178, x25179, x25180;
  wire x25181, x25182, x25183, x25184, x25185, x25186, x25187, x25188;
  wire x25189, x25190, x25191, x25192, x25193, x25194, x25195, x25196;
  wire x25197, x25198, x25199, x25200, x25201, x25202, x25203, x25204;
  wire x25205, x25206, x25207, x25208, x25209, x25210, x25211, x25212;
  wire x25213, x25214, x25215, x25216, x25217, x25218, x25219, x25220;
  wire x25221, x25222, x25223, x25224, x25225, x25226, x25227, x25228;
  wire x25229, x25230, x25231, x25232, x25233, x25234, x25235, x25236;
  wire x25237, x25238, x25239, x25240, x25241, x25242, x25243, x25244;
  wire x25245, x25246, x25247, x25248, x25249, x25250, x25251, x25252;
  wire x25253, x25254, x25255, x25256, x25257, x25258, x25259, x25260;
  wire x25261, x25262, x25263, x25264, x25265, x25266, x25267, x25268;
  wire x25269, x25270, x25271, x25272, x25273, x25274, x25275, x25276;
  wire x25277, x25278, x25279, x25280, x25281, x25282, x25283, x25284;
  wire x25285, x25286, x25287, x25288, x25289, x25290, x25291, x25292;
  wire x25293, x25294, x25295, x25296, x25297, x25298, x25299, x25300;
  wire x25301, x25302, x25303, x25304, x25305, x25306, x25307, x25308;
  wire x25309, x25310, x25311, x25312, x25313, x25314, x25315, x25316;
  wire x25317, x25318, x25319, x25320, x25321, x25322, x25323, x25324;
  wire x25325, x25326, x25327, x25328, x25329, x25330, x25331, x25332;
  wire x25333, x25334, x25335, x25336, x25337, x25338, x25339, x25340;
  wire x25341, x25342, x25343, x25344, x25345, x25346, x25347, x25348;
  wire x25349, x25350, x25351, x25352, x25353, x25354, x25355, x25356;
  wire x25357, x25358, x25359, x25360, x25361, x25362, x25363, x25364;
  wire x25365, x25366, x25367, x25368, x25369, x25370, x25371, x25372;
  wire x25373, x25374, x25375, x25376, x25377, x25378, x25379, x25380;
  wire x25381, x25382, x25383, x25384, x25385, x25386, x25387, x25388;
  wire x25389, x25390, x25391, x25392, x25393, x25394, x25395, x25396;
  wire x25397, x25398, x25399, x25400, x25401, x25402, x25403, x25404;
  wire x25405, x25406, x25407, x25408, x25409, x25410, x25411, x25412;
  wire x25413, x25414, x25415, x25416, x25417, x25418, x25419, x25420;
  wire x25421, x25422, x25423, x25424, x25425, x25426, x25427, x25428;
  wire x25429, x25430, x25431, x25432, x25433, x25434, x25435, x25436;
  wire x25437, x25438, x25439, x25440, x25441, x25442, x25443, x25444;
  wire x25445, x25446, x25447, x25448, x25449, x25450, x25451, x25452;
  wire x25453, x25454, x25455, x25456, x25457, x25458, x25459, x25460;
  wire x25461, x25462, x25463, x25464, x25465, x25466, x25467, x25468;
  wire x25469, x25470, x25471, x25472, x25473, x25474, x25475, x25476;
  wire x25477, x25478, x25479, x25480, x25481, x25482, x25483, x25484;
  wire x25485, x25486, x25487, x25488, x25489, x25490, x25491, x25492;
  wire x25493, x25494, x25495, x25496, x25497, x25498, x25499, x25500;
  wire x25501, x25502, x25503, x25504, x25505, x25506, x25507, x25508;
  wire x25509, x25510, x25511, x25512, x25513, x25514, x25515, x25516;
  wire x25517, x25518, x25519, x25520, x25521, x25522, x25523, x25524;
  wire x25525, x25526, x25527, x25528, x25529, x25530, x25531, x25532;
  wire x25533, x25534, x25535, x25536, x25537, x25538, x25539, x25540;
  wire x25541, x25542, x25543, x25544, x25545, x25546, x25547, x25548;
  wire x25549, x25550, x25551, x25552, x25553, x25554, x25555, x25556;
  wire x25557, x25558, x25559, x25560, x25561, x25562, x25563, x25564;
  wire x25565, x25566, x25567, x25568, x25569, x25570, x25571, x25572;
  wire x25573, x25574, x25575, x25576, x25577, x25578, x25579, x25580;
  wire x25581, x25582, x25583, x25584, x25585, x25586, x25587, x25588;
  wire x25589, x25590, x25591, x25592, x25593, x25594, x25595, x25596;
  wire x25597, x25598, x25599, x25600, x25601, x25602, x25603, x25604;
  wire x25605, x25606, x25607, x25608, x25609, x25610, x25611, x25612;
  wire x25613, x25614, x25615, x25616, x25617, x25618, x25619, x25620;
  wire x25621, x25622, x25623, x25624, x25625, x25626, x25627, x25628;
  wire x25629, x25630, x25631, x25632, x25633, x25634, x25635, x25636;
  wire x25637, x25638, x25639, x25640, x25641, x25642, x25643, x25644;
  wire x25645, x25646, x25647, x25648, x25649, x25650, x25651, x25652;
  wire x25653, x25654, x25655, x25656, x25657, x25658, x25659, x25660;
  wire x25661, x25662, x25663, x25664, x25665, x25666, x25667, x25668;
  wire x25669, x25670, x25671, x25672, x25673, x25674, x25675, x25676;
  wire x25677, x25678, x25679, x25680, x25681, x25682, x25683, x25684;
  wire x25685, x25686, x25687, x25688, x25689, x25690, x25691, x25692;
  wire x25693, x25694, x25695, x25696, x25697, x25698, x25699, x25700;
  wire x25701, x25702, x25703, x25704, x25705, x25706, x25707, x25708;
  wire x25709, x25710, x25711, x25712, x25713, x25714, x25715, x25716;
  wire x25717, x25718, x25719, x25720, x25721, x25722, x25723, x25724;
  wire x25725, x25726, x25727, x25728, x25729, x25730, x25731, x25732;
  wire x25733, x25734, x25735, x25736, x25737, x25738, x25739, x25740;
  wire x25741, x25742, x25743, x25744, x25745, x25746, x25747, x25748;
  wire x25750, x25751, x25752, x25753, x25754, x25755, x25756, x25757;
  wire x25758, x25759, x25760, x25761, x25762, x25763, x25764, x25765;
  wire x25766, x25767, x25768, x25769, x25770, x25771, x25773, x25774;
  wire x25775, x25776, x25777, x25778, x25779, x25780, x25781, x25783;
  wire x25784, x25785, x25786, x25787, x25788, x25789, x25791, x25792;
  wire x25793, x25794, x25795, x25797, x25798, x25799, x25800, x25801;
  wire x25802, x25803, x25804, x25805, x25806, x25807, x25808, x25809;
  wire x25810, x25811, x25812, x25813, x25814, x25815, x25816, x25817;
  wire x25818, x25819, x25820, x25821, x25822, x25823, x25824, x25825;
  wire x25826, x25827, x25828, x25829, x25830, x25831, x25832, x25833;
  wire x25834, x25835, x25836, x25837, x25838, x25839, x25840, x25841;
  wire x25842, x25843, x25844, x25845, x25846, x25847, x25848, x25849;
  wire x25850, x25851, x25852, x25853, x25854, x25855, x25856, x25857;
  wire x25858, x25859, x25860, x25861, x25862, x25863, x25864, x25865;
  wire x25866, x25867, x25868, x25869, x25870, x25871, x25872, x25873;
  wire x25874, x25875, x25876, x25877, x25878, x25879, x25880, x25881;
  wire x25882, x25883, x25884, x25885, x25886, x25887, x25888, x25889;
  wire x25890, x25891, x25892, x25893, x25894, x25895, x25896, x25897;
  wire x25898, x25899, x25900, x25901, x25902, x25903, x25904, x25905;
  wire x25906, x25907, x25908, x25909, x25910, x25911, x25912, x25913;
  wire x25914, x25915, x25916, x25917, x25918, x25919, x25920, x25921;
  wire x25922, x25923, x25924, x25925, x25926, x25927, x25928, x25929;
  wire x25930, x25931, x25932, x25933, x25934, x25935, x25936, x25937;
  wire x25938, x25939, x25940, x25941, x25942, x25943, x25944, x25945;
  wire x25946, x25947, x25948, x25949, x25950, x25951, x25952, x25953;
  wire x25954, x25955, x25956, x25957, x25958, x25959, x25960, x25961;
  wire x25962, x25963, x25964, x25965, x25966, x25967, x25968, x25969;
  wire x25970, x25971, x25972, x25973, x25974, x25975, x25976, x25977;
  wire x25978, x25979, x25980, x25981, x25982, x25983, x25984, x25985;
  wire x25986, x25987, x25988, x25989, x25990, x25991, x25992, x25993;
  wire x25994, x25995, x25996, x25997, x25998, x25999, x26000, x26001;
  wire x26002, x26003, x26004, x26005, x26006, x26007, x26008, x26009;
  wire x26010, x26011, x26012, x26013, x26014, x26015, x26016, x26017;
  wire x26018, x26019, x26020, x26021, x26022, x26023, x26024, x26025;
  wire x26026, x26027, x26028, x26029, x26030, x26031, x26032, x26033;
  wire x26034, x26035, x26036, x26037, x26038, x26039, x26040, x26041;
  wire x26042, x26043, x26044, x26045, x26046, x26047, x26048, x26049;
  wire x26050, x26051, x26052, x26053, x26054, x26055, x26056, x26057;
  wire x26058, x26059, x26060, x26061, x26062, x26063, x26064, x26065;
  wire x26066, x26067, x26068, x26069, x26070, x26071, x26072, x26073;
  wire x26074, x26075, x26076, x26077, x26078, x26079, x26080, x26081;
  wire x26082, x26083, x26084, x26085, x26086, x26087, x26088, x26089;
  wire x26090, x26091, x26092, x26093, x26094, x26095, x26096, x26097;
  wire x26098, x26099, x26100, x26101, x26102, x26103, x26104, x26105;
  wire x26106, x26107, x26108, x26109, x26110, x26111, x26112, x26113;
  wire x26114, x26115, x26116, x26117, x26118, x26119, x26120, x26121;
  wire x26122, x26123, x26124, x26125, x26126, x26127, x26128, x26129;
  wire x26130, x26131, x26132, x26133, x26134, x26135, x26136, x26137;
  wire x26138, x26139, x26140, x26141, x26142, x26143, x26144, x26145;
  wire x26146, x26147, x26148, x26149, x26150, x26151, x26152, x26153;
  wire x26154, x26155, x26156, x26157, x26158, x26159, x26160, x26161;
  wire x26162, x26163, x26164, x26165, x26166, x26167, x26168, x26169;
  wire x26170, x26171, x26172, x26173, x26174, x26175, x26176, x26177;
  wire x26178, x26179, x26180, x26181, x26182, x26183, x26184, x26185;
  wire x26186, x26187, x26188, x26189, x26190, x26191, x26192, x26193;
  wire x26194, x26195, x26196, x26197, x26198, x26199, x26200, x26201;
  wire x26202, x26203, x26204, x26205, x26206, x26207, x26208, x26209;
  wire x26210, x26211, x26212, x26213, x26214, x26215, x26216, x26217;
  wire x26218, x26219, x26220, x26221, x26222, x26223, x26224, x26225;
  wire x26226, x26227, x26228, x26229, x26230, x26231, x26232, x26233;
  wire x26234, x26235, x26236, x26237, x26238, x26239, x26240, x26241;
  wire x26242, x26243, x26244, x26245, x26246, x26247, x26248, x26249;
  wire x26250, x26251, x26252, x26253, x26254, x26255, x26256, x26257;
  wire x26258, x26259, x26260, x26261, x26262, x26263, x26264, x26265;
  wire x26266, x26267, x26268, x26269, x26270, x26271, x26272, x26273;
  wire x26274, x26275, x26276, x26277, x26278, x26279, x26280, x26281;
  wire x26282, x26283, x26284, x26285, x26286, x26287, x26288, x26289;
  wire x26290, x26291, x26292, x26293, x26294, x26295, x26296, x26297;
  wire x26298, x26299, x26300, x26301, x26302, x26303, x26304, x26305;
  wire x26306, x26307, x26308, x26309, x26310, x26311, x26312, x26313;
  wire x26314, x26315, x26316, x26317, x26318, x26319, x26320, x26321;
  wire x26322, x26323, x26324, x26325, x26326, x26327, x26328, x26329;
  wire x26330, x26331, x26332, x26333, x26334, x26335, x26336, x26337;
  wire x26338, x26339, x26340, x26341, x26342, x26343, x26344, x26345;
  wire x26346, x26347, x26348, x26349, x26350, x26351, x26352, x26353;
  wire x26354, x26355, x26356, x26357, x26358, x26359, x26360, x26361;
  wire x26362, x26363, x26364, x26365, x26366, x26367, x26368, x26369;
  wire x26370, x26371, x26372, x26373, x26374, x26375, x26376, x26377;
  wire x26378, x26379, x26380, x26381, x26382, x26383, x26384, x26385;
  wire x26386, x26387, x26388, x26389, x26390, x26391, x26392, x26393;
  wire x26394, x26395, x26396, x26397, x26398, x26399, x26400, x26401;
  wire x26402, x26403, x26404, x26405, x26406, x26407, x26408, x26409;
  wire x26410, x26411, x26412, x26413, x26414, x26415, x26416, x26417;
  wire x26418, x26419, x26420, x26421, x26422, x26423, x26424, x26425;
  wire x26426, x26427, x26428, x26429, x26430, x26431, x26432, x26433;
  wire x26434, x26435, x26436, x26437, x26438, x26439, x26440, x26441;
  wire x26442, x26443, x26444, x26445, x26446, x26447, x26448, x26449;
  wire x26450, x26451, x26452, x26453, x26454, x26455, x26456, x26457;
  wire x26458, x26459, x26460, x26461, x26462, x26463, x26464, x26465;
  wire x26466, x26467, x26468, x26469, x26470, x26471, x26472, x26473;
  wire x26474, x26475, x26476, x26477, x26478, x26479, x26480, x26481;
  wire x26482, x26483, x26484, x26485, x26486, x26487, x26488, x26489;
  wire x26490, x26491, x26492, x26493, x26494, x26495, x26496, x26497;
  wire x26498, x26499, x26500, x26501, x26502, x26503, x26504, x26505;
  wire x26506, x26507, x26508, x26509, x26510, x26511, x26512, x26513;
  wire x26514, x26515, x26516, x26517, x26518, x26519, x26520, x26521;
  wire x26522, x26523, x26524, x26525, x26526, x26527, x26528, x26529;
  wire x26530, x26531, x26532, x26533, x26534, x26535, x26536, x26537;
  wire x26538, x26539, x26540, x26541, x26542, x26543, x26544, x26545;
  wire x26546, x26547, x26548, x26549, x26550, x26551, x26552, x26553;
  wire x26554, x26555, x26556, x26557, x26558, x26559, x26560, x26561;
  wire x26562, x26563, x26564, x26565, x26566, x26567, x26568, x26569;
  wire x26570, x26571, x26572, x26573, x26574, x26575, x26576, x26577;
  wire x26578, x26579, x26580, x26581, x26582, x26583, x26584, x26585;
  wire x26586, x26587, x26588, x26589, x26590, x26591, x26592, x26593;
  wire x26594, x26595, x26596, x26597, x26598, x26599, x26600, x26601;
  wire x26602, x26603, x26604, x26605, x26606, x26607, x26608, x26609;
  wire x26610, x26611, x26612, x26613, x26614, x26615, x26616, x26617;
  wire x26618, x26619, x26620, x26621, x26622, x26623, x26624, x26625;
  wire x26626, x26627, x26628, x26629, x26630, x26631, x26632, x26633;
  wire x26634, x26635, x26636, x26637, x26638, x26639, x26640, x26641;
  wire x26642, x26643, x26644, x26645, x26646, x26647, x26648, x26649;
  wire x26650, x26651, x26652, x26653, x26654, x26655, x26656, x26657;
  wire x26658, x26659, x26660, x26661, x26662, x26663, x26664, x26665;
  wire x26666, x26667, x26668, x26669, x26670, x26671, x26672, x26673;
  wire x26674, x26675, x26676, x26677, x26678, x26679, x26680, x26681;
  wire x26682, x26683, x26684, x26685, x26686, x26687, x26688, x26689;
  wire x26690, x26691, x26692, x26693, x26694, x26695, x26696, x26697;
  wire x26698, x26699, x26700, x26701, x26702, x26703, x26704, x26705;
  wire x26706, x26707, x26708, x26709, x26710, x26711, x26712, x26713;
  wire x26714, x26715, x26716, x26717, x26718, x26719, x26720, x26721;
  wire x26722, x26723, x26724, x26725, x26726, x26727, x26728, x26729;
  wire x26730, x26731, x26732, x26733, x26734, x26735, x26736, x26737;
  wire x26738, x26739, x26740, x26741, x26742, x26743, x26744, x26745;
  wire x26746, x26747, x26748, x26749, x26750, x26751, x26752, x26753;
  wire x26754, x26755, x26756, x26757, x26758, x26759, x26760, x26761;
  wire x26762, x26763, x26764, x26765, x26766, x26767, x26768, x26769;
  wire x26770, x26771, x26772, x26773, x26774, x26775, x26776, x26777;
  wire x26778, x26779, x26780, x26781, x26782, x26783, x26784, x26785;
  wire x26786, x26787, x26788, x26789, x26790, x26791, x26792, x26793;
  wire x26794, x26795, x26796, x26797, x26798, x26799, x26800, x26801;
  wire x26802, x26803, x26804, x26805, x26806, x26807, x26808, x26809;
  wire x26810, x26811, x26812, x26813, x26814, x26815, x26816, x26817;
  wire x26818, x26819, x26820, x26821, x26822, x26823, x26824, x26825;
  wire x26826, x26827, x26828, x26829, x26830, x26831, x26832, x26833;
  wire x26834, x26835, x26836, x26837, x26838, x26839, x26840, x26841;
  wire x26842, x26843, x26844, x26845, x26846, x26847, x26848, x26849;
  wire x26850, x26851, x26852, x26853, x26854, x26855, x26856, x26857;
  wire x26858, x26859, x26860, x26861, x26862, x26863, x26864, x26865;
  wire x26866, x26867, x26868, x26869, x26870, x26871, x26872, x26873;
  wire x26874, x26875, x26876, x26877, x26878, x26879, x26880, x26881;
  wire x26882, x26883, x26884, x26885, x26886, x26887, x26888, x26889;
  wire x26890, x26891, x26892, x26893, x26894, x26895, x26896, x26897;
  wire x26898, x26899, x26900, x26901, x26902, x26903, x26904, x26905;
  wire x26906, x26907, x26908, x26909, x26910, x26911, x26912, x26913;
  wire x26914, x26915, x26916, x26917, x26918, x26919, x26920, x26921;
  wire x26922, x26923, x26924, x26925, x26926, x26927, x26928, x26929;
  wire x26930, x26931, x26932, x26933, x26934, x26935, x26936, x26937;
  wire x26938, x26939, x26940, x26941, x26942, x26943, x26944, x26945;
  wire x26946, x26947, x26948, x26949, x26950, x26951, x26952, x26953;
  wire x26954, x26955, x26956, x26957, x26958, x26959, x26960, x26961;
  wire x26962, x26963, x26964, x26965, x26966, x26967, x26968, x26969;
  wire x26970, x26971, x26972, x26973, x26974, x26975, x26976, x26977;
  wire x26978, x26979, x26980, x26981, x26982, x26983, x26984, x26985;
  wire x26986, x26987, x26988, x26989, x26990, x26991, x26992, x26993;
  wire x26994, x26995, x26996, x26997, x26998, x26999, x27000, x27001;
  wire x27002, x27003, x27004, x27005, x27006, x27007, x27008, x27009;
  wire x27010, x27011, x27012, x27013, x27014, x27015, x27016, x27017;
  wire x27018, x27019, x27020, x27021, x27022, x27023, x27024, x27025;
  wire x27026, x27027, x27028, x27029, x27030, x27031, x27032, x27033;
  wire x27034, x27035, x27036, x27037, x27038, x27039, x27040, x27041;
  wire x27042, x27043, x27044, x27045, x27046, x27047, x27048, x27049;
  wire x27050, x27051, x27052, x27053, x27054, x27055, x27056, x27057;
  wire x27058, x27059, x27060, x27061, x27062, x27063, x27064, x27065;
  wire x27066, x27067, x27068, x27069, x27070, x27071, x27072, x27073;
  wire x27074, x27075, x27076, x27077, x27078, x27079, x27080, x27081;
  wire x27082, x27083, x27084, x27085, x27086, x27087, x27088, x27089;
  wire x27090, x27091, x27092, x27093, x27094, x27095, x27096, x27097;
  wire x27098, x27099, x27100, x27101, x27102, x27103, x27104, x27105;
  wire x27106, x27107, x27108, x27109, x27110, x27111, x27112, x27113;
  wire x27114, x27115, x27116, x27117, x27118, x27119, x27120, x27121;
  wire x27122, x27123, x27124, x27125, x27126, x27127, x27128, x27129;
  wire x27130, x27131, x27132, x27133, x27134, x27135, x27136, x27137;
  wire x27138, x27139, x27140, x27141, x27142, x27143, x27144, x27145;
  wire x27146, x27147, x27148, x27149, x27150, x27151, x27152, x27153;
  wire x27154, x27155, x27156, x27157, x27158, x27159, x27160, x27161;
  wire x27162, x27163, x27164, x27165, x27166, x27167, x27168, x27169;
  wire x27170, x27171, x27172, x27173, x27174, x27175, x27176, x27177;
  wire x27178, x27179, x27180, x27181, x27182, x27183, x27184, x27185;
  wire x27186, x27187, x27188, x27189, x27190, x27191, x27192, x27193;
  wire x27194, x27195, x27196, x27197, x27198, x27199, x27200, x27201;
  wire x27202, x27203, x27204, x27205, x27206, x27207, x27208, x27209;
  wire x27210, x27211, x27212, x27213, x27214, x27215, x27216, x27217;
  wire x27218, x27219, x27220, x27221, x27222, x27223, x27224, x27225;
  wire x27226, x27227, x27228, x27229, x27230, x27231, x27232, x27233;
  wire x27234, x27235, x27236, x27237, x27238, x27239, x27240, x27241;
  wire x27242, x27243, x27244, x27245, x27246, x27247, x27248, x27249;
  wire x27250, x27251, x27252, x27253, x27254, x27255, x27256, x27257;
  wire x27258, x27259, x27260, x27261, x27262, x27263, x27264, x27265;
  wire x27266, x27267, x27268, x27269, x27270, x27271, x27272, x27273;
  wire x27274, x27275, x27276, x27277, x27278, x27279, x27280, x27281;
  wire x27282, x27283, x27284, x27285, x27286, x27287, x27288, x27289;
  wire x27290, x27291, x27292, x27293, x27294, x27295, x27296, x27297;
  wire x27298, x27299, x27300, x27301, x27302, x27303, x27304, x27305;
  wire x27306, x27307, x27308, x27309, x27310, x27311, x27312, x27313;
  wire x27314, x27315, x27316, x27317, x27318, x27319, x27320, x27321;
  wire x27322, x27323, x27324, x27325, x27326, x27327, x27328, x27329;
  wire x27330, x27331, x27332, x27333, x27334, x27335, x27336, x27337;
  wire x27338, x27339, x27340, x27341, x27342, x27343, x27344, x27345;
  wire x27346, x27347, x27348, x27349, x27350, x27351, x27352, x27353;
  wire x27354, x27355, x27356, x27357, x27358, x27359, x27360, x27361;
  wire x27362, x27363, x27364, x27365, x27366, x27367, x27368, x27369;
  wire x27370, x27371, x27372, x27373, x27374, x27375, x27376, x27377;
  wire x27378, x27379, x27380, x27381, x27382, x27383, x27384, x27385;
  wire x27386, x27387, x27388, x27389, x27390, x27391, x27392, x27393;
  wire x27394, x27395, x27396, x27397, x27398, x27399, x27400, x27401;
  wire x27402, x27403, x27404, x27405, x27406, x27407, x27408, x27409;
  wire x27410, x27411, x27412, x27413, x27414, x27415, x27416, x27417;
  wire x27418, x27419, x27420, x27421, x27422, x27423, x27424, x27425;
  wire x27426, x27427, x27428, x27429, x27430, x27431, x27432, x27433;
  wire x27434, x27435, x27436, x27437, x27438, x27439, x27440, x27441;
  wire x27442, x27443, x27444, x27445, x27446, x27447, x27448, x27449;
  wire x27450, x27451, x27452, x27453, x27454, x27455, x27456, x27457;
  wire x27458, x27459, x27460, x27461, x27462, x27463, x27464, x27465;
  wire x27466, x27467, x27468, x27469, x27470, x27471, x27472, x27473;
  wire x27474, x27475, x27476, x27477, x27478, x27479, x27480, x27481;
  wire x27482, x27483, x27484, x27485, x27486, x27487, x27488, x27489;
  wire x27490, x27491, x27492, x27493, x27494, x27495, x27496, x27497;
  wire x27498, x27499, x27500, x27501, x27502, x27503, x27504, x27505;
  wire x27506, x27507, x27508, x27509, x27510, x27511, x27512, x27513;
  wire x27514, x27515, x27516, x27517, x27518, x27519, x27520, x27521;
  wire x27522, x27523, x27524, x27525, x27526, x27527, x27528, x27529;
  wire x27530, x27531, x27532, x27533, x27534, x27535, x27536, x27537;
  wire x27538, x27539, x27540, x27541, x27542, x27543, x27544, x27545;
  wire x27546, x27547, x27548, x27549, x27550, x27551, x27552, x27553;
  wire x27554, x27555, x27556, x27557, x27558, x27559, x27560, x27561;
  wire x27562, x27563, x27564, x27565, x27566, x27567, x27568, x27569;
  wire x27570, x27571, x27572, x27573, x27574, x27575, x27576, x27577;
  wire x27578, x27579, x27580, x27581, x27582, x27583, x27584, x27585;
  wire x27586, x27587, x27588, x27589, x27590, x27591, x27592, x27593;
  wire x27594, x27595, x27596, x27597, x27598, x27599, x27600, x27601;
  wire x27602, x27603, x27604, x27605, x27606, x27607, x27608, x27609;
  wire x27610, x27611, x27612, x27613, x27614, x27615, x27616, x27617;
  wire x27618, x27619, x27620, x27621, x27622, x27623, x27624, x27625;
  wire x27626, x27627, x27628, x27629, x27630, x27631, x27632, x27633;
  wire x27634, x27635, x27636, x27637, x27638, x27639, x27640, x27641;
  wire x27642, x27643, x27644, x27645, x27646, x27647, x27648, x27649;
  wire x27650, x27651, x27652, x27653, x27654, x27655, x27656, x27657;
  wire x27658, x27659, x27660, x27661, x27662, x27663, x27664, x27665;
  wire x27666, x27667, x27668, x27669, x27670, x27671, x27672, x27673;
  wire x27674, x27675, x27676, x27677, x27678, x27679, x27680, x27681;
  wire x27682, x27683, x27684, x27685, x27686, x27687, x27688, x27689;
  wire x27690, x27691, x27692, x27693, x27694, x27695, x27696, x27697;
  wire x27698, x27699, x27700, x27701, x27702, x27703, x27704, x27705;
  wire x27706, x27707, x27708, x27709, x27710, x27711, x27712, x27713;
  wire x27714, x27715, x27716, x27717, x27718, x27719, x27720, x27721;
  wire x27722, x27723, x27724, x27725, x27726, x27727, x27728, x27729;
  wire x27730, x27731, x27732, x27733, x27734, x27735, x27736, x27737;
  wire x27738, x27739, x27740, x27741, x27742, x27743, x27744, x27745;
  wire x27746, x27747, x27748, x27749, x27750, x27751, x27752, x27753;
  wire x27754, x27756, x27757, x27758, x27760, x27761, x27762, x27764;
  wire x27765, x27766, x27768, x27769, x27770, x27772, x27773, x27774;
  wire x27776, x27777, x27778, x27780, x27781, x27782, x27784, x27785;
  wire x27786, x27788, x27789, x27790, x27792, x27793, x27794, x27796;
  wire x27797, x27798, x27800, x27801, x27802, x27804, x27805, x27806;
  wire x27808, x27809, x27810, x27812, x27813, x27814, x27816, x27817;
  wire x27818, x27820, x27821, x27822, x27824, x27825, x27826, x27828;
  wire x27829, x27830, x27832, x27833, x27834, x27836, x27837, x27838;
  wire x27840, x27841, x27842, x27844, x27845, x27846, x27848, x27849;
  wire x27850, x27852, x27853, x27854, x27856, x27857, x27858, x27860;
  wire x27861, x27862, x27864, x27865, x27866, x27868, x27869, x27870;
  wire x27872, x27873, x27874, x27876, x27877, x27878, x27880, x27881;
  wire x27882, x27883, x27884, x27885, x27886, x27887, x27888, x27889;
  wire x27890, x27891, x27892, x27893, x27894, x27895, x27896, x27897;
  wire x27898, x27899, x27900, x27901, x27902, x27903, x27904, x27905;
  wire x27906, x27907, x27908, x27909, x27910, x27911, x27912, x27913;
  wire x27914, x27915, x27916, x27917, x27918, x27919, x27920, x27921;
  wire x27922, x27923, x27924, x27925, x27926, x27927, x27928, x27929;
  wire x27930, x27931, x27932, x27933, x27934, x27935, x27936, x27937;
  wire x27938, x27939, x27940, x27941, x27942, x27943, x27976, x27977;
  wire x27978, x27979, x27980, x27981, x27982, x27983, x27984, x27985;
  wire x27986, x27987, x27988, x27989, x27990, x27991, x27992, x27993;
  wire x27994, x27995, x27996, x27997, x27998, x27999, x28000, x28001;
  wire x28002, x28003, x28004, x28005, x28006, x28007, x28008, x28009;
  wire x28010, x28011, x28012, x28013, x28014, x28015, x28016, x28017;
  wire x28018, x28019, x28020, x28021, x28022, x28023, x28024, x28025;
  wire x28026, x28027, x28028, x28029, x28030, x28031, x28032, x28033;
  wire x28034, x28035, x28036, x28037, x28038, x28039, x28040, x28041;
  wire x28042, x28043, x28044, x28045, x28046, x28047, x28048, x28049;
  wire x28050, x28051, x28052, x28053, x28054, x28055, x28056, x28057;
  wire x28058, x28059, x28060, x28061, x28062, x28063, x28064, x28065;
  wire x28066, x28067, x28068, x28069, x28070, x28071, x28072, x28075;
  wire x28076, x28078, x28081, x28082, x28084, x28087, x28088, x28090;
  wire x28093, x28094, x28096, x28099, x28100, x28102, x28105, x28106;
  wire x28108, x28111, x28112, x28114, x28117, x28118, x28120, x28123;
  wire x28124, x28126, x28129, x28130, x28132, x28135, x28136, x28138;
  wire x28141, x28142, x28144, x28147, x28148, x28150, x28153, x28154;
  wire x28156, x28159, x28160, x28162, x28165, x28166, x28168, x28171;
  wire x28172, x28174, x28177, x28178, x28180, x28183, x28184, x28186;
  wire x28189, x28190, x28192, x28195, x28196, x28198, x28201, x28202;
  wire x28204, x28207, x28208, x28210, x28213, x28214, x28216, x28219;
  wire x28220, x28222, x28225, x28226, x28228, x28231, x28232, x28234;
  wire x28237, x28238, x28240, x28243, x28244, x28246, x28249, x28250;
  wire x28252, x28255, x28256, x28258, x28261, x28262, x28294, x28295;
  wire x28296, x28297, x28298, x28300, x28301, x28302, x28304, x28305;
  wire x28306, x28308, x28309, x28310, x28312, x28313, x28314, x28316;
  wire x28317, x28318, x28320, x28321, x28322, x28324, x28325, x28326;
  wire x28328, x28329, x28330, x28332, x28333, x28334, x28336, x28337;
  wire x28338, x28340, x28341, x28342, x28344, x28345, x28346, x28348;
  wire x28349, x28350, x28352, x28353, x28354, x28356, x28357, x28358;
  wire x28360, x28361, x28362, x28364, x28365, x28366, x28368, x28369;
  wire x28370, x28372, x28373, x28374, x28376, x28377, x28378, x28380;
  wire x28381, x28382, x28384, x28385, x28386, x28388, x28389, x28390;
  wire x28392, x28393, x28394, x28396, x28397, x28398, x28400, x28401;
  wire x28402, x28404, x28405, x28406, x28408, x28409, x28410, x28412;
  wire x28413, x28414, x28416, x28418, x28419, x28421, x28422, x28424;
  wire x28425, x28427, x28429, x28430, x28432, x28434, x28435, x28437;
  wire x28439, x28440, x28442, x28444, x28445, x28447, x28449, x28450;
  wire x28452, x28454, x28455, x28457, x28459, x28460, x28462, x28464;
  wire x28465, x28467, x28469, x28470, x28472, x28474, x28475, x28477;
  wire x28479, x28480, x28482, x28484, x28485, x28487, x28489, x28490;
  wire x28492, x28494, x28495, x28497, x28499, x28500, x28502, x28504;
  wire x28505, x28507, x28509, x28510, x28512, x28514, x28515, x28517;
  wire x28519, x28520, x28522, x28524, x28525, x28527, x28529, x28530;
  wire x28532, x28534, x28535, x28537, x28539, x28540, x28542, x28544;
  wire x28545, x28547, x28549, x28550, x28552, x28554, x28555, x28557;
  wire x28559, x28560, x28562, x28564, x28565, x28567, x28568, x28570;
  wire x28571, x28573, x28574, x28576, x28577, x28579, x28581, x28582;
  wire x28584, x28586, x28587, x28589, x28591, x28592, x28594, x28596;
  wire x28597, x28599, x28601, x28602, x28604, x28606, x28607, x28609;
  wire x28611, x28612, x28614, x28616, x28617, x28619, x28621, x28622;
  wire x28624, x28626, x28627, x28629, x28631, x28632, x28634, x28636;
  wire x28637, x28639, x28641, x28642, x28644, x28646, x28647, x28649;
  wire x28651, x28652, x28654, x28656, x28657, x28659, x28661, x28662;
  wire x28664, x28666, x28667, x28669, x28671, x28672, x28674, x28676;
  wire x28677, x28679, x28681, x28682, x28684, x28686, x28687, x28689;
  wire x28691, x28692, x28694, x28696, x28697, x28699, x28700, x28702;
  wire x28703, x28705, x28706, x28708, x28709, x28711, x28712, x28714;
  wire x28715, x28717, x28718, x28720, x28721, x28723, x28725, x28726;
  wire x28728, x28730, x28731, x28733, x28735, x28736, x28738, x28740;
  wire x28741, x28743, x28745, x28746, x28748, x28750, x28751, x28753;
  wire x28755, x28756, x28758, x28760, x28761, x28763, x28765, x28766;
  wire x28768, x28770, x28771, x28773, x28775, x28776, x28778, x28780;
  wire x28781, x28783, x28785, x28786, x28788, x28790, x28791, x28793;
  wire x28795, x28796, x28798, x28800, x28801, x28803, x28804, x28806;
  wire x28807, x28809, x28810, x28812, x28813, x28815, x28816, x28818;
  wire x28819, x28821, x28822, x28824, x28825, x28827, x28828, x28830;
  wire x28831, x28833, x28834, x28836, x28837, x28839, x28840, x28842;
  wire x28843, x28845, x28846, x28847, x28849, x28851, x28852, x28854;
  wire x28856, x28857, x28859, x28861, x28862, x28864, x28866, x28867;
  wire x28869, x28871, x28872, x28874, x28876, x28877, x28879, x28881;
  wire x28882, x28884, x28886, x28887, x28889, x28891, x28892, x28894;
  wire x28896, x28897, x28899, x28901, x28902, x28904, x28906, x28907;
  wire x28909, x28911, x28912, x28914, x28916, x28917, x28919, x28921;
  wire x28922, x28924, x28926, x28927, x28929, x28931, x28932, x28934;
  wire x28936, x28937, x28939, x28941, x28942, x28944, x28946, x28947;
  wire x28949, x28951, x28952, x28954, x28956, x28957, x28959, x28961;
  wire x28962, x28964, x28966, x28967, x28969, x28971, x28972, x28974;
  wire x28976, x28977, x28979, x28981, x28982, x28984, x28986, x28987;
  wire x28989, x28991, x28992, x28994, x28996, x28997, x28999, x29001;
  wire x29002, x29004, x29005, x29007, x29009, x29011, x29013, x29015;
  wire x29017, x29019, x29021, x29022, x29024, x29026, x29028, x29030;
  wire x29032, x29034, x29036, x29038, x29040, x29042, x29044, x29046;
  wire x29048, x29050, x29052, x29054, x29056, x29057, x29059, x29061;
  wire x29063, x29065, x29067, x29069, x29071, x29073, x29075, x29077;
  wire x29079, x29081, x29083, x29085, x29087, x29089, x29091, x29093;
  wire x29095, x29097, x29099, x29101, x29103, x29105, x29107, x29109;
  wire x29110, x29112, x29114, x29116, x29118, x29120, x29122, x29124;
  wire x29126, x29128, x29130, x29132, x29134, x29136, x29138, x29140;
  wire x29142, x29144, x29146, x29148, x29150, x29152, x29154, x29156;
  wire x29158, x29160, x29162, x29164, x29166, x29168, x29170, x29172;
  wire x29174, x29176, x29178, x29180, x29181, x29183, x29185, x29187;
  wire x29189, x29191, x29193, x29195, x29197, x29199, x29201, x29203;
  wire x29205, x29207, x29209, x29211, x29213, x29215, x29217, x29219;
  wire x29221, x29223, x29225, x29227, x29229, x29231, x29233, x29235;
  wire x29237, x29239, x29241, x29243, x29245, x29247, x29249, x29251;
  wire x29253, x29255, x29257, x29259, x29261, x29263, x29265, x29267;
  wire x29269, x29270, x29272, x29274, x29276, x29278, x29280, x29282;
  wire x29284, x29286, x29288, x29290, x29292, x29294, x29296, x29298;
  wire x29300, x29302, x29304, x29306, x29308, x29310, x29312, x29314;
  wire x29316, x29318, x29320, x29322, x29324, x29326, x29328, x29330;
  wire x29332, x29334, x29336, x29338, x29340, x29342, x29344, x29346;
  wire x29348, x29350, x29352, x29354, x29356, x29358, x29360, x29362;
  wire x29364, x29366, x29368, x29370, x29372, x29374, x29376, x29377;
  wire x29379, x29381, x29383, x29385, x29387, x29389, x29391, x29393;
  wire x29395, x29397, x29399, x29401, x29403, x29405, x29407, x29409;
  wire x29411, x29413, x29415, x29417, x29419, x29421, x29423, x29425;
  wire x29427, x29429, x29431, x29433, x29435, x29437, x29439, x29441;
  wire x29443, x29445, x29447, x29449, x29451, x29453, x29455, x29457;
  wire x29459, x29461, x29463, x29465, x29467, x29469, x29471, x29473;
  wire x29475, x29477, x29479, x29481, x29483, x29485, x29487, x29489;
  wire x29491, x29493, x29495, x29497, x29499, x29501, x29502, x29504;
  wire x29506, x29508, x29510, x29512, x29514, x29516, x29518, x29520;
  wire x29522, x29524, x29526, x29528, x29530, x29532, x29534, x29536;
  wire x29538, x29540, x29542, x29544, x29546, x29548, x29550, x29552;
  wire x29554, x29556, x29558, x29560, x29562, x29564, x29566, x29568;
  wire x29570, x29572, x29574, x29576, x29578, x29580, x29582, x29584;
  wire x29586, x29588, x29590, x29592, x29594, x29596, x29598, x29600;
  wire x29602, x29604, x29606, x29608, x29610, x29612, x29614, x29616;
  wire x29618, x29620, x29622, x29624, x29626, x29628, x29630, x29632;
  wire x29634, x29636, x29638, x29640, x29642, x29644, x29645, x29647;
  wire x29649, x29651, x29653, x29655, x29657, x29659, x29661, x29663;
  wire x29665, x29667, x29669, x29671, x29673, x29675, x29677, x29679;
  wire x29681, x29683, x29685, x29687, x29689, x29691, x29693, x29695;
  wire x29697, x29699, x29701, x29703, x29705, x29707, x29709, x29711;
  wire x29713, x29715, x29717, x29719, x29721, x29723, x29725, x29727;
  wire x29729, x29731, x29733, x29735, x29737, x29739, x29741, x29743;
  wire x29745, x29747, x29749, x29751, x29753, x29755, x29757, x29759;
  wire x29761, x29763, x29765, x29767, x29769, x29771, x29773, x29775;
  wire x29777, x29779, x29781, x29783, x29785, x29787, x29789, x29791;
  wire x29793, x29795, x29797, x29799, x29801, x29803, x29805, x29806;
  wire x29808, x29810, x29812, x29814, x29816, x29818, x29820, x29822;
  wire x29824, x29826, x29828, x29830, x29832, x29834, x29836, x29838;
  wire x29840, x29842, x29844, x29846, x29848, x29850, x29852, x29854;
  wire x29856, x29858, x29860, x29862, x29864, x29866, x29868, x29870;
  wire x29872, x29874, x29876, x29878, x29880, x29882, x29884, x29886;
  wire x29888, x29890, x29892, x29894, x29896, x29898, x29900, x29902;
  wire x29904, x29906, x29908, x29910, x29912, x29914, x29916, x29918;
  wire x29920, x29922, x29924, x29926, x29928, x29930, x29932, x29934;
  wire x29936, x29938, x29940, x29942, x29944, x29946, x29948, x29950;
  wire x29952, x29954, x29956, x29958, x29960, x29962, x29964, x29966;
  wire x29968, x29970, x29972, x29974, x29976, x29978, x29980, x29982;
  wire x29984, x29985, x29987, x29989, x29991, x29993, x29995, x29997;
  wire x29999, x30001, x30003, x30005, x30007, x30009, x30011, x30013;
  wire x30015, x30017, x30019, x30021, x30023, x30025, x30027, x30029;
  wire x30031, x30033, x30035, x30037, x30039, x30041, x30043, x30045;
  wire x30047, x30049, x30050, x30051, x30052, x30053, x30054, x30056;
  wire x30057, x30058, x30059, x30060, x30061, x30062, x30064, x30065;
  wire x30066, x30067, x30068, x30069, x30070, x30072, x30073, x30074;
  wire x30075, x30076, x30077, x30078, x30079, x30080, x30081, x30083;
  wire x30084, x30085, x30086, x30087, x30088, x30089, x30091, x30092;
  wire x30093, x30094, x30095, x30096, x30097, x30099, x30100, x30101;
  wire x30102, x30103, x30104, x30105, x30107, x30108, x30109, x30111;
  wire x30112, x30113, x30114, x30116, x30117, x30118, x30119, x30120;
  wire x30121, x30122, x30124, x30125, x30126, x30128, x30129, x30130;
  wire x30131, x30132, x30133, x30134, x30136, x30137, x30138, x30139;
  wire x30140, x30141, x30142, x30144, x30145, x30146, x30148, x30149;
  wire x30150, x30151, x30153, x30154, x30155, x30157, x30158, x30159;
  wire x30160, x30162, x30163, x30164, x30165, x30166, x30167, x30168;
  wire x30170, x30171, x30172, x30174, x30175, x30176, x30177, x30179;
  wire x30180, x30181, x30183, x30184, x30185, x30186, x30188, x30189;
  wire x30190, x30191, x30192, x30193, x30194, x30196, x30197, x30198;
  wire x30200, x30201, x30202, x30203, x30205, x30206, x30207, x30209;
  wire x30210, x30211, x30212, x30213, x30214, x30215, x30217, x30218;
  wire x30219, x30220, x30221, x30222, x30223, x30225, x30226, x30227;
  wire x30229, x30230, x30231, x30232, x30234, x30235, x30236, x30238;
  wire x30239, x30240, x30241, x30243, x30244, x30245, x30247, x30248;
  wire x30249, x30250, x30252, x30253, x30254, x30255, x30256, x30257;
  wire x30258, x30260, x30261, x30262, x30264, x30265, x30266, x30267;
  wire x30269, x30270, x30271, x30273, x30274, x30275, x30276, x30278;
  wire x30279, x30280, x30282, x30283, x30284, x30285, x30287, x30288;
  wire x30289, x30290, x30291, x30292, x30293, x30295, x30296, x30297;
  wire x30299, x30300, x30301, x30302, x30304, x30305, x30306, x30308;
  wire x30309, x30310, x30311, x30313, x30314, x30315, x30317, x30318;
  wire x30319, x30320, x30321, x30322, x30323, x30325, x30326, x30327;
  wire x30328, x30329, x30330, x30331, x30333, x30334, x30335, x30337;
  wire x30338, x30339, x30340, x30342, x30343, x30344, x30346, x30347;
  wire x30348, x30349, x30351, x30352, x30353, x30355, x30356, x30357;
  wire x30358, x30360, x30361, x30362, x30363, x30364, x30365, x30366;
  wire x30368, x30369, x30370, x30371, x30372, x30373, x30374, x30376;
  wire x30377, x30378, x30380, x30381, x30382, x30383, x30385, x30386;
  wire x30387, x30389, x30390, x30391, x30392, x30394, x30395, x30396;
  wire x30398, x30399, x30400, x30401, x30403, x30404, x30405, x30407;
  wire x30408, x30409, x30410, x30412, x30413, x30414, x30415, x30416;
  wire x30417, x30418, x30420, x30421, x30422, x30424, x30425, x30426;
  wire x30427, x30429, x30430, x30431, x30433, x30434, x30435, x30436;
  wire x30438, x30439, x30440, x30442, x30443, x30444, x30445, x30447;
  wire x30448, x30449, x30451, x30452, x30453, x30454, x30455, x30456;
  wire x30457, x30459, x30460, x30461, x30462, x30463, x30464, x30465;
  wire x30467, x30468, x30469, x30471, x30472, x30473, x30474, x30476;
  wire x30477, x30478, x30480, x30481, x30482, x30483, x30485, x30486;
  wire x30487, x30489, x30490, x30491, x30492, x30494, x30495, x30496;
  wire x30498, x30499, x30500, x30501, x30503, x30504, x30505, x30507;
  wire x30508, x30509, x30510, x30512, x30513, x30514, x30515, x30516;
  wire x30517, x30518, x30520, x30521, x30522, x30524, x30525, x30526;
  wire x30527, x30529, x30530, x30531, x30533, x30534, x30535, x30536;
  wire x30538, x30539, x30540, x30542, x30543, x30544, x30545, x30547;
  wire x30548, x30549, x30551, x30552, x30553, x30554, x30556, x30557;
  wire x30558, x30560, x30561, x30562, x30563, x30565, x30566, x30567;
  wire x30568, x30569, x30570, x30571, x30573, x30574, x30575, x30577;
  wire x30578, x30579, x30580, x30582, x30583, x30584, x30586, x30587;
  wire x30588, x30589, x30591, x30592, x30593, x30595, x30596, x30597;
  wire x30598, x30600, x30601, x30602, x30604, x30605, x30606, x30607;
  wire x30609, x30610, x30611, x30613, x30614, x30615, x30616, x30617;
  wire x30618, x30619, x30621, x30622, x30623, x30624, x30625, x30626;
  wire x30627, x30629, x30630, x30631, x30633, x30634, x30635, x30636;
  wire x30638, x30639, x30640, x30642, x30643, x30644, x30645, x30647;
  wire x30648, x30649, x30651, x30652, x30653, x30654, x30656, x30657;
  wire x30658, x30660, x30661, x30662, x30663, x30665, x30666, x30667;
  wire x30669, x30670, x30671, x30672, x30674, x30675, x30676, x30678;
  wire x30679, x30680, x30681, x30683, x30684, x30685, x30686, x30687;
  wire x30688, x30689, x30691, x30692, x30693, x30695, x30696, x30697;
  wire x30698, x30700, x30701, x30702, x30704, x30705, x30706, x30707;
  wire x30709, x30710, x30711, x30713, x30714, x30715, x30716, x30718;
  wire x30719, x30720, x30722, x30723, x30724, x30725, x30727, x30728;
  wire x30729, x30731, x30732, x30733, x30734, x30736, x30737, x30738;
  wire x30740, x30741, x30742, x30743, x30745, x30746, x30747, x30748;
  wire x30749, x30750, x30751, x30753, x30754, x30755, x30757, x30758;
  wire x30759, x30760, x30762, x30763, x30764, x30766, x30767, x30768;
  wire x30769, x30771, x30772, x30773, x30775, x30776, x30777, x30778;
  wire x30780, x30781, x30782, x30784, x30785, x30786, x30787, x30789;
  wire x30790, x30791, x30793, x30794, x30795, x30796, x30798, x30799;
  wire x30800, x30802, x30803, x30804, x30805, x30806, x30807, x30808;
  wire x30810, x30811, x30812, x30813, x30814, x30815, x30816, x30818;
  wire x30819, x30820, x30822, x30823, x30824, x30825, x30827, x30828;
  wire x30829, x30831, x30832, x30833, x30834, x30836, x30837, x30838;
  wire x30840, x30841, x30842, x30843, x30845, x30846, x30847, x30849;
  wire x30850, x30851, x30852, x30854, x30855, x30856, x30858, x30859;
  wire x30860, x30861, x30863, x30864, x30865, x30867, x30868, x30869;
  wire x30870, x30872, x30873, x30874, x30875, x30876, x30877, x30878;
  wire x30880, x30881, x30882, x30883, x30884, x30885, x30886, x30888;
  wire x30889, x30890, x30892, x30893, x30894, x30895, x30897, x30898;
  wire x30899, x30901, x30902, x30903, x30904, x30906, x30907, x30908;
  wire x30910, x30911, x30912, x30913, x30915, x30916, x30917, x30919;
  wire x30920, x30921, x30922, x30924, x30925, x30926, x30928, x30929;
  wire x30930, x30931, x30933, x30934, x30935, x30937, x30938, x30939;
  wire x30940, x30942, x30943, x30944, x30946, x30947, x30948, x30949;
  wire x30951, x30952, x30953, x30954, x30955, x30956, x30957, x30959;
  wire x30960, x30961, x30963, x30964, x30965, x30966, x30968, x30969;
  wire x30970, x30972, x30973, x30974, x30975, x30977, x30978, x30979;
  wire x30981, x30982, x30983, x30984, x30986, x30987, x30988, x30990;
  wire x30991, x30992, x30993, x30995, x30996, x30997, x30999, x31000;
  wire x31001, x31002, x31004, x31005, x31006, x31008, x31009, x31010;
  wire x31011, x31013, x31014, x31015, x31017, x31018, x31019, x31020;
  wire x31021, x31022, x31023, x31025, x31026, x31027, x31028, x31029;
  wire x31030, x31031, x31033, x31034, x31035, x31037, x31038, x31039;
  wire x31040, x31042, x31043, x31044, x31046, x31047, x31048, x31049;
  wire x31051, x31052, x31053, x31055, x31056, x31057, x31058, x31060;
  wire x31061, x31062, x31064, x31065, x31066, x31067, x31069, x31070;
  wire x31071, x31073, x31074, x31075, x31076, x31078, x31079, x31080;
  wire x31082, x31083, x31084, x31085, x31087, x31088, x31089, x31091;
  wire x31092, x31093, x31094, x31096, x31097, x31098, x31100, x31101;
  wire x31102, x31103, x31105, x31106, x31107, x31108, x31109, x31110;
  wire x31111, x31113, x31114, x31115, x31117, x31118, x31119, x31120;
  wire x31122, x31123, x31124, x31126, x31127, x31128, x31129, x31131;
  wire x31132, x31133, x31135, x31136, x31137, x31138, x31140, x31141;
  wire x31142, x31144, x31145, x31146, x31147, x31149, x31150, x31151;
  wire x31153, x31154, x31155, x31156, x31158, x31159, x31160, x31162;
  wire x31163, x31164, x31165, x31167, x31168, x31169, x31171, x31172;
  wire x31173, x31174, x31176, x31177, x31178, x31180, x31181, x31182;
  wire x31183, x31185, x31186, x31187, x31188, x31189, x31190, x31191;
  wire x31193, x31194, x31195, x31197, x31198, x31199, x31200, x31202;
  wire x31203, x31204, x31206, x31207, x31208, x31209, x31211, x31212;
  wire x31213, x31215, x31216, x31217, x31218, x31220, x31221, x31222;
  wire x31224, x31225, x31226, x31227, x31229, x31230, x31231, x31233;
  wire x31234, x31235, x31236, x31238, x31239, x31240, x31242, x31243;
  wire x31244, x31245, x31247, x31248, x31249, x31251, x31252, x31253;
  wire x31254, x31256, x31257, x31258, x31260, x31261, x31262, x31263;
  wire x31264, x31265, x31266, x31268, x31269, x31270, x31272, x31273;
  wire x31274, x31275, x31277, x31278, x31279, x31281, x31282, x31283;
  wire x31284, x31286, x31287, x31288, x31290, x31291, x31292, x31293;
  wire x31295, x31296, x31297, x31299, x31300, x31301, x31302, x31304;
  wire x31305, x31306, x31308, x31309, x31310, x31311, x31313, x31314;
  wire x31315, x31317, x31318, x31319, x31320, x31322, x31323, x31324;
  wire x31326, x31327, x31328, x31329, x31331, x31332, x31333, x31335;
  wire x31336, x31337, x31338, x31340, x31341, x31342, x31344, x31345;
  wire x31346, x31347, x31349, x31350, x31351, x31353, x31354, x31355;
  wire x31356, x31358, x31359, x31360, x31362, x31363, x31364, x31365;
  wire x31367, x31368, x31369, x31371, x31372, x31373, x31374, x31376;
  wire x31377, x31378, x31380, x31381, x31382, x31383, x31385, x31386;
  wire x31387, x31389, x31390, x31391, x31392, x31394, x31395, x31396;
  wire x31398, x31399, x31400, x31401, x31403, x31404, x31405, x31407;
  wire x31408, x31409, x31410, x31412, x31413, x31414, x31416, x31417;
  wire x31418, x31419, x31421, x31422, x31423, x31425, x31426, x31427;
  wire x31428, x31430, x31431, x31432, x31434, x31435, x31436, x31437;
  wire x31439, x31440, x31441, x31443, x31444, x31445, x31446, x31448;
  wire x31449, x31450, x31452, x31453, x31454, x31456, x31457, x31458;
  wire x31460, x31461, x31462, x31464, x31465, x31466, x31468, x31469;
  wire x31470, x31472, x31473, x31474, x31476, x31477, x31478, x31480;
  wire x31481, x31482, x31484, x31485, x31486, x31488, x31489, x31490;
  wire x31492, x31493, x31494, x31496, x31497, x31498, x31500, x31501;
  wire x31502, x31504, x31505, x31506, x31508, x31509, x31510, x31512;
  wire x31513, x31514, x31516, x31517, x31518, x31520, x31521, x31522;
  wire x31524, x31525, x31526, x31530, x31532, x31533, x31534, x31537;
  wire x31538, x31539, x31540, x31541, x31542, x31545, x31546, x31547;
  wire x31548, x31549, x31550, x31553, x31554, x31556, x31557, x31558;
  wire x31559, x31560, x31561, x31562, x31563, x31566, x31567, x31569;
  wire x31571, x31572, x31573, x31574, x31575, x31576, x31578, x31579;
  wire x31580, x31582, x31583, x31586, x31587, x31589, x31591, x31592;
  wire x31593, x31594, x31595, x31596, x31598, x31599, x31600, x31602;
  wire x31603, x31606, x31607, x31609, x31611, x31612, x31613, x31614;
  wire x31615, x31616, x31618, x31619, x31620, x31622, x31623, x31626;
  wire x31627, x31629, x31631, x31632, x31633, x31635, x31636, x31637;
  wire x31639, x31640, x31641, x31643, x31644, x31647, x31648, x31650;
  wire x31652, x31653, x31654, x31656, x31657, x31658, x31660, x31661;
  wire x31662, x31664, x31665, x31668, x31669, x31671, x31673, x31674;
  wire x31675, x31676, x31678, x31679, x31680, x31681, x31682, x31684;
  wire x31685, x31686, x31688, x31689, x31692, x31693, x31695, x31697;
  wire x31698, x31699, x31700, x31703, x31704, x31705, x31706, x31707;
  wire x31709, x31710, x31711, x31713, x31714, x31715, x31716, x31717;
  wire x31720, x31721, x31723, x31725, x31726, x31727, x31728, x31731;
  wire x31732, x31733, x31734, x31735, x31737, x31738, x31739, x31741;
  wire x31742, x31743, x31744, x31745, x31748, x31749, x31751, x31753;
  wire x31754, x31755, x31756, x31759, x31760, x31762, x31763, x31764;
  wire x31766, x31767, x31768, x31769, x31771, x31772, x31773, x31775;
  wire x31776, x31777, x31778, x31779, x31782, x31783, x31785, x31787;
  wire x31788, x31789, x31790, x31793, x31794, x31796, x31798, x31799;
  wire x31801, x31802, x31803, x31804, x31806, x31807, x31808, x31810;
  wire x31811, x31812, x31813, x31815, x31816, x31817, x31818, x31819;
  wire x31822, x31823, x31825, x31827, x31828, x31829, x31830, x31833;
  wire x31834, x31836, x31838, x31839, x31841, x31842, x31843, x31844;
  wire x31846, x31847, x31848, x31850, x31851, x31852, x31853, x31855;
  wire x31856, x31857, x31858, x31859, x31862, x31863, x31865, x31867;
  wire x31868, x31869, x31870, x31873, x31874, x31876, x31878, x31879;
  wire x31881, x31882, x31883, x31884, x31886, x31887, x31888, x31890;
  wire x31891, x31892, x31893, x31895, x31896, x31897, x31898, x31899;
  wire x31902, x31903, x31905, x31907, x31908, x31909, x31910, x31913;
  wire x31914, x31916, x31918, x31919, x31921, x31923, x31924, x31925;
  wire x31927, x31928, x31929, x31931, x31932, x31933, x31934, x31936;
  wire x31937, x31938, x31940, x31941, x31944, x31945, x31947, x31949;
  wire x31950, x31951, x31952, x31955, x31956, x31958, x31960, x31961;
  wire x31963, x31965, x31966, x31967, x31969, x31970, x31971, x31973;
  wire x31974, x31975, x31976, x31978, x31979, x31980, x31982, x31983;
  wire x31986, x31987, x31989, x31991, x31992, x31993, x31994, x31997;
  wire x31998, x32000, x32002, x32003, x32005, x32006, x32008, x32009;
  wire x32010, x32011, x32012, x32014, x32015, x32016, x32018, x32019;
  wire x32020, x32021, x32023, x32024, x32025, x32027, x32028, x32031;
  wire x32032, x32034, x32036, x32037, x32038, x32039, x32042, x32043;
  wire x32045, x32047, x32048, x32050, x32051, x32054, x32055, x32056;
  wire x32057, x32058, x32060, x32061, x32062, x32064, x32065, x32066;
  wire x32067, x32069, x32070, x32071, x32073, x32074, x32075, x32076;
  wire x32077, x32080, x32081, x32083, x32085, x32086, x32088, x32089;
  wire x32092, x32093, x32095, x32097, x32098, x32100, x32101, x32104;
  wire x32105, x32106, x32107, x32108, x32110, x32111, x32112, x32114;
  wire x32115, x32116, x32117, x32119, x32120, x32121, x32123, x32124;
  wire x32125, x32126, x32127, x32130, x32131, x32133, x32135, x32136;
  wire x32138, x32139, x32142, x32143, x32145, x32147, x32148, x32150;
  wire x32151, x32154, x32155, x32157, x32158, x32159, x32161, x32162;
  wire x32163, x32164, x32166, x32167, x32168, x32170, x32171, x32172;
  wire x32173, x32175, x32176, x32177, x32179, x32180, x32181, x32182;
  wire x32183, x32186, x32187, x32189, x32191, x32192, x32194, x32195;
  wire x32198, x32199, x32201, x32203, x32204, x32206, x32207, x32210;
  wire x32211, x32213, x32215, x32216, x32218, x32219, x32220, x32221;
  wire x32223, x32224, x32225, x32227, x32228, x32229, x32230, x32232;
  wire x32233, x32234, x32236, x32237, x32238, x32239, x32241, x32242;
  wire x32243, x32245, x32246, x32249, x32250, x32252, x32254, x32255;
  wire x32257, x32258, x32261, x32262, x32264, x32266, x32267, x32269;
  wire x32270, x32273, x32274, x32276, x32278, x32279, x32281, x32282;
  wire x32283, x32284, x32286, x32287, x32288, x32290, x32291, x32292;
  wire x32293, x32295, x32296, x32297, x32299, x32300, x32301, x32302;
  wire x32304, x32305, x32306, x32308, x32309, x32312, x32313, x32315;
  wire x32317, x32318, x32320, x32321, x32324, x32325, x32327, x32329;
  wire x32330, x32332, x32333, x32336, x32337, x32339, x32341, x32342;
  wire x32344, x32345, x32346, x32347, x32349, x32350, x32351, x32353;
  wire x32354, x32355, x32357, x32358, x32359, x32360, x32362, x32363;
  wire x32364, x32366, x32367, x32368, x32369, x32371, x32372, x32373;
  wire x32375, x32376, x32379, x32380, x32382, x32384, x32385, x32387;
  wire x32388, x32391, x32392, x32394, x32396, x32397, x32399, x32400;
  wire x32403, x32404, x32406, x32408, x32409, x32411, x32413, x32414;
  wire x32415, x32417, x32418, x32419, x32421, x32422, x32423, x32425;
  wire x32426, x32427, x32428, x32430, x32431, x32432, x32434, x32435;
  wire x32436, x32437, x32439, x32440, x32441, x32443, x32444, x32447;
  wire x32448, x32450, x32452, x32453, x32455, x32458, x32459, x32461;
  wire x32463, x32464, x32466, x32469, x32470, x32472, x32474, x32475;
  wire x32478, x32479, x32480, x32482, x32483, x32484, x32486, x32487;
  wire x32488, x32490, x32491, x32492, x32494, x32495, x32496, x32498;
  wire x32499, x32500, x32502, x32503, x32504, x32506, x32507, x32508;
  wire x32510, x32511, x32512, x32514, x32515, x32516, x32518, x32519;
  wire x32520, x32522, x32523, x32524, x32526, x32527, x32528, x32531;
  wire x32532, x32533, x32537, x32538, x32539, x32543, x32544, x32545;
  wire x32547, x32548, x32549, x32553, x32554, x32555, x32557, x32558;
  wire x32559, x32563, x32564, x32565, x32567, x32568, x32569, x32573;
  wire x32574, x32575, x32577, x32578, x32579, x32581, x32583, x32584;
  wire x32586, x32587, x32588, x32590, x32591, x32592, x32594, x32596;
  wire x32597, x32599, x32600, x32601, x32603, x32604, x32605, x32607;
  wire x32608, x32609, x32611, x32613, x32614, x32616, x32617, x32618;
  wire x32620, x32621, x32622, x32624, x32625, x32626, x32628, x32631;
  wire x32632, x32634, x32635, x32636, x32638, x32639, x32640, x32642;
  wire x32643, x32644, x32646, x32649, x32650, x32652, x32654, x32655;
  wire x32657, x32658, x32659, x32661, x32662, x32663, x32665, x32668;
  wire x32669, x32671, x32673, x32674, x32676, x32677, x32678, x32680;
  wire x32681, x32682, x32684, x32685, x32686, x32688, x32689, x32692;
  wire x32693, x32695, x32697, x32698, x32700, x32701, x32702, x32704;
  wire x32705, x32706, x32708, x32709, x32710, x32712, x32713, x32714;
  wire x32715, x32716, x32719, x32720, x32722, x32724, x32725, x32727;
  wire x32728, x32729, x32731, x32732, x32733, x32735, x32736, x32737;
  wire x32739, x32740, x32741, x32742, x32743, x32746, x32747, x32749;
  wire x32751, x32752, x32754, x32755, x32756, x32758, x32759, x32760;
  wire x32762, x32763, x32764, x32766, x32767, x32768, x32769, x32770;
  wire x32773, x32774, x32776, x32777, x32778, x32780, x32782, x32784;
  wire x32785, x32787, x32788, x32789, x32791, x32792, x32793, x32795;
  wire x32796, x32797, x32799, x32800, x32801, x32802, x32803, x32806;
  wire x32807, x32809, x32810, x32811, x32813, x32815, x32817, x32818;
  wire x32820, x32821, x32822, x32824, x32825, x32826, x32828, x32829;
  wire x32830, x32831, x32833, x32834, x32835, x32837, x32838, x32839;
  wire x32840, x32841, x32844, x32845, x32847, x32848, x32849, x32851;
  wire x32853, x32855, x32856, x32858, x32859, x32860, x32862, x32863;
  wire x32864, x32866, x32867, x32868, x32869, x32871, x32872, x32873;
  wire x32875, x32876, x32877, x32878, x32879, x32882, x32883, x32885;
  wire x32887, x32888, x32890, x32892, x32894, x32895, x32897, x32898;
  wire x32899, x32901, x32902, x32903, x32905, x32906, x32907, x32908;
  wire x32910, x32911, x32912, x32914, x32915, x32916, x32917, x32918;
  wire x32921, x32922, x32924, x32926, x32927, x32929, x32931, x32933;
  wire x32934, x32936, x32938, x32939, x32941, x32942, x32943, x32945;
  wire x32946, x32947, x32948, x32950, x32951, x32952, x32954, x32955;
  wire x32956, x32957, x32958, x32961, x32962, x32964, x32966, x32967;
  wire x32969, x32971, x32973, x32974, x32976, x32978, x32979, x32981;
  wire x32982, x32983, x32985, x32986, x32987, x32988, x32990, x32991;
  wire x32992, x32994, x32995, x32996, x32997, x32998, x33001, x33002;
  wire x33004, x33006, x33007, x33009, x33010, x33012, x33013, x33015;
  wire x33017, x33018, x33020, x33021, x33023, x33024, x33026, x33027;
  wire x33028, x33030, x33031, x33032, x33033, x33035, x33036, x33037;
  wire x33039, x33040, x33041, x33042, x33044, x33045, x33046, x33048;
  wire x33049, x33052, x33053, x33055, x33057, x33058, x33060, x33062;
  wire x33063, x33065, x33067, x33068, x33070, x33072, x33073, x33075;
  wire x33076, x33077, x33079, x33080, x33081, x33083, x33084, x33085;
  wire x33087, x33088, x33089, x33091, x33092, x33093, x33095, x33096;
  wire x33097, x33098, x33099, x33100, x33101, x33102, x33103, x33105;
  wire x33106, x33107, x33109, x33110, x33111, x33112, x33113, x33114;
  wire x33116, x33117, x33118, x33119, x33120, x33121, x33123, x33124;
  wire x33125, x33127, x33128, x33129, x33130, x33131, x33132, x33133;
  wire x33135, x33136, x33137, x33139, x33140, x33141, x33142, x33143;
  wire x33144, x33145, x33147, x33148, x33149, x33151, x33152, x33153;
  wire x33154, x33155, x33156, x33157, x33159, x33160, x33161, x33163;
  wire x33164, x33165, x33166, x33167, x33168, x33169, x33171, x33172;
  wire x33173, x33175, x33176, x33177, x33178, x33180, x33181, x33182;
  wire x33184, x33185, x33186, x33188, x33189, x33190, x33191, x33193;
  wire x33194, x33195, x33197, x33198, x33199, x33201, x33202, x33203;
  wire x33204, x33206, x33207, x33208, x33210, x33211, x33212, x33214;
  wire x33215, x33216, x33217, x33219, x33220, x33221, x33223, x33224;
  wire x33225, x33227, x33228, x33229, x33230, x33232, x33233, x33234;
  wire x33236, x33237, x33238, x33240, x33241, x33242, x33244, x33245;
  wire x33246, x33247, x33249, x33250, x33251, x33253, x33254, x33255;
  wire x33256, x33258, x33259, x33260, x33262, x33263, x33264, x33266;
  wire x33267, x33268, x33269, x33271, x33272, x33273, x33275, x33276;
  wire x33277, x33278, x33280, x33281, x33282, x33284, x33285, x33286;
  wire x33288, x33289, x33290, x33291, x33293, x33294, x33295, x33297;
  wire x33298, x33299, x33300, x33302, x33303, x33304, x33306, x33307;
  wire x33308, x33310, x33311, x33312, x33313, x33315, x33316, x33317;
  wire x33319, x33320, x33321, x33322, x33324, x33325, x33326, x33328;
  wire x33329, x33330, x33332, x33333, x33334, x33335, x33337, x33338;
  wire x33339, x33341, x33343, x33344, x33345, x33347, x33348, x33349;
  wire x33351, x33352, x33353, x33355, x33356, x33357, x33358, x33360;
  wire x33361, x33362, x33364, x33365, x33367, x33368, x33370, x33371;
  wire x33372, x33374, x33375, x33376, x33377, x33379, x33380, x33381;
  wire x33383, x33384, x33385, x33386, x33388, x33389, x33390, x33392;
  wire x33393, x33395, x33396, x33398, x33399, x33400, x33402, x33403;
  wire x33404, x33405, x33407, x33408, x33409, x33411, x33412, x33413;
  wire x33414, x33416, x33417, x33418, x33420, x33421, x33423, x33424;
  wire x33426, x33427, x33428, x33430, x33431, x33432, x33433, x33435;
  wire x33436, x33437, x33439, x33440, x33442, x33443, x33445, x33446;
  wire x33447, x33449, x33450, x33452, x33453, x33455, x33456, x33457;
  wire x33459, x33460, x33461, x33462, x33464, x33465, x33466, x33468;
  wire x33469, x33471, x33472, x33474, x33476, x33477, x33479, x33480;
  wire x33482, x33483, x33485, x33486, x33487, x33489, x33490, x33491;
  wire x33492, x33494, x33495, x33496, x33498, x33499, x33501, x33502;
  wire x33504, x33506, x33507, x33509, x33510, x33512, x33513, x33515;
  wire x33516, x33517, x33519, x33520, x33521, x33522, x33524, x33525;
  wire x33526, x33528, x33529, x33531, x33532, x33534, x33536, x33537;
  wire x33539, x33540, x33542, x33543, x33545, x33546, x33547, x33549;
  wire x33550, x33551, x33552, x33554, x33555, x33556, x33558, x33559;
  wire x33561, x33562, x33564, x33566, x33567, x33569, x33570, x33572;
  wire x33573, x33575, x33576, x33577, x33579, x33580, x33581, x33582;
  wire x33584, x33585, x33586, x33588, x33589, x33591, x33592, x33594;
  wire x33596, x33597, x33599, x33600, x33602, x33603, x33605, x33606;
  wire x33607, x33609, x33610, x33611, x33612, x33614, x33615, x33616;
  wire x33618, x33619, x33622, x33623, x33625, x33627, x33628, x33630;
  wire x33633, x33634, x33636, x33637, x33638, x33640, x33641, x33642;
  wire x33644, x33645, x33646, x33648, x33649, x33650, x33651, x33652;
  wire x33653, x33654, x33655, x33656, x33657, x33658, x33659, x33661;
  wire x33662, x33663, x33664, x33666, x33667, x33669, x33670, x33671;
  wire x33672, x33674, x33675, x33677, x33678, x33679, x33680, x33682;
  wire x33683, x33685, x33686, x33687, x33688, x33690, x33691, x33693;
  wire x33694, x33695, x33696, x33698, x33699, x33701, x33702, x33703;
  wire x33705, x33706, x33707, x33709, x33710, x33712, x33713, x33715;
  wire x33716, x33717, x33719, x33720, x33721, x33723, x33724, x33726;
  wire x33727, x33729, x33730, x33731, x33733, x33734, x33735, x33737;
  wire x33738, x33740, x33741, x33743, x33744, x33745, x33747, x33748;
  wire x33749, x33751, x33752, x33754, x33755, x33757, x33758, x33759;
  wire x33761, x33762, x33763, x33765, x33766, x33767, x33768, x33770;
  wire x33772, x33773, x33775, x33776, x33777, x33778, x33780, x33781;
  wire x33782, x33784, x33785, x33787, x33788, x33790, x33792, x33793;
  wire x33795, x33796, x33797, x33798, x33800, x33801, x33802, x33804;
  wire x33805, x33807, x33808, x33810, x33812, x33813, x33815, x33816;
  wire x33817, x33818, x33820, x33821, x33822, x33824, x33825, x33827;
  wire x33828, x33830, x33832, x33833, x33835, x33836, x33837, x33838;
  wire x33840, x33841, x33842, x33844, x33845, x33847, x33848, x33850;
  wire x33852, x33853, x33855, x33856, x33857, x33858, x33860, x33861;
  wire x33862, x33864, x33865, x33867, x33868, x33870, x33872, x33873;
  wire x33875, x33876, x33877, x33878, x33880, x33881, x33882, x33884;
  wire x33885, x33888, x33889, x33891, x33893, x33894, x33896, x33897;
  wire x33898, x33899, x33901, x33902, x33903, x33905, x33906, x33909;
  wire x33910, x33912, x33914, x33915, x33917, x33918, x33919, x33920;
  wire x33922, x33923, x33924, x33926, x33927, x33930, x33931, x33933;
  wire x33935, x33936, x33938, x33939, x33940, x33941, x33943, x33944;
  wire x33945, x33947, x33948, x33951, x33952, x33954, x33956, x33957;
  wire x33959, x33960, x33961, x33962, x33964, x33965, x33966, x33968;
  wire x33969, x33972, x33973, x33975, x33977, x33978, x33980, x33981;
  wire x33982, x33983, x33985, x33986, x33987, x33989, x33990, x33993;
  wire x33994, x33996, x33998, x33999, x34001, x34002, x34003, x34004;
  wire x34006, x34007, x34008, x34010, x34011, x34014, x34015, x34017;
  wire x34019, x34020, x34022, x34023, x34024, x34025, x34027, x34028;
  wire x34029, x34031, x34032, x34035, x34036, x34038, x34040, x34041;
  wire x34043, x34044, x34045, x34046, x34048, x34049, x34050, x34052;
  wire x34053, x34056, x34057, x34059, x34061, x34062, x34064, x34065;
  wire x34066, x34068, x34069, x34070, x34072, x34073, x34074, x34075;
  wire x34076, x34077, x34079, x34080, x34081, x34083, x34084, x34085;
  wire x34087, x34088, x34089, x34091, x34092, x34093, x34094, x34096;
  wire x34097, x34098, x34100, x34101, x34102, x34103, x34105, x34106;
  wire x34107, x34109, x34110, x34111, x34112, x34114, x34115, x34116;
  wire x34118, x34119, x34120, x34121, x34123, x34124, x34125, x34127;
  wire x34128, x34129, x34130, x34133, x34135, x34136, x34138, x34139;
  wire x34140, x34142, x34143, x34144, x34145, x34148, x34150, x34151;
  wire x34153, x34154, x34155, x34157, x34158, x34159, x34160, x34163;
  wire x34165, x34166, x34168, x34169, x34170, x34172, x34173, x34174;
  wire x34175, x34178, x34180, x34181, x34183, x34184, x34185, x34187;
  wire x34188, x34189, x34190, x34193, x34195, x34196, x34198, x34199;
  wire x34200, x34202, x34203, x34204, x34205, x34208, x34211, x34212;
  wire x34214, x34215, x34216, x34218, x34219, x34220, x34221, x34224;
  wire x34227, x34228, x34230, x34231, x34232, x34234, x34235, x34236;
  wire x34237, x34240, x34243, x34244, x34246, x34247, x34248, x34250;
  wire x34251, x34252, x34253, x34256, x34259, x34260, x34262, x34263;
  wire x34264, x34266, x34267, x34268, x34269, x34272, x34275, x34276;
  wire x34278, x34279, x34280, x34282, x34283, x34284, x34285, x34288;
  wire x34291, x34292, x34294, x34295, x34296, x34298, x34299, x34300;
  wire x34301, x34304, x34307, x34308, x34310, x34311, x34312, x34314;
  wire x34315, x34316, x34317, x34320, x34323, x34324, x34326, x34327;
  wire x34328, x34330, x34331, x34332, x34333, x34336, x34339, x34340;
  wire x34342, x34343, x34344, x34346, x34347, x34348, x34349, x34352;
  wire x34355, x34356, x34358, x34359, x34360, x34362, x34363, x34364;
  wire x34365, x34368, x34371, x34372, x34374, x34375, x34376, x34378;
  wire x34379, x34380, x34381, x34384, x34387, x34388, x34390, x34391;
  wire x34392, x34394, x34395, x34396, x34397, x34400, x34403, x34404;
  wire x34406, x34407, x34408, x34410, x34411, x34412, x34413, x34416;
  wire x34419, x34420, x34422, x34423, x34424, x34426, x34427, x34428;
  wire x34430, x34431, x34432, x34433, x34434, x34435, x34436, x34437;
  wire x34438, x34440, x34441, x34442, x34445, x34446, x34447, x34450;
  wire x34451, x34452, x34455, x34456, x34457, x34460, x34461, x34462;
  wire x34464, x34466, x34467, x34469, x34470, x34471, x34473, x34474;
  wire x34476, x34477, x34479, x34480, x34481, x34483, x34484, x34486;
  wire x34487, x34489, x34490, x34491, x34493, x34494, x34496, x34497;
  wire x34499, x34500, x34501, x34503, x34504, x34506, x34507, x34509;
  wire x34510, x34511, x34513, x34514, x34516, x34517, x34519, x34520;
  wire x34521, x34523, x34524, x34526, x34527, x34529, x34530, x34531;
  wire x34533, x34534, x34536, x34537, x34539, x34540, x34541, x34543;
  wire x34544, x34546, x34547, x34549, x34550, x34551, x34553, x34554;
  wire x34556, x34557, x34559, x34560, x34561, x34563, x34564, x34566;
  wire x34567, x34569, x34570, x34571, x34573, x34574, x34576, x34577;
  wire x34579, x34580, x34581, x34583, x34584, x34586, x34587, x34589;
  wire x34590, x34591, x34593, x34594, x34596, x34597, x34599, x34600;
  wire x34601, x34603, x34604, x34606, x34607, x34609, x34610, x34611;
  wire x34613, x34614, x34616, x34617, x34619, x34620, x34621, x34623;
  wire x34624, x34626, x34627, x34629, x34630, x34631, x34633, x34634;
  wire x34636, x34637, x34639, x34640, x34641, x34643, x34644, x34646;
  wire x34647, x34649, x34650, x34651, x34653, x34654, x34655, x34657;
  wire x34658, x34659, x34660, x34661, x34662, x34663, x34665, x34666;
  wire x34667, x34669, x34670, x34671, x34673, x34674, x34675, x34677;
  wire x34678, x34679, x34680, x34682, x34683, x34684, x34686, x34687;
  wire x34688, x34689, x34691, x34692, x34693, x34695, x34696, x34697;
  wire x34698, x34700, x34701, x34702, x34704, x34705, x34706, x34707;
  wire x34709, x34710, x34711, x34713, x34714, x34715, x34716, x34718;
  wire x34719, x34720, x34722, x34723, x34724, x34725, x34727, x34728;
  wire x34729, x34731, x34732, x34734, x34735, x34737, x34738, x34739;
  wire x34741, x34742, x34744, x34745, x34747, x34748, x34749, x34751;
  wire x34752, x34754, x34755, x34757, x34758, x34759, x34761, x34762;
  wire x34764, x34765, x34767, x34768, x34769, x34771, x34772, x34774;
  wire x34775, x34777, x34778, x34779, x34781, x34782, x34784, x34785;
  wire x34787, x34788, x34789, x34791, x34792, x34794, x34795, x34797;
  wire x34798, x34799, x34801, x34802, x34804, x34805, x34807, x34808;
  wire x34809, x34811, x34812, x34814, x34815, x34817, x34818, x34819;
  wire x34821, x34822, x34824, x34825, x34827, x34828, x34829, x34831;
  wire x34832, x34834, x34835, x34837, x34838, x34839, x34841, x34842;
  wire x34844, x34845, x34847, x34848, x34849, x34851, x34852, x34854;
  wire x34855, x34857, x34858, x34859, x34861, x34862, x34864, x34865;
  wire x34867, x34868, x34869, x34871, x34872, x34874, x34875, x34877;
  wire x34878, x34879, x34881, x34882, x34884, x34885, x34887, x34888;
  wire x34889, x34891, x34892, x34894, x34895, x34897, x34898, x34899;
  wire x34901, x34902, x34904, x34905, x34907, x34908, x34909, x34911;
  wire x34913, x34914, x34915, x34916, x34917, x34919, x34920, x34921;
  wire x34923, x34925, x34926, x34928, x34930, x34931, x34933, x34935;
  wire x34936, x34938, x34940, x34941, x34943, x34945, x34946, x34948;
  wire x34950, x34951, x34953, x34955, x34956, x34958, x34960, x34961;
  wire x34963, x34965, x34966, x34968, x34970, x34971, x34973, x34975;
  wire x34976, x34978, x34980, x34981, x34983, x34985, x34986, x34988;
  wire x34990, x34991, x34993, x34995, x34996, x34998, x35000, x35001;
  wire x35003, x35005, x35006, x35008, x35010, x35011, x35013, x35015;
  wire x35016, x35018, x35020, x35021, x35023, x35025, x35026, x35028;
  wire x35030, x35031, x35033, x35035, x35036, x35038, x35040, x35041;
  wire x35068, x35069, x35070, x35071, x35072, x35074, x35075, x35076;
  wire x35078, x35079, x35080, x35082, x35083, x35084, x35086, x35087;
  wire x35088, x35090, x35091, x35092, x35094, x35095, x35096, x35098;
  wire x35099, x35100, x35102, x35103, x35104, x35106, x35107, x35108;
  wire x35110, x35111, x35112, x35114, x35115, x35116, x35118, x35119;
  wire x35120, x35122, x35123, x35124, x35126, x35127, x35128, x35130;
  wire x35131, x35132, x35134, x35135, x35136, x35138, x35139, x35140;
  wire x35142, x35143, x35144, x35146, x35147, x35148, x35150, x35151;
  wire x35152, x35154, x35155, x35156, x35158, x35159, x35160, x35162;
  wire x35163, x35164, x35167, x35169, x35170, x35172, x35173, x35175;
  wire x35176, x35178, x35180, x35181, x35183, x35185, x35186, x35188;
  wire x35190, x35191, x35193, x35195, x35196, x35198, x35200, x35201;
  wire x35203, x35205, x35206, x35208, x35210, x35211, x35213, x35215;
  wire x35216, x35218, x35220, x35221, x35223, x35225, x35226, x35228;
  wire x35230, x35231, x35233, x35235, x35236, x35238, x35240, x35241;
  wire x35243, x35245, x35246, x35248, x35250, x35251, x35253, x35255;
  wire x35256, x35258, x35260, x35261, x35263, x35265, x35266, x35268;
  wire x35270, x35271, x35273, x35275, x35276, x35278, x35280, x35281;
  wire x35285, x35287, x35288, x35290, x35291, x35293, x35294, x35296;
  wire x35297, x35299, x35300, x35302, x35304, x35305, x35307, x35309;
  wire x35310, x35312, x35314, x35315, x35317, x35319, x35320, x35322;
  wire x35324, x35325, x35327, x35329, x35330, x35332, x35334, x35335;
  wire x35337, x35339, x35340, x35342, x35344, x35345, x35347, x35349;
  wire x35350, x35352, x35354, x35355, x35357, x35359, x35360, x35362;
  wire x35364, x35365, x35367, x35369, x35370, x35372, x35374, x35375;
  wire x35377, x35379, x35380, x35382, x35384, x35385, x35391, x35393;
  wire x35394, x35396, x35397, x35399, x35400, x35402, x35403, x35405;
  wire x35406, x35408, x35409, x35411, x35412, x35414, x35415, x35417;
  wire x35418, x35420, x35422, x35423, x35425, x35427, x35428, x35430;
  wire x35432, x35433, x35435, x35437, x35438, x35440, x35442, x35443;
  wire x35445, x35447, x35448, x35450, x35452, x35453, x35455, x35457;
  wire x35458, x35460, x35462, x35463, x35471, x35473, x35474, x35476;
  wire x35477, x35479, x35480, x35482, x35483, x35485, x35486, x35488;
  wire x35489, x35491, x35492, x35494, x35495, x35497, x35498, x35500;
  wire x35501, x35502, x35504, x35505, x35506, x35508, x35509, x35510;
  wire x35512, x35513, x35514, x35516, x35517, x35518, x35520, x35521;
  wire x35522, x35524, x35525, x35526, x35528, x35529, x35530, x35532;
  wire x35534, x35535, x35537, x35539, x35540, x35542, x35543, x35544;
  wire x35546, x35547, x35548, x35550, x35551, x35552, x35554, x35555;
  wire x35556, x35558, x35559, x35560, x35562, x35563, x35564, x35566;
  wire x35568, x35569, x35571, x35573, x35574, x35576, x35578, x35579;
  wire x35581, x35583, x35584, x35586, x35588, x35589, x35591, x35593;
  wire x35594, x35596, x35598, x35599, x35601, x35603, x35604, x35606;
  wire x35608, x35609, x35611, x35613, x35614, x35616, x35618, x35620;
  wire x35622, x35624, x35626, x35628, x35630, x35632, x35634, x35636;
  wire x35638, x35640, x35642, x35644, x35646, x35648, x35650, x35652;
  wire x35654, x35656, x35658, x35660, x35662, x35664, x35666, x35668;
  wire x35670, x35672, x35674, x35676, x35677, x35679, x35681, x35683;
  wire x35685, x35687, x35689, x35691, x35693, x35695, x35697, x35699;
  wire x35701, x35703, x35705, x35707, x35709, x35711, x35713, x35715;
  wire x35717, x35719, x35721, x35723, x35725, x35727, x35729, x35731;
  wire x35733, x35734, x35735, x35736, x35738, x35740, x35742, x35744;
  wire x35746, x35748, x35750, x35752, x35754, x35756, x35758, x35760;
  wire x35762, x35764, x35766, x35768, x35770, x35772, x35774, x35776;
  wire x35778, x35780, x35782, x35784, x35785, x35786, x35787, x35788;
  wire x35789, x35790, x35791, x35792, x35794, x35796, x35798, x35800;
  wire x35802, x35804, x35806, x35808, x35810, x35812, x35814, x35816;
  wire x35818, x35820, x35822, x35823, x35824, x35825, x35826, x35827;
  wire x35828, x35829, x35830, x35831, x35832, x35833, x35834, x35835;
  wire x35836, x35837, x35838, x35840, x35841, x35842, x35844, x35845;
  wire x35846, x35848, x35849, x35850, x35852, x35853, x35854, x35856;
  wire x35857, x35858, x35860, x35861, x35862, x35864, x35865, x35866;
  wire x35868, x35869, x35870, x35872, x35873, x35874, x35876, x35877;
  wire x35878, x35880, x35881, x35882, x35884, x35885, x35886, x35888;
  wire x35889, x35890, x35892, x35893, x35894, x35896, x35897, x35898;
  wire x35900, x35901, x35902, x35904, x35905, x35906, x35908, x35909;
  wire x35910, x35912, x35913, x35914, x35916, x35917, x35918, x35920;
  wire x35921, x35922, x35924, x35925, x35926, x35928, x35929, x35930;
  wire x35932, x35933, x35934, x35936, x35937, x35938, x35940, x35941;
  wire x35942, x35944, x35945, x35946, x35948, x35949, x35950, x35952;
  wire x35953, x35954, x35956, x35957, x35958, x35961, x35963, x35965;
  wire x35967, x35969, x35971, x35973, x35975, x35977, x35979, x35981;
  wire x35983, x35985, x35987, x35989, x35991, x35993, x35994, x35995;
  wire x35996, x35997, x35998, x35999, x36000, x36001, x36002, x36003;
  wire x36004, x36005, x36006, x36007, x36008, x36009, x36010, x36011;
  wire x36012, x36013, x36014, x36015, x36016, x36017, x36018, x36019;
  wire x36020, x36021, x36022, x36023, x36024, x36025, x36027, x36029;
  wire x36031, x36033, x36035, x36037, x36039, x36041, x36043, x36045;
  wire x36047, x36049, x36051, x36053, x36055, x36057, x36059, x36061;
  wire x36063, x36065, x36067, x36069, x36071, x36073, x36075, x36077;
  wire x36079, x36081, x36083, x36085, x36087, x36089, x36090, x36091;
  wire x36092, x36093, x36094, x36095, x36096, x36097, x36098, x36099;
  wire x36100, x36101, x36102, x36103, x36104, x36105, x36106, x36107;
  wire x36108, x36109, x36110, x36111, x36112, x36113, x36114, x36115;
  wire x36116, x36117, x36118, x36119, x36120, x36121, x36122, x36123;
  wire x36124, x36125, x36126, x36127, x36128, x36129, x36130, x36131;
  wire x36132, x36133, x36134, x36135, x36136, x36137, x36138, x36139;
  wire x36140, x36141, x36142, x36143, x36144, x36145, x36146, x36147;
  wire x36148, x36149, x36150, x36151, x36152, x36153, x36154, x36155;
  wire x36156, x36157, x36158, x36159, x36160, x36161, x36162, x36163;
  wire x36164, x36165, x36166, x36167, x36168, x36169, x36170, x36171;
  wire x36172, x36173, x36174, x36175, x36176, x36177, x36178, x36179;
  wire x36180, x36181, x36182, x36183, x36184, x36185, x36186, x36187;
  wire x36188, x36189, x36190, x36191, x36192, x36193, x36194, x36195;
  wire x36196, x36197, x36198, x36199, x36200, x36201, x36202, x36203;
  wire x36204, x36205, x36206, x36207, x36208, x36209, x36210, x36211;
  wire x36212, x36213, x36214, x36215, x36216, x36217, x36218, x36219;
  wire x36220, x36221, x36222, x36223, x36224, x36225, x36226, x36227;
  wire x36228, x36229, x36230, x36231, x36232, x36233, x36234, x36235;
  wire x36236, x36237, x36238, x36239, x36240, x36241, x36242, x36243;
  wire x36244, x36245, x36246, x36247, x36248, x36249, x36250, x36251;
  wire x36252, x36253, x36254, x36255, x36256, x36257, x36258, x36259;
  wire x36260, x36261, x36262, x36263, x36264, x36265, x36266, x36267;
  wire x36268, x36269, x36270, x36271, x36272, x36273, x36274, x36275;
  wire x36276, x36277, x36278, x36279, x36280, x36281, x36282, x36283;
  wire x36284, x36285, x36286, x36287, x36288, x36289, x36290, x36291;
  wire x36292, x36293, x36294, x36295, x36296, x36297, x36298, x36299;
  wire x36300, x36301, x36302, x36303, x36304, x36305, x36306, x36307;
  wire x36308, x36309, x36310, x36311, x36312, x36313, x36314, x36315;
  wire x36316, x36317, x36318, x36319, x36320, x36321, x36322, x36323;
  wire x36324, x36325, x36326, x36327, x36328, x36329, x36330, x36331;
  wire x36332, x36333, x36334, x36335, x36336, x36337, x36338, x36339;
  wire x36340, x36341, x36342, x36343, x36344, x36345, x36346, x36347;
  wire x36348, x36349, x36350, x36351, x36352, x36353, x36354, x36355;
  wire x36356, x36357, x36358, x36359, x36360, x36361, x36362, x36363;
  wire x36364, x36365, x36366, x36367, x36368, x36369, x36370, x36371;
  wire x36372, x36373, x36374, x36375, x36376, x36377, x36378, x36379;
  wire x36380, x36381, x36382, x36383, x36384, x36385, x36386, x36387;
  wire x36388, x36389, x36390, x36391, x36392, x36393, x36394, x36395;
  wire x36396, x36397, x36398, x36399, x36400, x36401, x36402, x36403;
  wire x36404, x36405, x36406, x36407, x36408, x36409, x36410, x36411;
  wire x36412, x36413, x36414, x36415, x36416, x36417, x36418, x36419;
  wire x36420, x36421, x36422, x36423, x36424, x36425, x36426, x36427;
  wire x36428, x36429, x36430, x36431, x36432, x36433, x36434, x36435;
  wire x36436, x36437, x36438, x36439, x36440, x36441, x36442, x36443;
  wire x36444, x36445, x36446, x36447, x36448, x36449, x36450, x36451;
  wire x36452, x36453, x36454, x36455, x36456, x36457, x36458, x36459;
  wire x36460, x36461, x36462, x36463, x36464, x36465, x36466, x36467;
  wire x36468, x36469, x36470, x36471, x36472, x36473, x36474, x36475;
  wire x36476, x36477, x36478, x36479, x36480, x36481, x36482, x36483;
  wire x36484, x36485, x36486, x36487, x36488, x36489, x36490, x36491;
  wire x36492, x36493, x36494, x36495, x36496, x36497, x36498, x36499;
  wire x36500, x36501, x36502, x36503, x36504, x36505, x36506, x36507;
  wire x36508, x36509, x36510, x36511, x36512, x36513, x36514, x36515;
  wire x36516, x36517, x36518, x36519, x36520, x36521, x36522, x36523;
  wire x36524, x36525, x36526, x36527, x36528, x36529, x36530, x36531;
  wire x36532, x36533, x36534, x36535, x36536, x36537, x36538, x36539;
  wire x36540, x36541, x36542, x36543, x36544, x36545, x36546, x36547;
  wire x36548, x36549, x36550, x36551, x36552, x36553, x36554, x36555;
  wire x36556, x36557, x36558, x36559, x36560, x36561, x36562, x36563;
  wire x36564, x36565, x36566, x36567, x36568, x36569, x36570, x36571;
  wire x36572, x36573, x36574, x36575, x36576, x36577, x36578, x36579;
  wire x36580, x36581, x36582, x36583, x36584, x36585, x36586, x36587;
  wire x36588, x36589, x36590, x36591, x36592, x36593, x36594, x36595;
  wire x36596, x36597, x36598, x36599, x36600, x36601, x36602, x36603;
  wire x36604, x36605, x36606, x36607, x36608, x36609, x36610, x36611;
  wire x36612, x36613, x36614, x36615, x36616, x36617, x36618, x36619;
  wire x36620, x36621, x36622, x36623, x36624, x36625, x36626, x36627;
  wire x36628, x36629, x36630, x36631, x36632, x36633, x36634, x36635;
  wire x36636, x36637, x36638, x36639, x36640, x36641, x36642, x36643;
  wire x36644, x36645, x36646, x36647, x36648, x36649, x36650, x36651;
  wire x36652, x36653, x36654, x36655, x36656, x36657, x36658, x36659;
  wire x36660, x36661, x36662, x36663, x36664, x36665, x36666, x36667;
  wire x36668, x36669, x36670, x36671, x36672, x36673, x36674, x36675;
  wire x36676, x36677, x36678, x36679, x36680, x36681, x36682, x36683;
  wire x36684, x36685, x36686, x36687, x36688, x36689, x36690, x36691;
  wire x36692, x36693, x36694, x36695, x36696, x36697, x36698, x36699;
  wire x36700, x36701, x36702, x36703, x36704, x36705, x36706, x36707;
  wire x36708, x36709, x36710, x36711, x36712, x36713, x36714, x36715;
  wire x36716, x36717, x36718, x36719, x36720, x36721, x36722, x36723;
  wire x36724, x36725, x36726, x36727, x36728, x36729, x36730, x36731;
  wire x36732, x36733, x36734, x36735, x36736, x36737, x36738, x36739;
  wire x36740, x36741, x36742, x36743, x36744, x36745, x36746, x36747;
  wire x36748, x36749, x36750, x36751, x36752, x36753, x36754, x36755;
  wire x36756, x36757, x36758, x36759, x36760, x36761, x36762, x36763;
  wire x36764, x36765, x36766, x36767, x36768, x36769, x36770, x36771;
  wire x36772, x36773, x36774, x36775, x36776, x36777, x36778, x36779;
  wire x36780, x36781, x36782, x36783, x36784, x36785, x36786, x36787;
  wire x36788, x36789, x36790, x36791, x36792, x36793, x36794, x36795;
  wire x36796, x36797, x36798, x36799, x36800, x36801, x36802, x36803;
  wire x36804, x36805, x36806, x36807, x36808, x36809, x36810, x36811;
  wire x36812, x36813, x36814, x36815, x36816, x36817, x36818, x36819;
  wire x36820, x36821, x36822, x36823, x36824, x36825, x36826, x36827;
  wire x36828, x36829, x36830, x36831, x36832, x36833, x36834, x36835;
  wire x36836, x36837, x36838, x36839, x36840, x36841, x36842, x36843;
  wire x36844, x36845, x36846, x36847, x36848, x36849, x36850, x36851;
  wire x36852, x36853, x36854, x36855, x36856, x36857, x36858, x36859;
  wire x36860, x36861, x36862, x36863, x36864, x36865, x36866, x36867;
  wire x36868, x36869, x36870, x36871, x36872, x36873, x36874, x36875;
  wire x36876, x36877, x36878, x36879, x36880, x36881, x36882, x36883;
  wire x36884, x36885, x36886, x36887, x36888, x36889, x36890, x36891;
  wire x36892, x36893, x36894, x36895, x36896, x36897, x36898, x36899;
  wire x36900, x36901, x36902, x36903, x36904, x36905, x36906, x36907;
  wire x36908, x36909, x36910, x36911, x36912, x36913, x36914, x36915;
  wire x36916, x36917, x36918, x36919, x36920, x36921, x36922, x36923;
  wire x36924, x36925, x36926, x36927, x36928, x36929, x36930, x36931;
  wire x36932, x36933, x36934, x36935, x36936, x36937, x36938, x36939;
  wire x36940, x36941, x36942, x36943, x36944, x36945, x36946, x36947;
  wire x36948, x36949, x36950, x36951, x36952, x36953, x36954, x36955;
  wire x36956, x36957, x36958, x36959, x36960, x36961, x36962, x36963;
  wire x36964, x36965, x36966, x36967, x36968, x36969, x36970, x36971;
  wire x36972, x36973, x36974, x36975, x36976, x36977, x36978, x36979;
  wire x36980, x36981, x36982, x36983, x36984, x36985, x36986, x36987;
  wire x36988, x36989, x36990, x36991, x36992, x36993, x36994, x36995;
  wire x36996, x36997, x36998, x36999, x37000, x37001, x37002, x37003;
  wire x37004, x37005, x37006, x37007, x37008, x37009, x37010, x37011;
  wire x37012, x37013, x37014, x37015, x37016, x37017, x37018, x37019;
  wire x37020, x37021, x37022, x37023, x37024, x37025, x37026, x37027;
  wire x37028, x37029, x37030, x37031, x37032, x37033, x37034, x37035;
  wire x37036, x37037, x37038, x37039, x37040, x37041, x37042, x37043;
  wire x37044, x37045, x37046, x37047, x37048, x37049, x37050, x37051;
  wire x37052, x37053, x37054, x37055, x37056, x37057, x37058, x37059;
  wire x37060, x37061, x37062, x37063, x37064, x37065, x37066, x37067;
  wire x37068, x37069, x37070, x37071, x37072, x37073, x37074, x37075;
  wire x37076, x37077, x37078, x37079, x37080, x37081, x37082, x37083;
  wire x37084, x37085, x37086, x37087, x37088, x37089, x37090, x37091;
  wire x37092, x37093, x37094, x37095, x37096, x37097, x37098, x37099;
  wire x37100, x37101, x37102, x37103, x37104, x37105, x37106, x37107;
  wire x37108, x37109, x37110, x37111, x37112, x37113, x37114, x37115;
  wire x37116, x37117, x37118, x37119, x37120, x37121, x37122, x37123;
  wire x37124, x37125, x37126, x37127, x37128, x37129, x37130, x37131;
  wire x37132, x37133, x37134, x37135, x37136, x37137, x37138, x37139;
  wire x37140, x37141, x37142, x37143, x37144, x37145, x37146, x37147;
  wire x37148, x37149, x37150, x37151, x37152, x37153, x37154, x37155;
  wire x37156, x37157, x37158, x37159, x37160, x37161, x37162, x37163;
  wire x37164, x37165, x37166, x37167, x37168, x37169, x37170, x37171;
  wire x37172, x37173, x37174, x37175, x37176, x37177, x37178, x37179;
  wire x37180, x37181, x37182, x37183, x37184, x37185, x37186, x37187;
  wire x37188, x37189, x37190, x37191, x37192, x37193, x37194, x37195;
  wire x37196, x37197, x37198, x37199, x37200, x37201, x37202, x37203;
  wire x37204, x37205, x37206, x37207, x37208, x37209, x37210, x37211;
  wire x37212, x37213, x37214, x37215, x37216, x37217, x37218, x37219;
  wire x37220, x37221, x37222, x37223, x37224, x37225, x37226, x37227;
  wire x37228, x37229, x37230, x37231, x37232, x37233, x37234, x37235;
  wire x37236, x37237, x37238, x37239, x37240, x37241, x37242, x37243;
  wire x37244, x37245, x37246, x37247, x37248, x37249, x37250, x37251;
  wire x37252, x37253, x37254, x37255, x37256, x37257, x37258, x37259;
  wire x37260, x37261, x37262, x37263, x37264, x37265, x37266, x37267;
  wire x37268, x37269, x37270, x37271, x37272, x37273, x37274, x37275;
  wire x37276, x37277, x37278, x37279, x37280, x37281, x37282, x37283;
  wire x37284, x37285, x37286, x37287, x37288, x37289, x37290, x37291;
  wire x37292, x37293, x37294, x37295, x37296, x37297, x37298, x37299;
  wire x37300, x37301, x37302, x37303, x37304, x37305, x37306, x37307;
  wire x37308, x37309, x37310, x37311, x37312, x37313, x37314, x37315;
  wire x37316, x37317, x37318, x37319, x37320, x37321, x37322, x37323;
  wire x37324, x37325, x37326, x37327, x37328, x37329, x37330, x37331;
  wire x37332, x37333, x37334, x37335, x37336, x37337, x37338, x37339;
  wire x37340, x37341, x37342, x37343, x37344, x37345, x37346, x37347;
  wire x37348, x37349, x37350, x37351, x37352, x37353, x37354, x37355;
  wire x37356, x37357, x37358, x37359, x37360, x37361, x37362, x37363;
  wire x37364, x37365, x37366, x37367, x37368, x37369, x37370, x37371;
  wire x37372, x37373, x37374, x37375, x37376, x37377, x37378, x37379;
  wire x37380, x37381, x37382, x37383, x37384, x37385, x37386, x37387;
  wire x37388, x37389, x37390, x37391, x37392, x37393, x37394, x37395;
  wire x37396, x37397, x37398, x37399, x37400, x37401, x37402, x37403;
  wire x37404, x37405, x37406, x37407, x37408, x37409, x37410, x37411;
  wire x37412, x37413, x37414, x37415, x37416, x37417, x37418, x37419;
  wire x37420, x37421, x37422, x37423, x37424, x37425, x37426, x37427;
  wire x37428, x37429, x37430, x37431, x37432, x37433, x37434, x37435;
  wire x37436, x37437, x37438, x37439, x37440, x37441, x37442, x37443;
  wire x37444, x37445, x37446, x37447, x37448, x37449, x37450, x37451;
  wire x37452, x37453, x37454, x37455, x37456, x37457, x37458, x37459;
  wire x37460, x37461, x37462, x37463, x37464, x37465, x37466, x37467;
  wire x37468, x37469, x37470, x37471, x37472, x37473, x37474, x37475;
  wire x37476, x37477, x37478, x37479, x37480, x37481, x37482, x37483;
  wire x37484, x37485, x37486, x37487, x37488, x37489, x37490, x37491;
  wire x37492, x37493, x37494, x37495, x37496, x37497, x37498, x37499;
  wire x37500, x37501, x37502, x37503, x37504, x37505, x37506, x37507;
  wire x37508, x37509, x37510, x37511, x37512, x37513, x37514, x37515;
  wire x37516, x37517, x37518, x37519, x37520, x37521, x37522, x37523;
  wire x37524, x37525, x37526, x37527, x37528, x37529, x37530, x37531;
  wire x37532, x37533, x37534, x37535, x37536, x37537, x37538, x37539;
  wire x37540, x37541, x37542, x37543, x37544, x37545, x37546, x37547;
  wire x37548, x37549, x37550, x37551, x37552, x37553, x37554, x37555;
  wire x37556, x37557, x37558, x37559, x37560, x37561, x37562, x37563;
  wire x37564, x37565, x37566, x37567, x37568, x37569, x37570, x37571;
  wire x37572, x37573, x37574, x37575, x37576, x37577, x37578, x37579;
  wire x37580, x37581, x37582, x37583, x37584, x37585, x37586, x37587;
  wire x37588, x37589, x37590, x37591, x37592, x37593, x37594, x37595;
  wire x37596, x37597, x37598, x37599, x37600, x37601, x37602, x37603;
  wire x37604, x37605, x37606, x37607, x37608, x37609, x37610, x37611;
  wire x37612, x37613, x37614, x37615, x37616, x37617, x37618, x37619;
  wire x37620, x37621, x37622, x37623, x37624, x37625, x37626, x37627;
  wire x37628, x37629, x37630, x37631, x37632, x37633, x37634, x37635;
  wire x37636, x37637, x37638, x37639, x37640, x37641, x37642, x37643;
  wire x37644, x37645, x37646, x37647, x37648, x37649, x37650, x37651;
  wire x37652, x37653, x37654, x37655, x37656, x37657, x37658, x37659;
  wire x37660, x37661, x37662, x37663, x37664, x37665, x37666, x37667;
  wire x37668, x37669, x37670, x37671, x37672, x37673, x37674, x37675;
  wire x37676, x37677, x37678, x37679, x37680, x37681, x37682, x37683;
  wire x37684, x37685, x37686, x37687, x37688, x37689, x37690, x37691;
  wire x37692, x37693, x37694, x37695, x37696, x37697, x37698, x37699;
  wire x37700, x37701, x37702, x37703, x37704, x37705, x37706, x37707;
  wire x37708, x37709, x37710, x37711, x37712, x37713, x37714, x37715;
  wire x37716, x37717, x37718, x37719, x37720, x37721, x37722, x37723;
  wire x37724, x37725, x37726, x37727, x37728, x37729, x37730, x37731;
  wire x37732, x37733, x37734, x37735, x37736, x37737, x37738, x37739;
  wire x37740, x37741, x37742, x37743, x37744, x37745, x37746, x37747;
  wire x37748, x37749, x37750, x37751, x37752, x37753, x37754, x37755;
  wire x37756, x37757, x37758, x37759, x37760, x37761, x37762, x37763;
  wire x37764, x37765, x37766, x37767, x37768, x37769, x37770, x37771;
  wire x37772, x37773, x37774, x37775, x37776, x37777, x37778, x37779;
  wire x37780, x37781, x37782, x37783, x37784, x37785, x37786, x37787;
  wire x37788, x37789, x37790, x37791, x37792, x37793, x37794, x37795;
  wire x37796, x37797, x37798, x37799, x37800, x37801, x37802, x37803;
  wire x37804, x37805, x37806, x37807, x37808, x37809, x37810, x37811;
  wire x37812, x37813, x37814, x37815, x37816, x37817, x37818, x37819;
  wire x37820, x37821, x37822, x37823, x37824, x37825, x37826, x37827;
  wire x37828, x37829, x37830, x37831, x37832, x37833, x37834, x37835;
  wire x37836, x37837, x37838, x37839, x37840, x37841, x37842, x37843;
  wire x37844, x37845, x37846, x37847, x37848, x37849, x37850, x37851;
  wire x37852, x37853, x37854, x37855, x37856, x37857, x37858, x37859;
  wire x37860, x37861, x37862, x37863, x37864, x37865, x37866, x37867;
  wire x37868, x37869, x37870, x37871, x37872, x37873, x37874, x37875;
  wire x37876, x37877, x37878, x37879, x37880, x37881, x37882, x37883;
  wire x37884, x37885, x37886, x37887, x37888, x37889, x37890, x37891;
  wire x37892, x37893, x37894, x37895, x37896, x37897, x37898, x37899;
  wire x37900, x37901, x37902, x37903, x37904, x37905, x37906, x37907;
  wire x37908, x37909, x37910, x37911, x37912, x37913, x37914, x37915;
  wire x37916, x37917, x37918, x37919, x37920, x37921, x37922, x37923;
  wire x37924, x37925, x37926, x37927, x37928, x37929, x37930, x37931;
  wire x37932, x37933, x37934, x37935, x37936, x37937, x37938, x37939;
  wire x37940, x37941, x37942, x37943, x37944, x37945, x37946, x37947;
  wire x37948, x37949, x37950, x37951, x37952, x37953, x37954, x37955;
  wire x37956, x37957, x37958, x37959, x37960, x37961, x37962, x37963;
  wire x37964, x37965, x37966, x37967, x37968, x37969, x37970, x37971;
  wire x37972, x37973, x37974, x37975, x37976, x37977, x37978, x37979;
  wire x37980, x37981, x37982, x37983, x37984, x37985, x37986, x37987;
  wire x37988, x37989, x37990, x37991, x37992, x37993, x37994, x37995;
  wire x37996, x37997, x37998, x37999, x38000, x38001, x38002, x38003;
  wire x38004, x38005, x38006, x38007, x38008, x38009, x38010, x38011;
  wire x38012, x38013, x38014, x38015, x38016, x38017, x38018, x38019;
  wire x38020, x38021, x38022, x38023, x38024, x38025, x38026, x38027;
  wire x38028, x38029, x38030, x38031, x38032, x38033, x38034, x38035;
  wire x38036, x38037, x38038, x38039, x38040, x38041, x38042, x38043;
  wire x38044, x38045, x38046, x38047, x38048, x38049, x38050, x38051;
  wire x38052, x38053, x38054, x38055, x38056, x38057, x38058, x38059;
  wire x38060, x38061, x38062, x38063, x38064, x38065, x38066, x38067;
  wire x38068, x38069, x38070, x38071, x38072, x38073, x38074, x38075;
  wire x38076, x38077, x38078, x38079, x38080, x38081, x38082, x38083;
  wire x38084, x38085, x38086, x38087, x38088, x38089, x38090, x38091;
  wire x38092, x38093, x38094, x38095, x38096, x38097, x38098, x38099;
  wire x38100, x38101, x38102, x38103, x38104, x38105, x38106, x38107;
  wire x38108, x38109, x38110, x38111, x38112, x38113, x38114, x38115;
  wire x38116, x38117, x38118, x38119, x38120, x38121, x38122, x38123;
  wire x38124, x38125, x38126, x38127, x38128, x38129, x38130, x38131;
  wire x38132, x38133, x38134, x38135, x38136, x38137, x38138, x38139;
  wire x38140, x38141, x38142, x38143, x38144, x38145, x38146, x38147;
  wire x38148, x38149, x38150, x38151, x38152, x38153, x38154, x38155;
  wire x38156, x38157, x38158, x38159, x38160, x38161, x38162, x38163;
  wire x38164, x38165, x38166, x38167, x38168, x38169, x38170, x38171;
  wire x38172, x38173, x38174, x38175, x38176, x38177, x38178, x38179;
  wire x38180, x38181, x38182, x38183, x38184, x38185, x38186, x38187;
  wire x38188, x38189, x38190, x38191, x38192, x38193, x38194, x38195;
  wire x38196, x38197, x38198, x38199, x38200, x38201, x38202, x38203;
  wire x38204, x38205, x38206, x38207, x38208, x38209, x38210, x38211;
  wire x38212, x38213, x38214, x38215, x38216, x38217, x38218, x38219;
  wire x38220, x38221, x38222, x38223, x38224, x38225, x38226, x38227;
  wire x38228, x38229, x38230, x38231, x38232, x38233, x38234, x38235;
  wire x38236, x38237, x38238, x38239, x38240, x38241, x38242, x38243;
  wire x38244, x38245, x38246, x38247, x38248, x38249, x38250, x38251;
  wire x38252, x38253, x38254, x38255, x38256, x38257, x38258, x38259;
  wire x38260, x38261, x38262, x38263, x38264, x38265, x38266, x38267;
  wire x38268, x38269, x38270, x38271, x38272, x38273, x38274, x38275;
  wire x38276, x38277, x38278, x38279, x38280, x38281, x38282, x38283;
  wire x38284, x38285, x38286, x38287, x38288, x38289, x38290, x38291;
  wire x38292, x38293, x38294, x38295, x38296, x38297, x38298, x38299;
  wire x38300, x38301, x38302, x38303, x38304, x38305, x38306, x38307;
  wire x38308, x38309, x38310, x38311, x38312, x38313, x38314, x38315;
  wire x38316, x38317, x38318, x38319, x38320, x38321, x38322, x38323;
  wire x38324, x38325, x38326, x38327, x38328, x38329, x38330, x38331;
  wire x38332, x38333, x38334, x38335, x38336, x38337, x38338, x38339;
  wire x38340, x38341, x38342, x38343, x38344, x38345, x38346, x38347;
  wire x38348, x38349, x38350, x38351, x38352, x38353, x38354, x38355;
  wire x38356, x38357, x38358, x38359, x38360, x38361, x38362, x38363;
  wire x38364, x38365, x38366, x38367, x38368, x38369, x38370, x38371;
  wire x38372, x38373, x38374, x38375, x38376, x38377, x38378, x38379;
  wire x38380, x38381, x38382, x38383, x38384, x38385, x38386, x38387;
  wire x38388, x38389, x38390, x38391, x38392, x38393, x38394, x38395;
  wire x38396, x38397, x38398, x38399, x38400, x38401, x38402, x38403;
  wire x38404, x38405, x38406, x38407, x38408, x38409, x38410, x38411;
  wire x38412, x38413, x38414, x38415, x38416, x38417, x38418, x38419;
  wire x38420, x38421, x38422, x38423, x38424, x38425, x38426, x38427;
  wire x38428, x38429, x38430, x38431, x38432, x38433, x38434, x38435;
  wire x38436, x38437, x38438, x38439, x38440, x38441, x38442, x38443;
  wire x38444, x38445, x38446, x38447, x38448, x38449, x38450, x38451;
  wire x38452, x38453, x38454, x38455, x38456, x38457, x38458, x38459;
  wire x38460, x38461, x38462, x38463, x38464, x38465, x38466, x38467;
  wire x38468, x38469, x38470, x38471, x38472, x38473, x38474, x38475;
  wire x38476, x38477, x38478, x38479, x38480, x38481, x38482, x38483;
  wire x38484, x38485, x38486, x38487, x38488, x38489, x38490, x38491;
  wire x38492, x38493, x38494, x38495, x38496, x38497, x38498, x38499;
  wire x38500, x38501, x38502, x38503, x38504, x38505, x38506, x38507;
  wire x38508, x38509, x38510, x38511, x38512, x38513, x38514, x38515;
  wire x38516, x38517, x38518, x38519, x38520, x38521, x38522, x38523;
  wire x38524, x38525, x38526, x38527, x38528, x38529, x38530, x38531;
  wire x38532, x38533, x38534, x38535, x38536, x38537, x38538, x38539;
  wire x38540, x38541, x38542, x38543, x38544, x38545, x38546, x38547;
  wire x38548, x38549, x38550, x38551, x38552, x38553, x38554, x38555;
  wire x38556, x38557, x38558, x38559, x38560, x38561, x38562, x38563;
  wire x38564, x38565, x38566, x38567, x38568, x38569, x38570, x38571;
  wire x38572, x38573, x38574, x38575, x38576, x38577, x38578, x38579;
  wire x38580, x38581, x38582, x38583, x38584, x38585, x38586, x38587;
  wire x38588, x38589, x38590, x38591, x38592, x38593, x38594, x38595;
  wire x38596, x38597, x38598, x38599, x38600, x38601, x38602, x38603;
  wire x38604, x38605, x38606, x38607, x38608, x38609, x38610, x38611;
  wire x38612, x38613, x38614, x38615, x38616, x38617, x38618, x38619;
  wire x38620, x38621, x38622, x38623, x38624, x38625, x38626, x38627;
  wire x38628, x38629, x38630, x38631, x38632, x38633, x38634, x38635;
  wire x38636, x38637, x38638, x38639, x38640, x38641, x38642, x38643;
  wire x38644, x38645, x38646, x38647, x38648, x38649, x38650, x38651;
  wire x38652, x38653, x38654, x38655, x38656, x38657, x38658, x38659;
  wire x38660, x38661, x38662, x38663, x38664, x38665, x38666, x38667;
  wire x38668, x38669, x38670, x38671, x38672, x38673, x38674, x38675;
  wire x38676, x38677, x38678, x38679, x38680, x38681, x38682, x38683;
  wire x38684, x38685, x38686, x38687, x38688, x38689, x38690, x38691;
  wire x38692, x38693, x38694, x38695, x38696, x38697, x38698, x38699;
  wire x38700, x38701, x38702, x38703, x38704, x38705, x38706, x38707;
  wire x38708, x38709, x38710, x38711, x38712, x38713, x38714, x38715;
  wire x38716, x38717, x38718, x38719, x38720, x38721, x38723, x38724;
  wire x38725, x38727, x38728, x38729, x38731, x38732, x38733, x38735;
  wire x38736, x38737, x38739, x38740, x38741, x38743, x38744, x38745;
  wire x38747, x38748, x38749, x38751, x38752, x38753, x38755, x38756;
  wire x38757, x38759, x38760, x38761, x38763, x38764, x38765, x38767;
  wire x38768, x38769, x38771, x38772, x38773, x38775, x38776, x38777;
  wire x38779, x38780, x38781, x38783, x38784, x38785, x38787, x38788;
  wire x38789, x38791, x38792, x38793, x38795, x38796, x38797, x38799;
  wire x38800, x38801, x38803, x38804, x38805, x38807, x38808, x38809;
  wire x38811, x38812, x38813, x38815, x38816, x38817, x38819, x38820;
  wire x38821, x38823, x38824, x38825, x38827, x38828, x38829, x38831;
  wire x38832, x38833, x38835, x38836, x38837, x38839, x38840, x38841;
  wire x38843, x38844, x38845, x38847, x38848, x38849, x38850, x38851;
  wire x38852, x38853, x38854, x38855, x38856, x38857, x38858, x38859;
  wire x38860, x38861, x38862, x38863, x38864, x38865, x38866, x38867;
  wire x38868, x38869, x38870, x38871, x38872, x38873, x38874, x38875;
  wire x38876, x38877, x38878, x38879, x38880, x38881, x38882, x38883;
  wire x38884, x38885, x38886, x38887, x38888, x38889, x38890, x38891;
  wire x38892, x38893, x38894, x38895, x38896, x38897, x38898, x38899;
  wire x38900, x38901, x38902, x38903, x38904, x38905, x38906, x38907;
  wire x38908, x38909, x38910, x38943, x38944, x38945, x38946, x38947;
  wire x38948, x38949, x38950, x38951, x38952, x38953, x38954, x38955;
  wire x38956, x38957, x38958, x38959, x38960, x38961, x38962, x38963;
  wire x38964, x38965, x38966, x38967, x38968, x38969, x38970, x38971;
  wire x38972, x38973, x38974, x38975, x38976, x38977, x38978, x38979;
  wire x38980, x38981, x38982, x38983, x38984, x38985, x38986, x38987;
  wire x38988, x38989, x38990, x38991, x38992, x38993, x38994, x38995;
  wire x38996, x38997, x38998, x38999, x39000, x39001, x39002, x39003;
  wire x39004, x39005, x39006, x39007, x39008, x39009, x39010, x39011;
  wire x39012, x39013, x39014, x39015, x39016, x39017, x39018, x39019;
  wire x39020, x39021, x39022, x39023, x39024, x39025, x39026, x39027;
  wire x39028, x39029, x39030, x39031, x39032, x39033, x39034, x39035;
  wire x39036, x39037, x39038, x39039, x39042, x39043, x39045, x39048;
  wire x39049, x39051, x39054, x39055, x39057, x39060, x39061, x39063;
  wire x39066, x39067, x39069, x39072, x39073, x39075, x39078, x39079;
  wire x39081, x39084, x39085, x39087, x39090, x39091, x39093, x39096;
  wire x39097, x39099, x39102, x39103, x39105, x39108, x39109, x39111;
  wire x39114, x39115, x39117, x39120, x39121, x39123, x39126, x39127;
  wire x39129, x39132, x39133, x39135, x39138, x39139, x39141, x39144;
  wire x39145, x39147, x39150, x39151, x39153, x39156, x39157, x39159;
  wire x39162, x39163, x39165, x39168, x39169, x39171, x39174, x39175;
  wire x39177, x39180, x39181, x39183, x39186, x39187, x39189, x39192;
  wire x39193, x39195, x39198, x39199, x39201, x39204, x39205, x39207;
  wire x39210, x39211, x39213, x39216, x39217, x39219, x39222, x39223;
  wire x39225, x39228, x39229, x39261, x39262, x39263, x39264, x39265;
  wire x39267, x39268, x39269, x39271, x39272, x39273, x39275, x39276;
  wire x39277, x39279, x39280, x39281, x39283, x39284, x39285, x39287;
  wire x39288, x39289, x39291, x39292, x39293, x39295, x39296, x39297;
  wire x39299, x39300, x39301, x39303, x39304, x39305, x39307, x39308;
  wire x39309, x39311, x39312, x39313, x39315, x39316, x39317, x39319;
  wire x39320, x39321, x39323, x39324, x39325, x39327, x39328, x39329;
  wire x39331, x39332, x39333, x39335, x39336, x39337, x39339, x39340;
  wire x39341, x39343, x39344, x39345, x39347, x39348, x39349, x39351;
  wire x39352, x39353, x39355, x39356, x39357, x39359, x39360, x39361;
  wire x39363, x39364, x39365, x39367, x39368, x39369, x39371, x39372;
  wire x39373, x39375, x39376, x39377, x39379, x39380, x39381, x39383;
  wire x39385, x39386, x39388, x39389, x39391, x39392, x39394, x39396;
  wire x39397, x39399, x39401, x39402, x39404, x39406, x39407, x39409;
  wire x39411, x39412, x39414, x39416, x39417, x39419, x39421, x39422;
  wire x39424, x39426, x39427, x39429, x39431, x39432, x39434, x39436;
  wire x39437, x39439, x39441, x39442, x39444, x39446, x39447, x39449;
  wire x39451, x39452, x39454, x39456, x39457, x39459, x39461, x39462;
  wire x39464, x39466, x39467, x39469, x39471, x39472, x39474, x39476;
  wire x39477, x39479, x39481, x39482, x39484, x39486, x39487, x39489;
  wire x39491, x39492, x39494, x39496, x39497, x39499, x39501, x39502;
  wire x39504, x39506, x39507, x39509, x39511, x39512, x39514, x39516;
  wire x39517, x39519, x39521, x39522, x39524, x39526, x39527, x39529;
  wire x39531, x39532, x39534, x39535, x39537, x39538, x39540, x39541;
  wire x39543, x39544, x39546, x39548, x39549, x39551, x39553, x39554;
  wire x39556, x39558, x39559, x39561, x39563, x39564, x39566, x39568;
  wire x39569, x39571, x39573, x39574, x39576, x39578, x39579, x39581;
  wire x39583, x39584, x39586, x39588, x39589, x39591, x39593, x39594;
  wire x39596, x39598, x39599, x39601, x39603, x39604, x39606, x39608;
  wire x39609, x39611, x39613, x39614, x39616, x39618, x39619, x39621;
  wire x39623, x39624, x39626, x39628, x39629, x39631, x39633, x39634;
  wire x39636, x39638, x39639, x39641, x39643, x39644, x39646, x39648;
  wire x39649, x39651, x39653, x39654, x39656, x39658, x39659, x39661;
  wire x39663, x39664, x39666, x39667, x39669, x39670, x39672, x39673;
  wire x39675, x39676, x39678, x39679, x39681, x39682, x39684, x39685;
  wire x39687, x39688, x39690, x39692, x39693, x39695, x39697, x39698;
  wire x39700, x39702, x39703, x39705, x39707, x39708, x39710, x39712;
  wire x39713, x39715, x39717, x39718, x39720, x39722, x39723, x39725;
  wire x39727, x39728, x39730, x39732, x39733, x39735, x39737, x39738;
  wire x39740, x39742, x39743, x39745, x39747, x39748, x39750, x39752;
  wire x39753, x39755, x39757, x39758, x39760, x39762, x39763, x39765;
  wire x39767, x39768, x39770, x39771, x39773, x39774, x39776, x39777;
  wire x39779, x39780, x39782, x39783, x39785, x39786, x39788, x39789;
  wire x39791, x39792, x39794, x39795, x39797, x39798, x39800, x39801;
  wire x39803, x39804, x39806, x39807, x39809, x39810, x39812, x39813;
  wire x39814, x39816, x39818, x39819, x39821, x39823, x39824, x39826;
  wire x39828, x39829, x39831, x39833, x39834, x39836, x39838, x39839;
  wire x39841, x39843, x39844, x39846, x39848, x39849, x39851, x39853;
  wire x39854, x39856, x39858, x39859, x39861, x39863, x39864, x39866;
  wire x39868, x39869, x39871, x39873, x39874, x39876, x39878, x39879;
  wire x39881, x39883, x39884, x39886, x39888, x39889, x39891, x39893;
  wire x39894, x39896, x39898, x39899, x39901, x39903, x39904, x39906;
  wire x39908, x39909, x39911, x39913, x39914, x39916, x39918, x39919;
  wire x39921, x39923, x39924, x39926, x39928, x39929, x39931, x39933;
  wire x39934, x39936, x39938, x39939, x39941, x39943, x39944, x39946;
  wire x39948, x39949, x39951, x39953, x39954, x39956, x39958, x39959;
  wire x39961, x39963, x39964, x39966, x39968, x39969, x39971, x39972;
  wire x39974, x39976, x39978, x39980, x39982, x39984, x39986, x39988;
  wire x39989, x39991, x39993, x39995, x39997, x39999, x40001, x40003;
  wire x40005, x40007, x40009, x40011, x40013, x40015, x40017, x40019;
  wire x40021, x40023, x40024, x40026, x40028, x40030, x40032, x40034;
  wire x40036, x40038, x40040, x40042, x40044, x40046, x40048, x40050;
  wire x40052, x40054, x40056, x40058, x40060, x40062, x40064, x40066;
  wire x40068, x40070, x40072, x40074, x40076, x40077, x40079, x40081;
  wire x40083, x40085, x40087, x40089, x40091, x40093, x40095, x40097;
  wire x40099, x40101, x40103, x40105, x40107, x40109, x40111, x40113;
  wire x40115, x40117, x40119, x40121, x40123, x40125, x40127, x40129;
  wire x40131, x40133, x40135, x40137, x40139, x40141, x40143, x40145;
  wire x40147, x40148, x40150, x40152, x40154, x40156, x40158, x40160;
  wire x40162, x40164, x40166, x40168, x40170, x40172, x40174, x40176;
  wire x40178, x40180, x40182, x40184, x40186, x40188, x40190, x40192;
  wire x40194, x40196, x40198, x40200, x40202, x40204, x40206, x40208;
  wire x40210, x40212, x40214, x40216, x40218, x40220, x40222, x40224;
  wire x40226, x40228, x40230, x40232, x40234, x40236, x40237, x40239;
  wire x40241, x40243, x40245, x40247, x40249, x40251, x40253, x40255;
  wire x40257, x40259, x40261, x40263, x40265, x40267, x40269, x40271;
  wire x40273, x40275, x40277, x40279, x40281, x40283, x40285, x40287;
  wire x40289, x40291, x40293, x40295, x40297, x40299, x40301, x40303;
  wire x40305, x40307, x40309, x40311, x40313, x40315, x40317, x40319;
  wire x40321, x40323, x40325, x40327, x40329, x40331, x40333, x40335;
  wire x40337, x40339, x40341, x40343, x40344, x40346, x40348, x40350;
  wire x40352, x40354, x40356, x40358, x40360, x40362, x40364, x40366;
  wire x40368, x40370, x40372, x40374, x40376, x40378, x40380, x40382;
  wire x40384, x40386, x40388, x40390, x40392, x40394, x40396, x40398;
  wire x40400, x40402, x40404, x40406, x40408, x40410, x40412, x40414;
  wire x40416, x40418, x40420, x40422, x40424, x40426, x40428, x40430;
  wire x40432, x40434, x40436, x40438, x40440, x40442, x40444, x40446;
  wire x40448, x40450, x40452, x40454, x40456, x40458, x40460, x40462;
  wire x40464, x40466, x40468, x40469, x40471, x40473, x40475, x40477;
  wire x40479, x40481, x40483, x40485, x40487, x40489, x40491, x40493;
  wire x40495, x40497, x40499, x40501, x40503, x40505, x40507, x40509;
  wire x40511, x40513, x40515, x40517, x40519, x40521, x40523, x40525;
  wire x40527, x40529, x40531, x40533, x40535, x40537, x40539, x40541;
  wire x40543, x40545, x40547, x40549, x40551, x40553, x40555, x40557;
  wire x40559, x40561, x40563, x40565, x40567, x40569, x40571, x40573;
  wire x40575, x40577, x40579, x40581, x40583, x40585, x40587, x40589;
  wire x40591, x40593, x40595, x40597, x40599, x40601, x40603, x40605;
  wire x40607, x40609, x40611, x40612, x40614, x40616, x40618, x40620;
  wire x40622, x40624, x40626, x40628, x40630, x40632, x40634, x40636;
  wire x40638, x40640, x40642, x40644, x40646, x40648, x40650, x40652;
  wire x40654, x40656, x40658, x40660, x40662, x40664, x40666, x40668;
  wire x40670, x40672, x40674, x40676, x40678, x40680, x40682, x40684;
  wire x40686, x40688, x40690, x40692, x40694, x40696, x40698, x40700;
  wire x40702, x40704, x40706, x40708, x40710, x40712, x40714, x40716;
  wire x40718, x40720, x40722, x40724, x40726, x40728, x40730, x40732;
  wire x40734, x40736, x40738, x40740, x40742, x40744, x40746, x40748;
  wire x40750, x40752, x40754, x40756, x40758, x40760, x40762, x40764;
  wire x40766, x40768, x40770, x40772, x40773, x40775, x40777, x40779;
  wire x40781, x40783, x40785, x40787, x40789, x40791, x40793, x40795;
  wire x40797, x40799, x40801, x40803, x40805, x40807, x40809, x40811;
  wire x40813, x40815, x40817, x40819, x40821, x40823, x40825, x40827;
  wire x40829, x40831, x40833, x40835, x40837, x40839, x40841, x40843;
  wire x40845, x40847, x40849, x40851, x40853, x40855, x40857, x40859;
  wire x40861, x40863, x40865, x40867, x40869, x40871, x40873, x40875;
  wire x40877, x40879, x40881, x40883, x40885, x40887, x40889, x40891;
  wire x40893, x40895, x40897, x40899, x40901, x40903, x40905, x40907;
  wire x40909, x40911, x40913, x40915, x40917, x40919, x40921, x40923;
  wire x40925, x40927, x40929, x40931, x40933, x40935, x40937, x40939;
  wire x40941, x40943, x40945, x40947, x40949, x40951, x40952, x40954;
  wire x40956, x40958, x40960, x40962, x40964, x40966, x40968, x40970;
  wire x40972, x40974, x40976, x40978, x40980, x40982, x40984, x40986;
  wire x40988, x40990, x40992, x40994, x40996, x40998, x41000, x41002;
  wire x41004, x41006, x41008, x41010, x41012, x41014, x41016, x41017;
  wire x41018, x41019, x41020, x41021, x41023, x41024, x41025, x41026;
  wire x41027, x41028, x41029, x41031, x41032, x41033, x41034, x41035;
  wire x41036, x41037, x41039, x41040, x41041, x41042, x41043, x41044;
  wire x41045, x41046, x41047, x41048, x41050, x41051, x41052, x41053;
  wire x41054, x41055, x41056, x41058, x41059, x41060, x41061, x41062;
  wire x41063, x41064, x41066, x41067, x41068, x41069, x41070, x41071;
  wire x41072, x41074, x41075, x41076, x41078, x41079, x41080, x41081;
  wire x41083, x41084, x41085, x41086, x41087, x41088, x41089, x41091;
  wire x41092, x41093, x41095, x41096, x41097, x41098, x41099, x41100;
  wire x41101, x41103, x41104, x41105, x41106, x41107, x41108, x41109;
  wire x41111, x41112, x41113, x41115, x41116, x41117, x41118, x41120;
  wire x41121, x41122, x41124, x41125, x41126, x41127, x41129, x41130;
  wire x41131, x41132, x41133, x41134, x41135, x41137, x41138, x41139;
  wire x41141, x41142, x41143, x41144, x41146, x41147, x41148, x41150;
  wire x41151, x41152, x41153, x41155, x41156, x41157, x41158, x41159;
  wire x41160, x41161, x41163, x41164, x41165, x41167, x41168, x41169;
  wire x41170, x41172, x41173, x41174, x41176, x41177, x41178, x41179;
  wire x41180, x41181, x41182, x41184, x41185, x41186, x41187, x41188;
  wire x41189, x41190, x41192, x41193, x41194, x41196, x41197, x41198;
  wire x41199, x41201, x41202, x41203, x41205, x41206, x41207, x41208;
  wire x41210, x41211, x41212, x41214, x41215, x41216, x41217, x41219;
  wire x41220, x41221, x41222, x41223, x41224, x41225, x41227, x41228;
  wire x41229, x41231, x41232, x41233, x41234, x41236, x41237, x41238;
  wire x41240, x41241, x41242, x41243, x41245, x41246, x41247, x41249;
  wire x41250, x41251, x41252, x41254, x41255, x41256, x41257, x41258;
  wire x41259, x41260, x41262, x41263, x41264, x41266, x41267, x41268;
  wire x41269, x41271, x41272, x41273, x41275, x41276, x41277, x41278;
  wire x41280, x41281, x41282, x41284, x41285, x41286, x41287, x41288;
  wire x41289, x41290, x41292, x41293, x41294, x41295, x41296, x41297;
  wire x41298, x41300, x41301, x41302, x41304, x41305, x41306, x41307;
  wire x41309, x41310, x41311, x41313, x41314, x41315, x41316, x41318;
  wire x41319, x41320, x41322, x41323, x41324, x41325, x41327, x41328;
  wire x41329, x41330, x41331, x41332, x41333, x41335, x41336, x41337;
  wire x41338, x41339, x41340, x41341, x41343, x41344, x41345, x41347;
  wire x41348, x41349, x41350, x41352, x41353, x41354, x41356, x41357;
  wire x41358, x41359, x41361, x41362, x41363, x41365, x41366, x41367;
  wire x41368, x41370, x41371, x41372, x41374, x41375, x41376, x41377;
  wire x41379, x41380, x41381, x41382, x41383, x41384, x41385, x41387;
  wire x41388, x41389, x41391, x41392, x41393, x41394, x41396, x41397;
  wire x41398, x41400, x41401, x41402, x41403, x41405, x41406, x41407;
  wire x41409, x41410, x41411, x41412, x41414, x41415, x41416, x41418;
  wire x41419, x41420, x41421, x41422, x41423, x41424, x41426, x41427;
  wire x41428, x41429, x41430, x41431, x41432, x41434, x41435, x41436;
  wire x41438, x41439, x41440, x41441, x41443, x41444, x41445, x41447;
  wire x41448, x41449, x41450, x41452, x41453, x41454, x41456, x41457;
  wire x41458, x41459, x41461, x41462, x41463, x41465, x41466, x41467;
  wire x41468, x41470, x41471, x41472, x41474, x41475, x41476, x41477;
  wire x41479, x41480, x41481, x41482, x41483, x41484, x41485, x41487;
  wire x41488, x41489, x41491, x41492, x41493, x41494, x41496, x41497;
  wire x41498, x41500, x41501, x41502, x41503, x41505, x41506, x41507;
  wire x41509, x41510, x41511, x41512, x41514, x41515, x41516, x41518;
  wire x41519, x41520, x41521, x41523, x41524, x41525, x41527, x41528;
  wire x41529, x41530, x41532, x41533, x41534, x41535, x41536, x41537;
  wire x41538, x41540, x41541, x41542, x41544, x41545, x41546, x41547;
  wire x41549, x41550, x41551, x41553, x41554, x41555, x41556, x41558;
  wire x41559, x41560, x41562, x41563, x41564, x41565, x41567, x41568;
  wire x41569, x41571, x41572, x41573, x41574, x41576, x41577, x41578;
  wire x41580, x41581, x41582, x41583, x41584, x41585, x41586, x41588;
  wire x41589, x41590, x41591, x41592, x41593, x41594, x41596, x41597;
  wire x41598, x41600, x41601, x41602, x41603, x41605, x41606, x41607;
  wire x41609, x41610, x41611, x41612, x41614, x41615, x41616, x41618;
  wire x41619, x41620, x41621, x41623, x41624, x41625, x41627, x41628;
  wire x41629, x41630, x41632, x41633, x41634, x41636, x41637, x41638;
  wire x41639, x41641, x41642, x41643, x41645, x41646, x41647, x41648;
  wire x41650, x41651, x41652, x41653, x41654, x41655, x41656, x41658;
  wire x41659, x41660, x41662, x41663, x41664, x41665, x41667, x41668;
  wire x41669, x41671, x41672, x41673, x41674, x41676, x41677, x41678;
  wire x41680, x41681, x41682, x41683, x41685, x41686, x41687, x41689;
  wire x41690, x41691, x41692, x41694, x41695, x41696, x41698, x41699;
  wire x41700, x41701, x41703, x41704, x41705, x41707, x41708, x41709;
  wire x41710, x41712, x41713, x41714, x41715, x41716, x41717, x41718;
  wire x41720, x41721, x41722, x41724, x41725, x41726, x41727, x41729;
  wire x41730, x41731, x41733, x41734, x41735, x41736, x41738, x41739;
  wire x41740, x41742, x41743, x41744, x41745, x41747, x41748, x41749;
  wire x41751, x41752, x41753, x41754, x41756, x41757, x41758, x41760;
  wire x41761, x41762, x41763, x41765, x41766, x41767, x41769, x41770;
  wire x41771, x41772, x41773, x41774, x41775, x41777, x41778, x41779;
  wire x41780, x41781, x41782, x41783, x41785, x41786, x41787, x41789;
  wire x41790, x41791, x41792, x41794, x41795, x41796, x41798, x41799;
  wire x41800, x41801, x41803, x41804, x41805, x41807, x41808, x41809;
  wire x41810, x41812, x41813, x41814, x41816, x41817, x41818, x41819;
  wire x41821, x41822, x41823, x41825, x41826, x41827, x41828, x41830;
  wire x41831, x41832, x41834, x41835, x41836, x41837, x41839, x41840;
  wire x41841, x41842, x41843, x41844, x41845, x41847, x41848, x41849;
  wire x41850, x41851, x41852, x41853, x41855, x41856, x41857, x41859;
  wire x41860, x41861, x41862, x41864, x41865, x41866, x41868, x41869;
  wire x41870, x41871, x41873, x41874, x41875, x41877, x41878, x41879;
  wire x41880, x41882, x41883, x41884, x41886, x41887, x41888, x41889;
  wire x41891, x41892, x41893, x41895, x41896, x41897, x41898, x41900;
  wire x41901, x41902, x41904, x41905, x41906, x41907, x41909, x41910;
  wire x41911, x41913, x41914, x41915, x41916, x41918, x41919, x41920;
  wire x41921, x41922, x41923, x41924, x41926, x41927, x41928, x41930;
  wire x41931, x41932, x41933, x41935, x41936, x41937, x41939, x41940;
  wire x41941, x41942, x41944, x41945, x41946, x41948, x41949, x41950;
  wire x41951, x41953, x41954, x41955, x41957, x41958, x41959, x41960;
  wire x41962, x41963, x41964, x41966, x41967, x41968, x41969, x41971;
  wire x41972, x41973, x41975, x41976, x41977, x41978, x41980, x41981;
  wire x41982, x41984, x41985, x41986, x41987, x41988, x41989, x41990;
  wire x41992, x41993, x41994, x41995, x41996, x41997, x41998, x42000;
  wire x42001, x42002, x42004, x42005, x42006, x42007, x42009, x42010;
  wire x42011, x42013, x42014, x42015, x42016, x42018, x42019, x42020;
  wire x42022, x42023, x42024, x42025, x42027, x42028, x42029, x42031;
  wire x42032, x42033, x42034, x42036, x42037, x42038, x42040, x42041;
  wire x42042, x42043, x42045, x42046, x42047, x42049, x42050, x42051;
  wire x42052, x42054, x42055, x42056, x42058, x42059, x42060, x42061;
  wire x42063, x42064, x42065, x42067, x42068, x42069, x42070, x42072;
  wire x42073, x42074, x42075, x42076, x42077, x42078, x42080, x42081;
  wire x42082, x42084, x42085, x42086, x42087, x42089, x42090, x42091;
  wire x42093, x42094, x42095, x42096, x42098, x42099, x42100, x42102;
  wire x42103, x42104, x42105, x42107, x42108, x42109, x42111, x42112;
  wire x42113, x42114, x42116, x42117, x42118, x42120, x42121, x42122;
  wire x42123, x42125, x42126, x42127, x42129, x42130, x42131, x42132;
  wire x42134, x42135, x42136, x42138, x42139, x42140, x42141, x42143;
  wire x42144, x42145, x42147, x42148, x42149, x42150, x42152, x42153;
  wire x42154, x42155, x42156, x42157, x42158, x42160, x42161, x42162;
  wire x42164, x42165, x42166, x42167, x42169, x42170, x42171, x42173;
  wire x42174, x42175, x42176, x42178, x42179, x42180, x42182, x42183;
  wire x42184, x42185, x42187, x42188, x42189, x42191, x42192, x42193;
  wire x42194, x42196, x42197, x42198, x42200, x42201, x42202, x42203;
  wire x42205, x42206, x42207, x42209, x42210, x42211, x42212, x42214;
  wire x42215, x42216, x42218, x42219, x42220, x42221, x42223, x42224;
  wire x42225, x42227, x42228, x42229, x42230, x42231, x42232, x42233;
  wire x42235, x42236, x42237, x42239, x42240, x42241, x42242, x42244;
  wire x42245, x42246, x42248, x42249, x42250, x42251, x42253, x42254;
  wire x42255, x42257, x42258, x42259, x42260, x42262, x42263, x42264;
  wire x42266, x42267, x42268, x42269, x42271, x42272, x42273, x42275;
  wire x42276, x42277, x42278, x42280, x42281, x42282, x42284, x42285;
  wire x42286, x42287, x42289, x42290, x42291, x42293, x42294, x42295;
  wire x42296, x42298, x42299, x42300, x42302, x42303, x42304, x42305;
  wire x42307, x42308, x42309, x42311, x42312, x42313, x42314, x42316;
  wire x42317, x42318, x42320, x42321, x42322, x42323, x42325, x42326;
  wire x42327, x42329, x42330, x42331, x42332, x42334, x42335, x42336;
  wire x42338, x42339, x42340, x42341, x42343, x42344, x42345, x42347;
  wire x42348, x42349, x42350, x42352, x42353, x42354, x42356, x42357;
  wire x42358, x42359, x42361, x42362, x42363, x42365, x42366, x42367;
  wire x42368, x42370, x42371, x42372, x42374, x42375, x42376, x42377;
  wire x42379, x42380, x42381, x42383, x42384, x42385, x42386, x42388;
  wire x42389, x42390, x42392, x42393, x42394, x42395, x42397, x42398;
  wire x42399, x42401, x42402, x42403, x42404, x42406, x42407, x42408;
  wire x42410, x42411, x42412, x42413, x42415, x42416, x42417, x42419;
  wire x42420, x42421, x42423, x42424, x42425, x42427, x42428, x42429;
  wire x42431, x42432, x42433, x42435, x42436, x42437, x42439, x42440;
  wire x42441, x42443, x42444, x42445, x42447, x42448, x42449, x42451;
  wire x42452, x42453, x42455, x42456, x42457, x42459, x42460, x42461;
  wire x42463, x42464, x42465, x42467, x42468, x42469, x42471, x42472;
  wire x42473, x42475, x42476, x42477, x42479, x42480, x42481, x42483;
  wire x42484, x42485, x42487, x42488, x42489, x42491, x42492, x42493;
  wire x42497, x42499, x42500, x42501, x42504, x42505, x42506, x42507;
  wire x42508, x42509, x42512, x42513, x42514, x42515, x42516, x42517;
  wire x42520, x42521, x42523, x42524, x42525, x42526, x42527, x42528;
  wire x42529, x42530, x42533, x42534, x42536, x42538, x42539, x42540;
  wire x42541, x42542, x42543, x42545, x42546, x42547, x42549, x42550;
  wire x42553, x42554, x42556, x42558, x42559, x42560, x42561, x42562;
  wire x42563, x42565, x42566, x42567, x42569, x42570, x42573, x42574;
  wire x42576, x42578, x42579, x42580, x42581, x42582, x42583, x42585;
  wire x42586, x42587, x42589, x42590, x42593, x42594, x42596, x42598;
  wire x42599, x42600, x42602, x42603, x42604, x42606, x42607, x42608;
  wire x42610, x42611, x42614, x42615, x42617, x42619, x42620, x42621;
  wire x42623, x42624, x42625, x42627, x42628, x42629, x42631, x42632;
  wire x42635, x42636, x42638, x42640, x42641, x42642, x42643, x42645;
  wire x42646, x42647, x42648, x42649, x42651, x42652, x42653, x42655;
  wire x42656, x42659, x42660, x42662, x42664, x42665, x42666, x42667;
  wire x42670, x42671, x42672, x42673, x42674, x42676, x42677, x42678;
  wire x42680, x42681, x42682, x42683, x42684, x42687, x42688, x42690;
  wire x42692, x42693, x42694, x42695, x42698, x42699, x42700, x42701;
  wire x42702, x42704, x42705, x42706, x42708, x42709, x42710, x42711;
  wire x42712, x42715, x42716, x42718, x42720, x42721, x42722, x42723;
  wire x42726, x42727, x42729, x42730, x42731, x42733, x42734, x42735;
  wire x42736, x42738, x42739, x42740, x42742, x42743, x42744, x42745;
  wire x42746, x42749, x42750, x42752, x42754, x42755, x42756, x42757;
  wire x42760, x42761, x42763, x42765, x42766, x42768, x42769, x42770;
  wire x42771, x42773, x42774, x42775, x42777, x42778, x42779, x42780;
  wire x42782, x42783, x42784, x42785, x42786, x42789, x42790, x42792;
  wire x42794, x42795, x42796, x42797, x42800, x42801, x42803, x42805;
  wire x42806, x42808, x42809, x42810, x42811, x42813, x42814, x42815;
  wire x42817, x42818, x42819, x42820, x42822, x42823, x42824, x42825;
  wire x42826, x42829, x42830, x42832, x42834, x42835, x42836, x42837;
  wire x42840, x42841, x42843, x42845, x42846, x42848, x42849, x42850;
  wire x42851, x42853, x42854, x42855, x42857, x42858, x42859, x42860;
  wire x42862, x42863, x42864, x42865, x42866, x42869, x42870, x42872;
  wire x42874, x42875, x42876, x42877, x42880, x42881, x42883, x42885;
  wire x42886, x42888, x42890, x42891, x42892, x42894, x42895, x42896;
  wire x42898, x42899, x42900, x42901, x42903, x42904, x42905, x42907;
  wire x42908, x42911, x42912, x42914, x42916, x42917, x42918, x42919;
  wire x42922, x42923, x42925, x42927, x42928, x42930, x42932, x42933;
  wire x42934, x42936, x42937, x42938, x42940, x42941, x42942, x42943;
  wire x42945, x42946, x42947, x42949, x42950, x42953, x42954, x42956;
  wire x42958, x42959, x42960, x42961, x42964, x42965, x42967, x42969;
  wire x42970, x42972, x42973, x42975, x42976, x42977, x42978, x42979;
  wire x42981, x42982, x42983, x42985, x42986, x42987, x42988, x42990;
  wire x42991, x42992, x42994, x42995, x42998, x42999, x43001, x43003;
  wire x43004, x43005, x43006, x43009, x43010, x43012, x43014, x43015;
  wire x43017, x43018, x43021, x43022, x43023, x43024, x43025, x43027;
  wire x43028, x43029, x43031, x43032, x43033, x43034, x43036, x43037;
  wire x43038, x43040, x43041, x43042, x43043, x43044, x43047, x43048;
  wire x43050, x43052, x43053, x43055, x43056, x43059, x43060, x43062;
  wire x43064, x43065, x43067, x43068, x43071, x43072, x43073, x43074;
  wire x43075, x43077, x43078, x43079, x43081, x43082, x43083, x43084;
  wire x43086, x43087, x43088, x43090, x43091, x43092, x43093, x43094;
  wire x43097, x43098, x43100, x43102, x43103, x43105, x43106, x43109;
  wire x43110, x43112, x43114, x43115, x43117, x43118, x43121, x43122;
  wire x43124, x43125, x43126, x43128, x43129, x43130, x43131, x43133;
  wire x43134, x43135, x43137, x43138, x43139, x43140, x43142, x43143;
  wire x43144, x43146, x43147, x43148, x43149, x43150, x43153, x43154;
  wire x43156, x43158, x43159, x43161, x43162, x43165, x43166, x43168;
  wire x43170, x43171, x43173, x43174, x43177, x43178, x43180, x43182;
  wire x43183, x43185, x43186, x43187, x43188, x43190, x43191, x43192;
  wire x43194, x43195, x43196, x43197, x43199, x43200, x43201, x43203;
  wire x43204, x43205, x43206, x43208, x43209, x43210, x43212, x43213;
  wire x43216, x43217, x43219, x43221, x43222, x43224, x43225, x43228;
  wire x43229, x43231, x43233, x43234, x43236, x43237, x43240, x43241;
  wire x43243, x43245, x43246, x43248, x43249, x43250, x43251, x43253;
  wire x43254, x43255, x43257, x43258, x43259, x43260, x43262, x43263;
  wire x43264, x43266, x43267, x43268, x43269, x43271, x43272, x43273;
  wire x43275, x43276, x43279, x43280, x43282, x43284, x43285, x43287;
  wire x43288, x43291, x43292, x43294, x43296, x43297, x43299, x43300;
  wire x43303, x43304, x43306, x43308, x43309, x43311, x43312, x43313;
  wire x43314, x43316, x43317, x43318, x43320, x43321, x43322, x43324;
  wire x43325, x43326, x43327, x43329, x43330, x43331, x43333, x43334;
  wire x43335, x43336, x43338, x43339, x43340, x43342, x43343, x43346;
  wire x43347, x43349, x43351, x43352, x43354, x43355, x43358, x43359;
  wire x43361, x43363, x43364, x43366, x43367, x43370, x43371, x43373;
  wire x43375, x43376, x43378, x43380, x43381, x43382, x43384, x43385;
  wire x43386, x43388, x43389, x43390, x43392, x43393, x43394, x43395;
  wire x43397, x43398, x43399, x43401, x43402, x43403, x43404, x43406;
  wire x43407, x43408, x43410, x43411, x43414, x43415, x43417, x43419;
  wire x43420, x43422, x43425, x43426, x43428, x43430, x43431, x43433;
  wire x43436, x43437, x43439, x43441, x43442, x43445, x43446, x43447;
  wire x43449, x43450, x43451, x43453, x43454, x43455, x43457, x43458;
  wire x43459, x43461, x43462, x43463, x43465, x43466, x43467, x43469;
  wire x43470, x43471, x43473, x43474, x43475, x43477, x43478, x43479;
  wire x43481, x43482, x43483, x43485, x43486, x43487, x43489, x43490;
  wire x43491, x43493, x43494, x43495, x43498, x43499, x43500, x43504;
  wire x43505, x43506, x43510, x43511, x43512, x43514, x43515, x43516;
  wire x43520, x43521, x43522, x43524, x43525, x43526, x43530, x43531;
  wire x43532, x43534, x43535, x43536, x43540, x43541, x43542, x43544;
  wire x43545, x43546, x43548, x43550, x43551, x43553, x43554, x43555;
  wire x43557, x43558, x43559, x43561, x43563, x43564, x43566, x43567;
  wire x43568, x43570, x43571, x43572, x43574, x43575, x43576, x43578;
  wire x43580, x43581, x43583, x43584, x43585, x43587, x43588, x43589;
  wire x43591, x43592, x43593, x43595, x43598, x43599, x43601, x43602;
  wire x43603, x43605, x43606, x43607, x43609, x43610, x43611, x43613;
  wire x43616, x43617, x43619, x43621, x43622, x43624, x43625, x43626;
  wire x43628, x43629, x43630, x43632, x43635, x43636, x43638, x43640;
  wire x43641, x43643, x43644, x43645, x43647, x43648, x43649, x43651;
  wire x43652, x43653, x43655, x43656, x43659, x43660, x43662, x43664;
  wire x43665, x43667, x43668, x43669, x43671, x43672, x43673, x43675;
  wire x43676, x43677, x43679, x43680, x43681, x43682, x43683, x43686;
  wire x43687, x43689, x43691, x43692, x43694, x43695, x43696, x43698;
  wire x43699, x43700, x43702, x43703, x43704, x43706, x43707, x43708;
  wire x43709, x43710, x43713, x43714, x43716, x43718, x43719, x43721;
  wire x43722, x43723, x43725, x43726, x43727, x43729, x43730, x43731;
  wire x43733, x43734, x43735, x43736, x43737, x43740, x43741, x43743;
  wire x43744, x43745, x43747, x43749, x43751, x43752, x43754, x43755;
  wire x43756, x43758, x43759, x43760, x43762, x43763, x43764, x43766;
  wire x43767, x43768, x43769, x43770, x43773, x43774, x43776, x43777;
  wire x43778, x43780, x43782, x43784, x43785, x43787, x43788, x43789;
  wire x43791, x43792, x43793, x43795, x43796, x43797, x43798, x43800;
  wire x43801, x43802, x43804, x43805, x43806, x43807, x43808, x43811;
  wire x43812, x43814, x43815, x43816, x43818, x43820, x43822, x43823;
  wire x43825, x43826, x43827, x43829, x43830, x43831, x43833, x43834;
  wire x43835, x43836, x43838, x43839, x43840, x43842, x43843, x43844;
  wire x43845, x43846, x43849, x43850, x43852, x43854, x43855, x43857;
  wire x43859, x43861, x43862, x43864, x43865, x43866, x43868, x43869;
  wire x43870, x43872, x43873, x43874, x43875, x43877, x43878, x43879;
  wire x43881, x43882, x43883, x43884, x43885, x43888, x43889, x43891;
  wire x43893, x43894, x43896, x43898, x43900, x43901, x43903, x43905;
  wire x43906, x43908, x43909, x43910, x43912, x43913, x43914, x43915;
  wire x43917, x43918, x43919, x43921, x43922, x43923, x43924, x43925;
  wire x43928, x43929, x43931, x43933, x43934, x43936, x43938, x43940;
  wire x43941, x43943, x43945, x43946, x43948, x43949, x43950, x43952;
  wire x43953, x43954, x43955, x43957, x43958, x43959, x43961, x43962;
  wire x43963, x43964, x43965, x43968, x43969, x43971, x43973, x43974;
  wire x43976, x43977, x43979, x43980, x43982, x43984, x43985, x43987;
  wire x43988, x43990, x43991, x43993, x43994, x43995, x43997, x43998;
  wire x43999, x44000, x44002, x44003, x44004, x44006, x44007, x44008;
  wire x44009, x44011, x44012, x44013, x44015, x44016, x44019, x44020;
  wire x44022, x44024, x44025, x44027, x44029, x44030, x44032, x44034;
  wire x44035, x44037, x44039, x44040, x44042, x44043, x44044, x44046;
  wire x44047, x44048, x44050, x44051, x44052, x44054, x44055, x44056;
  wire x44058, x44059, x44060, x44062, x44063, x44064, x44065, x44066;
  wire x44067, x44068, x44069, x44070, x44072, x44073, x44074, x44076;
  wire x44077, x44078, x44079, x44080, x44081, x44083, x44084, x44085;
  wire x44086, x44087, x44088, x44090, x44091, x44092, x44094, x44095;
  wire x44096, x44097, x44098, x44099, x44100, x44102, x44103, x44104;
  wire x44106, x44107, x44108, x44109, x44110, x44111, x44112, x44114;
  wire x44115, x44116, x44118, x44119, x44120, x44121, x44122, x44123;
  wire x44124, x44126, x44127, x44128, x44130, x44131, x44132, x44133;
  wire x44134, x44135, x44136, x44138, x44139, x44140, x44142, x44143;
  wire x44144, x44145, x44147, x44148, x44149, x44151, x44152, x44153;
  wire x44155, x44156, x44157, x44158, x44160, x44161, x44162, x44164;
  wire x44165, x44166, x44168, x44169, x44170, x44171, x44173, x44174;
  wire x44175, x44177, x44178, x44179, x44181, x44182, x44183, x44184;
  wire x44186, x44187, x44188, x44190, x44191, x44192, x44194, x44195;
  wire x44196, x44197, x44199, x44200, x44201, x44203, x44204, x44205;
  wire x44207, x44208, x44209, x44211, x44212, x44213, x44214, x44216;
  wire x44217, x44218, x44220, x44221, x44222, x44223, x44225, x44226;
  wire x44227, x44229, x44230, x44231, x44233, x44234, x44235, x44236;
  wire x44238, x44239, x44240, x44242, x44243, x44244, x44245, x44247;
  wire x44248, x44249, x44251, x44252, x44253, x44255, x44256, x44257;
  wire x44258, x44260, x44261, x44262, x44264, x44265, x44266, x44267;
  wire x44269, x44270, x44271, x44273, x44274, x44275, x44277, x44278;
  wire x44279, x44280, x44282, x44283, x44284, x44286, x44287, x44288;
  wire x44289, x44291, x44292, x44293, x44295, x44296, x44297, x44299;
  wire x44300, x44301, x44302, x44304, x44305, x44306, x44308, x44310;
  wire x44311, x44312, x44314, x44315, x44316, x44318, x44319, x44320;
  wire x44322, x44323, x44324, x44325, x44327, x44328, x44329, x44331;
  wire x44332, x44334, x44335, x44337, x44338, x44339, x44341, x44342;
  wire x44343, x44344, x44346, x44347, x44348, x44350, x44351, x44352;
  wire x44353, x44355, x44356, x44357, x44359, x44360, x44362, x44363;
  wire x44365, x44366, x44367, x44369, x44370, x44371, x44372, x44374;
  wire x44375, x44376, x44378, x44379, x44380, x44381, x44383, x44384;
  wire x44385, x44387, x44388, x44390, x44391, x44393, x44394, x44395;
  wire x44397, x44398, x44399, x44400, x44402, x44403, x44404, x44406;
  wire x44407, x44409, x44410, x44412, x44413, x44414, x44416, x44417;
  wire x44419, x44420, x44422, x44423, x44424, x44426, x44427, x44428;
  wire x44429, x44431, x44432, x44433, x44435, x44436, x44438, x44439;
  wire x44441, x44443, x44444, x44446, x44447, x44449, x44450, x44452;
  wire x44453, x44454, x44456, x44457, x44458, x44459, x44461, x44462;
  wire x44463, x44465, x44466, x44468, x44469, x44471, x44473, x44474;
  wire x44476, x44477, x44479, x44480, x44482, x44483, x44484, x44486;
  wire x44487, x44488, x44489, x44491, x44492, x44493, x44495, x44496;
  wire x44498, x44499, x44501, x44503, x44504, x44506, x44507, x44509;
  wire x44510, x44512, x44513, x44514, x44516, x44517, x44518, x44519;
  wire x44521, x44522, x44523, x44525, x44526, x44528, x44529, x44531;
  wire x44533, x44534, x44536, x44537, x44539, x44540, x44542, x44543;
  wire x44544, x44546, x44547, x44548, x44549, x44551, x44552, x44553;
  wire x44555, x44556, x44558, x44559, x44561, x44563, x44564, x44566;
  wire x44567, x44569, x44570, x44572, x44573, x44574, x44576, x44577;
  wire x44578, x44579, x44581, x44582, x44583, x44585, x44586, x44589;
  wire x44590, x44592, x44594, x44595, x44597, x44600, x44601, x44603;
  wire x44604, x44605, x44607, x44608, x44609, x44611, x44612, x44613;
  wire x44615, x44616, x44617, x44618, x44619, x44620, x44621, x44622;
  wire x44623, x44624, x44625, x44626, x44628, x44629, x44630, x44631;
  wire x44633, x44634, x44636, x44637, x44638, x44639, x44641, x44642;
  wire x44644, x44645, x44646, x44647, x44649, x44650, x44652, x44653;
  wire x44654, x44655, x44657, x44658, x44660, x44661, x44662, x44663;
  wire x44665, x44666, x44668, x44669, x44670, x44672, x44673, x44674;
  wire x44676, x44677, x44679, x44680, x44682, x44683, x44684, x44686;
  wire x44687, x44688, x44690, x44691, x44693, x44694, x44696, x44697;
  wire x44698, x44700, x44701, x44702, x44704, x44705, x44707, x44708;
  wire x44710, x44711, x44712, x44714, x44715, x44716, x44718, x44719;
  wire x44721, x44722, x44724, x44725, x44726, x44728, x44729, x44730;
  wire x44732, x44733, x44734, x44735, x44737, x44739, x44740, x44742;
  wire x44743, x44744, x44745, x44747, x44748, x44749, x44751, x44752;
  wire x44754, x44755, x44757, x44759, x44760, x44762, x44763, x44764;
  wire x44765, x44767, x44768, x44769, x44771, x44772, x44774, x44775;
  wire x44777, x44779, x44780, x44782, x44783, x44784, x44785, x44787;
  wire x44788, x44789, x44791, x44792, x44794, x44795, x44797, x44799;
  wire x44800, x44802, x44803, x44804, x44805, x44807, x44808, x44809;
  wire x44811, x44812, x44814, x44815, x44817, x44819, x44820, x44822;
  wire x44823, x44824, x44825, x44827, x44828, x44829, x44831, x44832;
  wire x44834, x44835, x44837, x44839, x44840, x44842, x44843, x44844;
  wire x44845, x44847, x44848, x44849, x44851, x44852, x44855, x44856;
  wire x44858, x44860, x44861, x44863, x44864, x44865, x44866, x44868;
  wire x44869, x44870, x44872, x44873, x44876, x44877, x44879, x44881;
  wire x44882, x44884, x44885, x44886, x44887, x44889, x44890, x44891;
  wire x44893, x44894, x44897, x44898, x44900, x44902, x44903, x44905;
  wire x44906, x44907, x44908, x44910, x44911, x44912, x44914, x44915;
  wire x44918, x44919, x44921, x44923, x44924, x44926, x44927, x44928;
  wire x44929, x44931, x44932, x44933, x44935, x44936, x44939, x44940;
  wire x44942, x44944, x44945, x44947, x44948, x44949, x44950, x44952;
  wire x44953, x44954, x44956, x44957, x44960, x44961, x44963, x44965;
  wire x44966, x44968, x44969, x44970, x44971, x44973, x44974, x44975;
  wire x44977, x44978, x44981, x44982, x44984, x44986, x44987, x44989;
  wire x44990, x44991, x44992, x44994, x44995, x44996, x44998, x44999;
  wire x45002, x45003, x45005, x45007, x45008, x45010, x45011, x45012;
  wire x45013, x45015, x45016, x45017, x45019, x45020, x45023, x45024;
  wire x45026, x45028, x45029, x45031, x45032, x45033, x45035, x45036;
  wire x45037, x45039, x45040, x45041, x45042, x45043, x45044, x45046;
  wire x45047, x45048, x45050, x45051, x45052, x45054, x45055, x45056;
  wire x45058, x45059, x45060, x45061, x45063, x45064, x45065, x45067;
  wire x45068, x45069, x45070, x45072, x45073, x45074, x45076, x45077;
  wire x45078, x45079, x45081, x45082, x45083, x45085, x45086, x45087;
  wire x45088, x45090, x45091, x45092, x45094, x45095, x45096, x45097;
  wire x45100, x45102, x45103, x45105, x45106, x45107, x45109, x45110;
  wire x45111, x45112, x45115, x45117, x45118, x45120, x45121, x45122;
  wire x45124, x45125, x45126, x45127, x45130, x45132, x45133, x45135;
  wire x45136, x45137, x45139, x45140, x45141, x45142, x45145, x45147;
  wire x45148, x45150, x45151, x45152, x45154, x45155, x45156, x45157;
  wire x45160, x45162, x45163, x45165, x45166, x45167, x45169, x45170;
  wire x45171, x45172, x45175, x45178, x45179, x45181, x45182, x45183;
  wire x45185, x45186, x45187, x45188, x45191, x45194, x45195, x45197;
  wire x45198, x45199, x45201, x45202, x45203, x45204, x45207, x45210;
  wire x45211, x45213, x45214, x45215, x45217, x45218, x45219, x45220;
  wire x45223, x45226, x45227, x45229, x45230, x45231, x45233, x45234;
  wire x45235, x45236, x45239, x45242, x45243, x45245, x45246, x45247;
  wire x45249, x45250, x45251, x45252, x45255, x45258, x45259, x45261;
  wire x45262, x45263, x45265, x45266, x45267, x45268, x45271, x45274;
  wire x45275, x45277, x45278, x45279, x45281, x45282, x45283, x45284;
  wire x45287, x45290, x45291, x45293, x45294, x45295, x45297, x45298;
  wire x45299, x45300, x45303, x45306, x45307, x45309, x45310, x45311;
  wire x45313, x45314, x45315, x45316, x45319, x45322, x45323, x45325;
  wire x45326, x45327, x45329, x45330, x45331, x45332, x45335, x45338;
  wire x45339, x45341, x45342, x45343, x45345, x45346, x45347, x45348;
  wire x45351, x45354, x45355, x45357, x45358, x45359, x45361, x45362;
  wire x45363, x45364, x45367, x45370, x45371, x45373, x45374, x45375;
  wire x45377, x45378, x45379, x45380, x45383, x45386, x45387, x45389;
  wire x45390, x45391, x45393, x45394, x45395, x45397, x45398, x45399;
  wire x45400, x45401, x45402, x45403, x45404, x45405, x45407, x45408;
  wire x45409, x45412, x45413, x45414, x45417, x45418, x45419, x45422;
  wire x45423, x45424, x45427, x45428, x45429, x45431, x45433, x45434;
  wire x45436, x45437, x45438, x45440, x45441, x45443, x45444, x45446;
  wire x45447, x45448, x45450, x45451, x45453, x45454, x45456, x45457;
  wire x45458, x45460, x45461, x45463, x45464, x45466, x45467, x45468;
  wire x45470, x45471, x45473, x45474, x45476, x45477, x45478, x45480;
  wire x45481, x45483, x45484, x45486, x45487, x45488, x45490, x45491;
  wire x45493, x45494, x45496, x45497, x45498, x45500, x45501, x45503;
  wire x45504, x45506, x45507, x45508, x45510, x45511, x45513, x45514;
  wire x45516, x45517, x45518, x45520, x45521, x45523, x45524, x45526;
  wire x45527, x45528, x45530, x45531, x45533, x45534, x45536, x45537;
  wire x45538, x45540, x45541, x45543, x45544, x45546, x45547, x45548;
  wire x45550, x45551, x45553, x45554, x45556, x45557, x45558, x45560;
  wire x45561, x45563, x45564, x45566, x45567, x45568, x45570, x45571;
  wire x45573, x45574, x45576, x45577, x45578, x45580, x45581, x45583;
  wire x45584, x45586, x45587, x45588, x45590, x45591, x45593, x45594;
  wire x45596, x45597, x45598, x45600, x45601, x45603, x45604, x45606;
  wire x45607, x45608, x45610, x45611, x45613, x45614, x45616, x45617;
  wire x45618, x45620, x45621, x45622, x45624, x45625, x45626, x45627;
  wire x45628, x45629, x45630, x45632, x45633, x45634, x45636, x45637;
  wire x45638, x45640, x45641, x45642, x45644, x45645, x45646, x45647;
  wire x45649, x45650, x45651, x45653, x45654, x45655, x45656, x45658;
  wire x45659, x45660, x45662, x45663, x45664, x45665, x45667, x45668;
  wire x45669, x45671, x45672, x45673, x45674, x45676, x45677, x45678;
  wire x45680, x45681, x45682, x45683, x45685, x45686, x45687, x45689;
  wire x45690, x45691, x45692, x45694, x45695, x45696, x45698, x45699;
  wire x45701, x45702, x45704, x45705, x45706, x45708, x45709, x45711;
  wire x45712, x45714, x45715, x45716, x45718, x45719, x45721, x45722;
  wire x45724, x45725, x45726, x45728, x45729, x45731, x45732, x45734;
  wire x45735, x45736, x45738, x45739, x45741, x45742, x45744, x45745;
  wire x45746, x45748, x45749, x45751, x45752, x45754, x45755, x45756;
  wire x45758, x45759, x45761, x45762, x45764, x45765, x45766, x45768;
  wire x45769, x45771, x45772, x45774, x45775, x45776, x45778, x45779;
  wire x45781, x45782, x45784, x45785, x45786, x45788, x45789, x45791;
  wire x45792, x45794, x45795, x45796, x45798, x45799, x45801, x45802;
  wire x45804, x45805, x45806, x45808, x45809, x45811, x45812, x45814;
  wire x45815, x45816, x45818, x45819, x45821, x45822, x45824, x45825;
  wire x45826, x45828, x45829, x45831, x45832, x45834, x45835, x45836;
  wire x45838, x45839, x45841, x45842, x45844, x45845, x45846, x45848;
  wire x45849, x45851, x45852, x45854, x45855, x45856, x45858, x45859;
  wire x45861, x45862, x45864, x45865, x45866, x45868, x45869, x45871;
  wire x45872, x45874, x45875, x45876, x45878, x45880, x45881, x45882;
  wire x45883, x45884, x45886, x45887, x45888, x45890, x45892, x45893;
  wire x45895, x45897, x45898, x45900, x45902, x45903, x45905, x45907;
  wire x45908, x45910, x45912, x45913, x45915, x45917, x45918, x45920;
  wire x45922, x45923, x45925, x45927, x45928, x45930, x45932, x45933;
  wire x45935, x45937, x45938, x45940, x45942, x45943, x45945, x45947;
  wire x45948, x45950, x45952, x45953, x45955, x45957, x45958, x45960;
  wire x45962, x45963, x45965, x45967, x45968, x45970, x45972, x45973;
  wire x45975, x45977, x45978, x45980, x45982, x45983, x45985, x45987;
  wire x45988, x45990, x45992, x45993, x45995, x45997, x45998, x46000;
  wire x46002, x46003, x46005, x46007, x46008, x46035, x46036, x46037;
  wire x46038, x46039, x46041, x46042, x46043, x46045, x46046, x46047;
  wire x46049, x46050, x46051, x46053, x46054, x46055, x46057, x46058;
  wire x46059, x46061, x46062, x46063, x46065, x46066, x46067, x46069;
  wire x46070, x46071, x46073, x46074, x46075, x46077, x46078, x46079;
  wire x46081, x46082, x46083, x46085, x46086, x46087, x46089, x46090;
  wire x46091, x46093, x46094, x46095, x46097, x46098, x46099, x46101;
  wire x46102, x46103, x46105, x46106, x46107, x46109, x46110, x46111;
  wire x46113, x46114, x46115, x46117, x46118, x46119, x46121, x46122;
  wire x46123, x46125, x46126, x46127, x46129, x46130, x46131, x46134;
  wire x46136, x46137, x46139, x46140, x46142, x46143, x46145, x46147;
  wire x46148, x46150, x46152, x46153, x46155, x46157, x46158, x46160;
  wire x46162, x46163, x46165, x46167, x46168, x46170, x46172, x46173;
  wire x46175, x46177, x46178, x46180, x46182, x46183, x46185, x46187;
  wire x46188, x46190, x46192, x46193, x46195, x46197, x46198, x46200;
  wire x46202, x46203, x46205, x46207, x46208, x46210, x46212, x46213;
  wire x46215, x46217, x46218, x46220, x46222, x46223, x46225, x46227;
  wire x46228, x46230, x46232, x46233, x46235, x46237, x46238, x46240;
  wire x46242, x46243, x46245, x46247, x46248, x46252, x46254, x46255;
  wire x46257, x46258, x46260, x46261, x46263, x46264, x46266, x46267;
  wire x46269, x46271, x46272, x46274, x46276, x46277, x46279, x46281;
  wire x46282, x46284, x46286, x46287, x46289, x46291, x46292, x46294;
  wire x46296, x46297, x46299, x46301, x46302, x46304, x46306, x46307;
  wire x46309, x46311, x46312, x46314, x46316, x46317, x46319, x46321;
  wire x46322, x46324, x46326, x46327, x46329, x46331, x46332, x46334;
  wire x46336, x46337, x46339, x46341, x46342, x46344, x46346, x46347;
  wire x46349, x46351, x46352, x46358, x46360, x46361, x46363, x46364;
  wire x46366, x46367, x46369, x46370, x46372, x46373, x46375, x46376;
  wire x46378, x46379, x46381, x46382, x46384, x46385, x46387, x46389;
  wire x46390, x46392, x46394, x46395, x46397, x46399, x46400, x46402;
  wire x46404, x46405, x46407, x46409, x46410, x46412, x46414, x46415;
  wire x46417, x46419, x46420, x46422, x46424, x46425, x46427, x46429;
  wire x46430, x46438, x46440, x46441, x46443, x46444, x46446, x46447;
  wire x46449, x46450, x46452, x46453, x46455, x46456, x46458, x46459;
  wire x46461, x46462, x46464, x46465, x46467, x46468, x46469, x46471;
  wire x46472, x46473, x46475, x46476, x46477, x46479, x46480, x46481;
  wire x46483, x46484, x46485, x46487, x46488, x46489, x46491, x46492;
  wire x46493, x46495, x46496, x46497, x46499, x46501, x46502, x46504;
  wire x46506, x46507, x46509, x46510, x46511, x46513, x46514, x46515;
  wire x46517, x46518, x46519, x46521, x46522, x46523, x46525, x46526;
  wire x46527, x46529, x46530, x46531, x46533, x46535, x46536, x46538;
  wire x46540, x46541, x46543, x46545, x46546, x46548, x46550, x46551;
  wire x46553, x46555, x46556, x46558, x46560, x46561, x46563, x46565;
  wire x46566, x46568, x46570, x46571, x46573, x46575, x46576, x46578;
  wire x46580, x46581, x46583, x46585, x46587, x46589, x46591, x46593;
  wire x46595, x46597, x46599, x46601, x46603, x46605, x46607, x46609;
  wire x46611, x46613, x46615, x46617, x46619, x46621, x46623, x46625;
  wire x46627, x46629, x46631, x46633, x46635, x46637, x46639, x46641;
  wire x46643, x46644, x46646, x46648, x46650, x46652, x46654, x46656;
  wire x46658, x46660, x46662, x46664, x46666, x46668, x46670, x46672;
  wire x46674, x46676, x46678, x46680, x46682, x46684, x46686, x46688;
  wire x46690, x46692, x46694, x46696, x46698, x46700, x46701, x46702;
  wire x46703, x46705, x46707, x46709, x46711, x46713, x46715, x46717;
  wire x46719, x46721, x46723, x46725, x46727, x46729, x46731, x46733;
  wire x46735, x46737, x46739, x46741, x46743, x46745, x46747, x46749;
  wire x46751, x46752, x46753, x46754, x46755, x46756, x46757, x46758;
  wire x46759, x46761, x46763, x46765, x46767, x46769, x46771, x46773;
  wire x46775, x46777, x46779, x46781, x46783, x46785, x46787, x46789;
  wire x46790, x46791, x46792, x46793, x46794, x46795, x46796, x46797;
  wire x46798, x46799, x46800, x46801, x46802, x46803, x46804, x46805;
  wire x46807, x46808, x46809, x46811, x46812, x46813, x46815, x46816;
  wire x46817, x46819, x46820, x46821, x46823, x46824, x46825, x46827;
  wire x46828, x46829, x46831, x46832, x46833, x46835, x46836, x46837;
  wire x46839, x46840, x46841, x46843, x46844, x46845, x46847, x46848;
  wire x46849, x46851, x46852, x46853, x46855, x46856, x46857, x46859;
  wire x46860, x46861, x46863, x46864, x46865, x46867, x46868, x46869;
  wire x46871, x46872, x46873, x46875, x46876, x46877, x46879, x46880;
  wire x46881, x46883, x46884, x46885, x46887, x46888, x46889, x46891;
  wire x46892, x46893, x46895, x46896, x46897, x46899, x46900, x46901;
  wire x46903, x46904, x46905, x46907, x46908, x46909, x46911, x46912;
  wire x46913, x46915, x46916, x46917, x46919, x46920, x46921, x46923;
  wire x46924, x46925, x46928, x46930, x46932, x46934, x46936, x46938;
  wire x46940, x46942, x46944, x46946, x46948, x46950, x46952, x46954;
  wire x46956, x46958, x46960, x46961, x46962, x46963, x46964, x46965;
  wire x46966, x46967, x46968, x46969, x46970, x46971, x46972, x46973;
  wire x46974, x46975, x46976, x46977, x46978, x46979, x46980, x46981;
  wire x46982, x46983, x46984, x46985, x46986, x46987, x46988, x46989;
  wire x46990, x46991, x46992, x46994, x46996, x46998, x47000, x47002;
  wire x47004, x47006, x47008, x47010, x47012, x47014, x47016, x47018;
  wire x47020, x47022, x47024, x47026, x47028, x47030, x47032, x47034;
  wire x47036, x47038, x47040, x47042, x47044, x47046, x47048, x47050;
  wire x47052, x47054, x47056, x47057, x47058, x47059, x47060, x47061;
  wire x47062, x47063, x47064, x47065, x47066, x47067, x47068, x47069;
  wire x47070, x47071, x47072, x47073, x47074, x47075, x47076, x47077;
  wire x47078, x47079, x47080, x47081, x47082, x47083, x47084, x47085;
  wire x47086, x47087, x47088, x47089, x47090, x47091, x47092, x47093;
  wire x47094, x47095, x47096, x47097, x47098, x47099, x47100, x47101;
  wire x47102, x47103, x47104, x47105, x47106, x47107, x47108, x47109;
  wire x47110, x47111, x47112, x47113, x47114, x47115, x47116, x47117;
  wire x47118, x47119, x47120, x47121, x47122, x47123, x47124, x47125;
  wire x47126, x47127, x47128, x47129, x47130, x47131, x47132, x47133;
  wire x47134, x47135, x47136, x47137, x47138, x47139, x47140, x47141;
  wire x47142, x47143, x47144, x47145, x47146, x47147, x47148, x47149;
  wire x47150, x47151, x47152, x47153, x47154, x47155, x47156, x47157;
  wire x47158, x47159, x47160, x47161, x47162, x47163, x47164, x47165;
  wire x47166, x47167, x47168, x47169, x47170, x47171, x47172, x47173;
  wire x47174, x47175, x47176, x47177, x47178, x47179, x47180, x47181;
  wire x47182, x47183, x47184, x47185, x47186, x47187, x47188, x47189;
  wire x47190, x47191, x47192, x47193, x47194, x47195, x47196, x47197;
  wire x47198, x47199, x47200, x47201, x47202, x47203, x47204, x47205;
  wire x47206, x47207, x47208, x47209, x47210, x47211, x47212, x47213;
  wire x47214, x47215, x47216, x47217, x47218, x47219, x47220, x47221;
  wire x47222, x47223, x47224, x47225, x47226, x47227, x47228, x47229;
  wire x47230, x47231, x47232, x47233, x47234, x47235, x47236, x47237;
  wire x47238, x47239, x47240, x47241, x47242, x47243, x47244, x47245;
  wire x47246, x47247, x47248, x47249, x47250, x47251, x47252, x47253;
  wire x47254, x47255, x47256, x47257, x47258, x47259, x47260, x47261;
  wire x47262, x47263, x47264, x47265, x47266, x47267, x47268, x47269;
  wire x47270, x47271, x47272, x47273, x47274, x47275, x47276, x47277;
  wire x47278, x47279, x47280, x47281, x47282, x47283, x47284, x47285;
  wire x47286, x47287, x47288, x47289, x47290, x47291, x47292, x47293;
  wire x47294, x47295, x47296, x47297, x47298, x47299, x47300, x47301;
  wire x47302, x47303, x47304, x47305, x47306, x47307, x47308, x47309;
  wire x47310, x47311, x47312, x47313, x47314, x47315, x47316, x47317;
  wire x47318, x47319, x47320, x47321, x47322, x47323, x47324, x47325;
  wire x47326, x47327, x47328, x47329, x47330, x47331, x47332, x47333;
  wire x47334, x47335, x47336, x47337, x47338, x47339, x47340, x47341;
  wire x47342, x47343, x47344, x47345, x47346, x47347, x47348, x47349;
  wire x47350, x47351, x47352, x47353, x47354, x47355, x47356, x47357;
  wire x47358, x47359, x47360, x47361, x47362, x47363, x47364, x47365;
  wire x47366, x47367, x47368, x47369, x47370, x47371, x47372, x47373;
  wire x47374, x47375, x47376, x47377, x47378, x47379, x47380, x47381;
  wire x47382, x47383, x47384, x47385, x47386, x47387, x47388, x47389;
  wire x47390, x47391, x47392, x47393, x47394, x47395, x47396, x47397;
  wire x47398, x47399, x47400, x47401, x47402, x47403, x47404, x47405;
  wire x47406, x47407, x47408, x47409, x47410, x47411, x47412, x47413;
  wire x47414, x47415, x47416, x47417, x47418, x47419, x47420, x47421;
  wire x47422, x47423, x47424, x47425, x47426, x47427, x47428, x47429;
  wire x47430, x47431, x47432, x47433, x47434, x47435, x47436, x47437;
  wire x47438, x47439, x47440, x47441, x47442, x47443, x47444, x47445;
  wire x47446, x47447, x47448, x47449, x47450, x47451, x47452, x47453;
  wire x47454, x47455, x47456, x47457, x47458, x47459, x47460, x47461;
  wire x47462, x47463, x47464, x47465, x47466, x47467, x47468, x47469;
  wire x47470, x47471, x47472, x47473, x47474, x47475, x47476, x47477;
  wire x47478, x47479, x47480, x47481, x47482, x47483, x47484, x47485;
  wire x47486, x47487, x47488, x47489, x47490, x47491, x47492, x47493;
  wire x47494, x47495, x47496, x47497, x47498, x47499, x47500, x47501;
  wire x47502, x47503, x47504, x47505, x47506, x47507, x47508, x47509;
  wire x47510, x47511, x47512, x47513, x47514, x47515, x47516, x47517;
  wire x47518, x47519, x47520, x47521, x47522, x47523, x47524, x47525;
  wire x47526, x47527, x47528, x47529, x47530, x47531, x47532, x47533;
  wire x47534, x47535, x47536, x47537, x47538, x47539, x47540, x47541;
  wire x47542, x47543, x47544, x47545, x47546, x47547, x47548, x47549;
  wire x47550, x47551, x47552, x47553, x47554, x47555, x47556, x47557;
  wire x47558, x47559, x47560, x47561, x47562, x47563, x47564, x47565;
  wire x47566, x47567, x47568, x47569, x47570, x47571, x47572, x47573;
  wire x47574, x47575, x47576, x47577, x47578, x47579, x47580, x47581;
  wire x47582, x47583, x47584, x47585, x47586, x47587, x47588, x47589;
  wire x47590, x47591, x47592, x47593, x47594, x47595, x47596, x47597;
  wire x47598, x47599, x47600, x47601, x47602, x47603, x47604, x47605;
  wire x47606, x47607, x47608, x47609, x47610, x47611, x47612, x47613;
  wire x47614, x47615, x47616, x47617, x47618, x47619, x47620, x47621;
  wire x47622, x47623, x47624, x47625, x47626, x47627, x47628, x47629;
  wire x47630, x47631, x47632, x47633, x47634, x47635, x47636, x47637;
  wire x47638, x47639, x47640, x47641, x47642, x47643, x47644, x47645;
  wire x47646, x47647, x47648, x47649, x47650, x47651, x47652, x47653;
  wire x47654, x47655, x47656, x47657, x47658, x47659, x47660, x47661;
  wire x47662, x47663, x47664, x47665, x47666, x47667, x47668, x47669;
  wire x47670, x47671, x47672, x47673, x47674, x47675, x47676, x47677;
  wire x47678, x47679, x47680, x47681, x47682, x47683, x47684, x47685;
  wire x47686, x47687, x47688, x47689, x47690, x47691, x47692, x47693;
  wire x47694, x47695, x47696, x47697, x47698, x47699, x47700, x47701;
  wire x47702, x47703, x47704, x47705, x47706, x47707, x47708, x47709;
  wire x47710, x47711, x47712, x47713, x47714, x47715, x47716, x47717;
  wire x47718, x47719, x47720, x47721, x47722, x47723, x47724, x47725;
  wire x47726, x47727, x47728, x47729, x47730, x47731, x47732, x47733;
  wire x47734, x47735, x47736, x47737, x47738, x47739, x47740, x47741;
  wire x47742, x47743, x47744, x47745, x47746, x47747, x47748, x47749;
  wire x47750, x47751, x47752, x47753, x47754, x47755, x47756, x47757;
  wire x47758, x47759, x47760, x47761, x47762, x47763, x47764, x47765;
  wire x47766, x47767, x47768, x47769, x47770, x47771, x47772, x47773;
  wire x47774, x47775, x47776, x47777, x47778, x47779, x47780, x47781;
  wire x47782, x47783, x47784, x47785, x47786, x47787, x47788, x47789;
  wire x47790, x47791, x47792, x47793, x47794, x47795, x47796, x47797;
  wire x47798, x47799, x47800, x47801, x47802, x47803, x47804, x47805;
  wire x47806, x47807, x47808, x47809, x47810, x47811, x47812, x47813;
  wire x47814, x47815, x47816, x47817, x47818, x47819, x47820, x47821;
  wire x47822, x47823, x47824, x47825, x47826, x47827, x47828, x47829;
  wire x47830, x47831, x47832, x47833, x47834, x47835, x47836, x47837;
  wire x47838, x47839, x47840, x47841, x47842, x47843, x47844, x47845;
  wire x47846, x47847, x47848, x47849, x47850, x47851, x47852, x47853;
  wire x47854, x47855, x47856, x47857, x47858, x47859, x47860, x47861;
  wire x47862, x47863, x47864, x47865, x47866, x47867, x47868, x47869;
  wire x47870, x47871, x47872, x47873, x47874, x47875, x47876, x47877;
  wire x47878, x47879, x47880, x47881, x47882, x47883, x47884, x47885;
  wire x47886, x47887, x47888, x47889, x47890, x47891, x47892, x47893;
  wire x47894, x47895, x47896, x47897, x47898, x47899, x47900, x47901;
  wire x47902, x47903, x47904, x47905, x47906, x47907, x47908, x47909;
  wire x47910, x47911, x47912, x47913, x47914, x47915, x47916, x47917;
  wire x47918, x47919, x47920, x47921, x47922, x47923, x47924, x47925;
  wire x47926, x47927, x47928, x47929, x47930, x47931, x47932, x47933;
  wire x47934, x47935, x47936, x47937, x47938, x47939, x47940, x47941;
  wire x47942, x47943, x47944, x47945, x47946, x47947, x47948, x47949;
  wire x47950, x47951, x47952, x47953, x47954, x47955, x47956, x47957;
  wire x47958, x47959, x47960, x47961, x47962, x47963, x47964, x47965;
  wire x47966, x47967, x47968, x47969, x47970, x47971, x47972, x47973;
  wire x47974, x47975, x47976, x47977, x47978, x47979, x47980, x47981;
  wire x47982, x47983, x47984, x47985, x47986, x47987, x47988, x47989;
  wire x47990, x47991, x47992, x47993, x47994, x47995, x47996, x47997;
  wire x47998, x47999, x48000, x48001, x48002, x48003, x48004, x48005;
  wire x48006, x48007, x48008, x48009, x48010, x48011, x48012, x48013;
  wire x48014, x48015, x48016, x48017, x48018, x48019, x48020, x48021;
  wire x48022, x48023, x48024, x48025, x48026, x48027, x48028, x48029;
  wire x48030, x48031, x48032, x48033, x48034, x48035, x48036, x48037;
  wire x48038, x48039, x48040, x48041, x48042, x48043, x48044, x48045;
  wire x48046, x48047, x48048, x48049, x48050, x48051, x48052, x48053;
  wire x48054, x48055, x48056, x48057, x48058, x48059, x48060, x48061;
  wire x48062, x48063, x48064, x48065, x48066, x48067, x48068, x48069;
  wire x48070, x48071, x48072, x48073, x48074, x48075, x48076, x48077;
  wire x48078, x48079, x48080, x48081, x48082, x48083, x48084, x48085;
  wire x48086, x48087, x48088, x48089, x48090, x48091, x48092, x48093;
  wire x48094, x48095, x48096, x48097, x48098, x48099, x48100, x48101;
  wire x48102, x48103, x48104, x48105, x48106, x48107, x48108, x48109;
  wire x48110, x48111, x48112, x48113, x48114, x48115, x48116, x48117;
  wire x48118, x48119, x48120, x48121, x48122, x48123, x48124, x48125;
  wire x48126, x48127, x48128, x48129, x48130, x48131, x48132, x48133;
  wire x48134, x48135, x48136, x48137, x48138, x48139, x48140, x48141;
  wire x48142, x48143, x48144, x48145, x48146, x48147, x48148, x48149;
  wire x48150, x48151, x48152, x48153, x48154, x48155, x48156, x48157;
  wire x48158, x48159, x48160, x48161, x48162, x48163, x48164, x48165;
  wire x48166, x48167, x48168, x48169, x48170, x48171, x48172, x48173;
  wire x48174, x48175, x48176, x48177, x48178, x48179, x48180, x48181;
  wire x48182, x48183, x48184, x48185, x48186, x48187, x48188, x48189;
  wire x48190, x48191, x48192, x48193, x48194, x48195, x48196, x48197;
  wire x48198, x48199, x48200, x48201, x48202, x48203, x48204, x48205;
  wire x48206, x48207, x48208, x48209, x48210, x48211, x48212, x48213;
  wire x48214, x48215, x48216, x48217, x48218, x48219, x48220, x48221;
  wire x48222, x48223, x48224, x48225, x48226, x48227, x48228, x48229;
  wire x48230, x48231, x48232, x48233, x48234, x48235, x48236, x48237;
  wire x48238, x48239, x48240, x48241, x48242, x48243, x48244, x48245;
  wire x48246, x48247, x48248, x48249, x48250, x48251, x48252, x48253;
  wire x48254, x48255, x48256, x48257, x48258, x48259, x48260, x48261;
  wire x48262, x48263, x48264, x48265, x48266, x48267, x48268, x48269;
  wire x48270, x48271, x48272, x48273, x48274, x48275, x48276, x48277;
  wire x48278, x48279, x48280, x48281, x48282, x48283, x48284, x48285;
  wire x48286, x48287, x48288, x48289, x48290, x48291, x48292, x48293;
  wire x48294, x48295, x48296, x48297, x48298, x48299, x48300, x48301;
  wire x48302, x48303, x48304, x48305, x48306, x48307, x48308, x48309;
  wire x48310, x48311, x48312, x48313, x48314, x48315, x48316, x48317;
  wire x48318, x48319, x48320, x48321, x48322, x48323, x48324, x48325;
  wire x48326, x48327, x48328, x48329, x48330, x48331, x48332, x48333;
  wire x48334, x48335, x48336, x48337, x48338, x48339, x48340, x48341;
  wire x48342, x48343, x48344, x48345, x48346, x48347, x48348, x48349;
  wire x48350, x48351, x48352, x48353, x48354, x48355, x48356, x48357;
  wire x48358, x48359, x48360, x48361, x48362, x48363, x48364, x48365;
  wire x48366, x48367, x48368, x48369, x48370, x48371, x48372, x48373;
  wire x48374, x48375, x48376, x48377, x48378, x48379, x48380, x48381;
  wire x48382, x48383, x48384, x48385, x48386, x48387, x48388, x48389;
  wire x48390, x48391, x48392, x48393, x48394, x48395, x48396, x48397;
  wire x48398, x48399, x48400, x48401, x48402, x48403, x48404, x48405;
  wire x48406, x48407, x48408, x48409, x48410, x48411, x48412, x48413;
  wire x48414, x48415, x48416, x48417, x48418, x48419, x48420, x48421;
  wire x48422, x48423, x48424, x48425, x48426, x48427, x48428, x48429;
  wire x48430, x48431, x48432, x48433, x48434, x48435, x48436, x48437;
  wire x48438, x48439, x48440, x48441, x48442, x48443, x48444, x48445;
  wire x48446, x48447, x48448, x48449, x48450, x48451, x48452, x48453;
  wire x48454, x48455, x48456, x48457, x48458, x48459, x48460, x48461;
  wire x48462, x48463, x48464, x48465, x48466, x48467, x48468, x48469;
  wire x48470, x48471, x48472, x48473, x48474, x48475, x48476, x48477;
  wire x48478, x48479, x48480, x48481, x48482, x48483, x48484, x48485;
  wire x48486, x48487, x48488, x48489, x48490, x48491, x48492, x48493;
  wire x48494, x48495, x48496, x48497, x48498, x48499, x48500, x48501;
  wire x48502, x48503, x48504, x48505, x48506, x48507, x48508, x48509;
  wire x48510, x48511, x48512, x48513, x48514, x48515, x48516, x48517;
  wire x48518, x48519, x48520, x48521, x48522, x48523, x48524, x48525;
  wire x48526, x48527, x48528, x48529, x48530, x48531, x48532, x48533;
  wire x48534, x48535, x48536, x48537, x48538, x48539, x48540, x48541;
  wire x48542, x48543, x48544, x48545, x48546, x48547, x48548, x48549;
  wire x48550, x48551, x48552, x48553, x48554, x48555, x48556, x48557;
  wire x48558, x48559, x48560, x48561, x48562, x48563, x48564, x48565;
  wire x48566, x48567, x48568, x48569, x48570, x48571, x48572, x48573;
  wire x48574, x48575, x48576, x48577, x48578, x48579, x48580, x48581;
  wire x48582, x48583, x48584, x48585, x48586, x48587, x48588, x48589;
  wire x48590, x48591, x48592, x48593, x48594, x48595, x48596, x48597;
  wire x48598, x48599, x48600, x48601, x48602, x48603, x48604, x48605;
  wire x48606, x48607, x48608, x48609, x48610, x48611, x48612, x48613;
  wire x48614, x48615, x48616, x48617, x48618, x48619, x48620, x48621;
  wire x48622, x48623, x48624, x48625, x48626, x48627, x48628, x48629;
  wire x48630, x48631, x48632, x48633, x48634, x48635, x48636, x48637;
  wire x48638, x48639, x48640, x48641, x48642, x48643, x48644, x48645;
  wire x48646, x48647, x48648, x48649, x48650, x48651, x48652, x48653;
  wire x48654, x48655, x48656, x48657, x48658, x48659, x48660, x48661;
  wire x48662, x48663, x48664, x48665, x48666, x48667, x48668, x48669;
  wire x48670, x48671, x48672, x48673, x48674, x48675, x48676, x48677;
  wire x48678, x48679, x48680, x48681, x48682, x48683, x48684, x48685;
  wire x48686, x48687, x48688, x48689, x48690, x48691, x48692, x48693;
  wire x48694, x48695, x48696, x48697, x48698, x48699, x48700, x48701;
  wire x48702, x48703, x48704, x48705, x48706, x48707, x48708, x48709;
  wire x48710, x48711, x48712, x48713, x48714, x48715, x48716, x48717;
  wire x48718, x48719, x48720, x48721, x48722, x48723, x48724, x48725;
  wire x48726, x48727, x48728, x48729, x48730, x48731, x48732, x48733;
  wire x48734, x48735, x48736, x48737, x48738, x48739, x48740, x48741;
  wire x48742, x48743, x48744, x48745, x48746, x48747, x48748, x48749;
  wire x48750, x48751, x48752, x48753, x48754, x48755, x48756, x48757;
  wire x48758, x48759, x48760, x48761, x48762, x48763, x48764, x48765;
  wire x48766, x48767, x48768, x48769, x48770, x48771, x48772, x48773;
  wire x48774, x48775, x48776, x48777, x48778, x48779, x48780, x48781;
  wire x48782, x48783, x48784, x48785, x48786, x48787, x48788, x48789;
  wire x48790, x48791, x48792, x48793, x48794, x48795, x48796, x48797;
  wire x48798, x48799, x48800, x48801, x48802, x48803, x48804, x48805;
  wire x48806, x48807, x48808, x48809, x48810, x48811, x48812, x48813;
  wire x48814, x48815, x48816, x48817, x48818, x48819, x48820, x48821;
  wire x48822, x48823, x48824, x48825, x48826, x48827, x48828, x48829;
  wire x48830, x48831, x48832, x48833, x48834, x48835, x48836, x48837;
  wire x48838, x48839, x48840, x48841, x48842, x48843, x48844, x48845;
  wire x48846, x48847, x48848, x48849, x48850, x48851, x48852, x48853;
  wire x48854, x48855, x48856, x48857, x48858, x48859, x48860, x48861;
  wire x48862, x48863, x48864, x48865, x48866, x48867, x48868, x48869;
  wire x48870, x48871, x48872, x48873, x48874, x48875, x48876, x48877;
  wire x48878, x48879, x48880, x48881, x48882, x48883, x48884, x48885;
  wire x48886, x48887, x48888, x48889, x48890, x48891, x48892, x48893;
  wire x48894, x48895, x48896, x48897, x48898, x48899, x48900, x48901;
  wire x48902, x48903, x48904, x48905, x48906, x48907, x48908, x48909;
  wire x48910, x48911, x48912, x48913, x48914, x48915, x48916, x48917;
  wire x48918, x48919, x48920, x48921, x48922, x48923, x48924, x48925;
  wire x48926, x48927, x48928, x48929, x48930, x48931, x48932, x48933;
  wire x48934, x48935, x48936, x48937, x48938, x48939, x48940, x48941;
  wire x48942, x48943, x48944, x48945, x48946, x48947, x48948, x48949;
  wire x48950, x48951, x48952, x48953, x48954, x48955, x48956, x48957;
  wire x48958, x48959, x48960, x48961, x48962, x48963, x48964, x48965;
  wire x48966, x48967, x48968, x48969, x48970, x48971, x48972, x48973;
  wire x48974, x48975, x48976, x48977, x48978, x48979, x48980, x48981;
  wire x48982, x48983, x48984, x48985, x48986, x48987, x48988, x48989;
  wire x48990, x48991, x48992, x48993, x48994, x48995, x48996, x48997;
  wire x48998, x48999, x49000, x49001, x49002, x49003, x49004, x49005;
  wire x49006, x49007, x49008, x49009, x49010, x49011, x49012, x49013;
  wire x49014, x49015, x49016, x49017, x49018, x49019, x49020, x49021;
  wire x49022, x49023, x49024, x49025, x49026, x49027, x49028, x49029;
  wire x49030, x49031, x49032, x49033, x49034, x49035, x49036, x49037;
  wire x49038, x49039, x49040, x49041, x49042, x49043, x49044, x49045;
  wire x49046, x49047, x49048, x49049, x49050, x49051, x49052, x49053;
  wire x49054, x49055, x49056, x49057, x49058, x49059, x49060, x49061;
  wire x49062, x49063, x49064, x49065, x49066, x49067, x49068, x49069;
  wire x49070, x49071, x49072, x49073, x49074, x49075, x49076, x49077;
  wire x49078, x49079, x49080, x49081, x49082, x49083, x49084, x49085;
  wire x49086, x49087, x49088, x49089, x49090, x49091, x49092, x49093;
  wire x49094, x49095, x49096, x49097, x49098, x49099, x49100, x49101;
  wire x49102, x49103, x49104, x49105, x49106, x49107, x49108, x49109;
  wire x49110, x49111, x49112, x49113, x49114, x49115, x49116, x49117;
  wire x49118, x49119, x49120, x49121, x49122, x49123, x49124, x49125;
  wire x49126, x49127, x49128, x49129, x49130, x49131, x49132, x49133;
  wire x49134, x49135, x49136, x49137, x49138, x49139, x49140, x49141;
  wire x49142, x49143, x49144, x49145, x49146, x49147, x49148, x49149;
  wire x49150, x49151, x49152, x49153, x49154, x49155, x49156, x49157;
  wire x49158, x49159, x49160, x49161, x49162, x49163, x49164, x49165;
  wire x49166, x49167, x49168, x49169, x49170, x49171, x49172, x49173;
  wire x49174, x49175, x49176, x49177, x49178, x49179, x49180, x49181;
  wire x49182, x49183, x49184, x49185, x49186, x49187, x49188, x49189;
  wire x49190, x49191, x49192, x49193, x49194, x49195, x49196, x49197;
  wire x49198, x49199, x49200, x49201, x49202, x49203, x49204, x49205;
  wire x49206, x49207, x49208, x49209, x49210, x49211, x49212, x49213;
  wire x49214, x49215, x49216, x49217, x49218, x49219, x49220, x49221;
  wire x49222, x49223, x49224, x49225, x49226, x49227, x49228, x49229;
  wire x49230, x49231, x49232, x49233, x49234, x49235, x49236, x49237;
  wire x49238, x49239, x49240, x49241, x49242, x49243, x49244, x49245;
  wire x49246, x49247, x49248, x49249, x49250, x49251, x49252, x49253;
  wire x49254, x49255, x49256, x49257, x49258, x49259, x49260, x49261;
  wire x49262, x49263, x49264, x49265, x49266, x49267, x49268, x49269;
  wire x49270, x49271, x49272, x49273, x49274, x49275, x49276, x49277;
  wire x49278, x49279, x49280, x49281, x49282, x49283, x49284, x49285;
  wire x49286, x49287, x49288, x49289, x49290, x49291, x49292, x49293;
  wire x49294, x49295, x49296, x49297, x49298, x49299, x49300, x49301;
  wire x49302, x49303, x49304, x49305, x49306, x49307, x49308, x49309;
  wire x49310, x49311, x49312, x49313, x49314, x49315, x49316, x49317;
  wire x49318, x49319, x49320, x49321, x49322, x49323, x49324, x49325;
  wire x49326, x49327, x49328, x49329, x49330, x49331, x49332, x49333;
  wire x49334, x49335, x49336, x49337, x49338, x49339, x49340, x49341;
  wire x49342, x49343, x49344, x49345, x49346, x49347, x49348, x49349;
  wire x49350, x49351, x49352, x49353, x49354, x49355, x49356, x49357;
  wire x49358, x49359, x49360, x49361, x49362, x49363, x49364, x49365;
  wire x49366, x49367, x49368, x49369, x49370, x49371, x49372, x49373;
  wire x49374, x49375, x49376, x49377, x49378, x49379, x49380, x49381;
  wire x49382, x49383, x49384, x49385, x49386, x49387, x49388, x49389;
  wire x49390, x49391, x49392, x49393, x49394, x49395, x49396, x49397;
  wire x49398, x49399, x49400, x49401, x49402, x49403, x49404, x49405;
  wire x49406, x49407, x49408, x49409, x49410, x49411, x49412, x49413;
  wire x49414, x49415, x49416, x49417, x49418, x49419, x49420, x49421;
  wire x49422, x49423, x49424, x49425, x49426, x49427, x49428, x49429;
  wire x49430, x49431, x49432, x49433, x49434, x49435, x49436, x49437;
  wire x49438, x49439, x49440, x49441, x49442, x49443, x49444, x49445;
  wire x49446, x49447, x49448, x49449, x49450, x49451, x49452, x49453;
  wire x49454, x49455, x49456, x49457, x49458, x49459, x49460, x49461;
  wire x49462, x49463, x49464, x49465, x49466, x49467, x49468, x49469;
  wire x49470, x49471, x49472, x49473, x49474, x49475, x49476, x49477;
  wire x49478, x49479, x49480, x49481, x49482, x49483, x49484, x49485;
  wire x49486, x49487, x49488, x49489, x49490, x49491, x49492, x49493;
  wire x49494, x49495, x49496, x49497, x49498, x49499, x49500, x49501;
  wire x49502, x49503, x49504, x49505, x49506, x49507, x49508, x49509;
  wire x49510, x49511, x49512, x49513, x49514, x49515, x49516, x49517;
  wire x49518, x49519, x49520, x49521, x49522, x49523, x49524, x49525;
  wire x49526, x49527, x49528, x49529, x49530, x49531, x49532, x49533;
  wire x49534, x49535, x49536, x49537, x49538, x49539, x49540, x49541;
  wire x49542, x49543, x49544, x49545, x49546, x49547, x49548, x49549;
  wire x49550, x49551, x49552, x49553, x49554, x49555, x49556, x49557;
  wire x49558, x49559, x49560, x49561, x49562, x49563, x49564, x49565;
  wire x49566, x49567, x49568, x49569, x49570, x49571, x49572, x49573;
  wire x49574, x49575, x49576, x49577, x49578, x49579, x49580, x49581;
  wire x49582, x49583, x49584, x49585, x49586, x49587, x49588, x49589;
  wire x49590, x49591, x49592, x49593, x49594, x49595, x49596, x49597;
  wire x49598, x49599, x49600, x49601, x49602, x49603, x49604, x49605;
  wire x49606, x49607, x49608, x49609, x49610, x49611, x49612, x49613;
  wire x49614, x49615, x49616, x49617, x49618, x49619, x49620, x49621;
  wire x49622, x49623, x49624, x49625, x49626, x49627, x49628, x49629;
  wire x49630, x49631, x49632, x49633, x49634, x49635, x49636, x49637;
  wire x49638, x49639, x49640, x49641, x49642, x49643, x49644, x49645;
  wire x49646, x49647, x49648, x49649, x49650, x49651, x49652, x49653;
  wire x49654, x49655, x49656, x49657, x49658, x49659, x49660, x49661;
  wire x49662, x49663, x49664, x49665, x49666, x49667, x49668, x49669;
  wire x49670, x49671, x49672, x49673, x49674, x49675, x49676, x49677;
  wire x49678, x49679, x49680, x49681, x49682, x49683, x49684, x49685;
  wire x49686, x49687, x49688, x49690, x49691, x49692, x49694, x49695;
  wire x49696, x49698, x49699, x49700, x49702, x49703, x49704, x49706;
  wire x49707, x49708, x49710, x49711, x49712, x49714, x49715, x49716;
  wire x49718, x49719, x49720, x49722, x49723, x49724, x49726, x49727;
  wire x49728, x49730, x49731, x49732, x49734, x49735, x49736, x49738;
  wire x49739, x49740, x49742, x49743, x49744, x49746, x49747, x49748;
  wire x49750, x49751, x49752, x49754, x49755, x49756, x49758, x49759;
  wire x49760, x49762, x49763, x49764, x49766, x49767, x49768, x49770;
  wire x49771, x49772, x49774, x49775, x49776, x49778, x49779, x49780;
  wire x49782, x49783, x49784, x49786, x49787, x49788, x49790, x49791;
  wire x49792, x49794, x49795, x49796, x49798, x49799, x49800, x49802;
  wire x49803, x49804, x49806, x49807, x49808, x49810, x49811, x49812;
  wire x49814, x49815, x49816, x49817, x49818, x49819, x49820, x49821;
  wire x49822, x49823, x49824, x49825, x49826, x49827, x49828, x49829;
  wire x49830, x49831, x49832, x49833, x49834, x49835, x49836, x49837;
  wire x49838, x49839, x49840, x49841, x49842, x49843, x49844, x49845;
  wire x49846, x49847, x49848, x49849, x49850, x49851, x49852, x49853;
  wire x49854, x49855, x49856, x49857, x49858, x49859, x49860, x49861;
  wire x49862, x49863, x49864, x49865, x49866, x49867, x49868, x49869;
  wire x49870, x49871, x49872, x49873, x49874, x49875, x49876, x49877;
  wire x49910, x49911, x49912, x49913, x49914, x49915, x49916, x49917;
  wire x49918, x49919, x49920, x49921, x49922, x49923, x49924, x49925;
  wire x49926, x49927, x49928, x49929, x49930, x49931, x49932, x49933;
  wire x49934, x49935, x49936, x49937, x49938, x49939, x49940, x49941;
  wire x49942, x49943, x49944, x49945, x49946, x49947, x49948, x49949;
  wire x49950, x49951, x49952, x49953, x49954, x49955, x49956, x49957;
  wire x49958, x49959, x49960, x49961, x49962, x49963, x49964, x49965;
  wire x49966, x49967, x49968, x49969, x49970, x49971, x49972, x49973;
  wire x49974, x49975, x49976, x49977, x49978, x49979, x49980, x49981;
  wire x49982, x49983, x49984, x49985, x49986, x49987, x49988, x49989;
  wire x49990, x49991, x49992, x49993, x49994, x49995, x49996, x49997;
  wire x49998, x49999, x50000, x50001, x50002, x50003, x50004, x50005;
  wire x50006, x50009, x50010, x50012, x50015, x50016, x50018, x50021;
  wire x50022, x50024, x50027, x50028, x50030, x50033, x50034, x50036;
  wire x50039, x50040, x50042, x50045, x50046, x50048, x50051, x50052;
  wire x50054, x50057, x50058, x50060, x50063, x50064, x50066, x50069;
  wire x50070, x50072, x50075, x50076, x50078, x50081, x50082, x50084;
  wire x50087, x50088, x50090, x50093, x50094, x50096, x50099, x50100;
  wire x50102, x50105, x50106, x50108, x50111, x50112, x50114, x50117;
  wire x50118, x50120, x50123, x50124, x50126, x50129, x50130, x50132;
  wire x50135, x50136, x50138, x50141, x50142, x50144, x50147, x50148;
  wire x50150, x50153, x50154, x50156, x50159, x50160, x50162, x50165;
  wire x50166, x50168, x50171, x50172, x50174, x50177, x50178, x50180;
  wire x50183, x50184, x50186, x50189, x50190, x50192, x50195, x50196;
  wire x50228, x50229, x50230, x50231, x50232, x50234, x50235, x50236;
  wire x50238, x50239, x50240, x50242, x50243, x50244, x50246, x50247;
  wire x50248, x50250, x50251, x50252, x50254, x50255, x50256, x50258;
  wire x50259, x50260, x50262, x50263, x50264, x50266, x50267, x50268;
  wire x50270, x50271, x50272, x50274, x50275, x50276, x50278, x50279;
  wire x50280, x50282, x50283, x50284, x50286, x50287, x50288, x50290;
  wire x50291, x50292, x50294, x50295, x50296, x50298, x50299, x50300;
  wire x50302, x50303, x50304, x50306, x50307, x50308, x50310, x50311;
  wire x50312, x50314, x50315, x50316, x50318, x50319, x50320, x50322;
  wire x50323, x50324, x50326, x50327, x50328, x50330, x50331, x50332;
  wire x50334, x50335, x50336, x50338, x50339, x50340, x50342, x50343;
  wire x50344, x50346, x50347, x50348, x50350, x50352, x50353, x50355;
  wire x50356, x50358, x50359, x50361, x50363, x50364, x50366, x50368;
  wire x50369, x50371, x50373, x50374, x50376, x50378, x50379, x50381;
  wire x50383, x50384, x50386, x50388, x50389, x50391, x50393, x50394;
  wire x50396, x50398, x50399, x50401, x50403, x50404, x50406, x50408;
  wire x50409, x50411, x50413, x50414, x50416, x50418, x50419, x50421;
  wire x50423, x50424, x50426, x50428, x50429, x50431, x50433, x50434;
  wire x50436, x50438, x50439, x50441, x50443, x50444, x50446, x50448;
  wire x50449, x50451, x50453, x50454, x50456, x50458, x50459, x50461;
  wire x50463, x50464, x50466, x50468, x50469, x50471, x50473, x50474;
  wire x50476, x50478, x50479, x50481, x50483, x50484, x50486, x50488;
  wire x50489, x50491, x50493, x50494, x50496, x50498, x50499, x50501;
  wire x50502, x50504, x50505, x50507, x50508, x50510, x50511, x50513;
  wire x50515, x50516, x50518, x50520, x50521, x50523, x50525, x50526;
  wire x50528, x50530, x50531, x50533, x50535, x50536, x50538, x50540;
  wire x50541, x50543, x50545, x50546, x50548, x50550, x50551, x50553;
  wire x50555, x50556, x50558, x50560, x50561, x50563, x50565, x50566;
  wire x50568, x50570, x50571, x50573, x50575, x50576, x50578, x50580;
  wire x50581, x50583, x50585, x50586, x50588, x50590, x50591, x50593;
  wire x50595, x50596, x50598, x50600, x50601, x50603, x50605, x50606;
  wire x50608, x50610, x50611, x50613, x50615, x50616, x50618, x50620;
  wire x50621, x50623, x50625, x50626, x50628, x50630, x50631, x50633;
  wire x50634, x50636, x50637, x50639, x50640, x50642, x50643, x50645;
  wire x50646, x50648, x50649, x50651, x50652, x50654, x50655, x50657;
  wire x50659, x50660, x50662, x50664, x50665, x50667, x50669, x50670;
  wire x50672, x50674, x50675, x50677, x50679, x50680, x50682, x50684;
  wire x50685, x50687, x50689, x50690, x50692, x50694, x50695, x50697;
  wire x50699, x50700, x50702, x50704, x50705, x50707, x50709, x50710;
  wire x50712, x50714, x50715, x50717, x50719, x50720, x50722, x50724;
  wire x50725, x50727, x50729, x50730, x50732, x50734, x50735, x50737;
  wire x50738, x50740, x50741, x50743, x50744, x50746, x50747, x50749;
  wire x50750, x50752, x50753, x50755, x50756, x50758, x50759, x50761;
  wire x50762, x50764, x50765, x50767, x50768, x50770, x50771, x50773;
  wire x50774, x50776, x50777, x50779, x50780, x50781, x50783, x50785;
  wire x50786, x50788, x50790, x50791, x50793, x50795, x50796, x50798;
  wire x50800, x50801, x50803, x50805, x50806, x50808, x50810, x50811;
  wire x50813, x50815, x50816, x50818, x50820, x50821, x50823, x50825;
  wire x50826, x50828, x50830, x50831, x50833, x50835, x50836, x50838;
  wire x50840, x50841, x50843, x50845, x50846, x50848, x50850, x50851;
  wire x50853, x50855, x50856, x50858, x50860, x50861, x50863, x50865;
  wire x50866, x50868, x50870, x50871, x50873, x50875, x50876, x50878;
  wire x50880, x50881, x50883, x50885, x50886, x50888, x50890, x50891;
  wire x50893, x50895, x50896, x50898, x50900, x50901, x50903, x50905;
  wire x50906, x50908, x50910, x50911, x50913, x50915, x50916, x50918;
  wire x50920, x50921, x50923, x50925, x50926, x50928, x50930, x50931;
  wire x50933, x50935, x50936, x50938, x50939, x50941, x50943, x50945;
  wire x50947, x50949, x50951, x50953, x50955, x50956, x50958, x50960;
  wire x50962, x50964, x50966, x50968, x50970, x50972, x50974, x50976;
  wire x50978, x50980, x50982, x50984, x50986, x50988, x50990, x50991;
  wire x50993, x50995, x50997, x50999, x51001, x51003, x51005, x51007;
  wire x51009, x51011, x51013, x51015, x51017, x51019, x51021, x51023;
  wire x51025, x51027, x51029, x51031, x51033, x51035, x51037, x51039;
  wire x51041, x51043, x51044, x51046, x51048, x51050, x51052, x51054;
  wire x51056, x51058, x51060, x51062, x51064, x51066, x51068, x51070;
  wire x51072, x51074, x51076, x51078, x51080, x51082, x51084, x51086;
  wire x51088, x51090, x51092, x51094, x51096, x51098, x51100, x51102;
  wire x51104, x51106, x51108, x51110, x51112, x51114, x51115, x51117;
  wire x51119, x51121, x51123, x51125, x51127, x51129, x51131, x51133;
  wire x51135, x51137, x51139, x51141, x51143, x51145, x51147, x51149;
  wire x51151, x51153, x51155, x51157, x51159, x51161, x51163, x51165;
  wire x51167, x51169, x51171, x51173, x51175, x51177, x51179, x51181;
  wire x51183, x51185, x51187, x51189, x51191, x51193, x51195, x51197;
  wire x51199, x51201, x51203, x51204, x51206, x51208, x51210, x51212;
  wire x51214, x51216, x51218, x51220, x51222, x51224, x51226, x51228;
  wire x51230, x51232, x51234, x51236, x51238, x51240, x51242, x51244;
  wire x51246, x51248, x51250, x51252, x51254, x51256, x51258, x51260;
  wire x51262, x51264, x51266, x51268, x51270, x51272, x51274, x51276;
  wire x51278, x51280, x51282, x51284, x51286, x51288, x51290, x51292;
  wire x51294, x51296, x51298, x51300, x51302, x51304, x51306, x51308;
  wire x51310, x51311, x51313, x51315, x51317, x51319, x51321, x51323;
  wire x51325, x51327, x51329, x51331, x51333, x51335, x51337, x51339;
  wire x51341, x51343, x51345, x51347, x51349, x51351, x51353, x51355;
  wire x51357, x51359, x51361, x51363, x51365, x51367, x51369, x51371;
  wire x51373, x51375, x51377, x51379, x51381, x51383, x51385, x51387;
  wire x51389, x51391, x51393, x51395, x51397, x51399, x51401, x51403;
  wire x51405, x51407, x51409, x51411, x51413, x51415, x51417, x51419;
  wire x51421, x51423, x51425, x51427, x51429, x51431, x51433, x51435;
  wire x51436, x51438, x51440, x51442, x51444, x51446, x51448, x51450;
  wire x51452, x51454, x51456, x51458, x51460, x51462, x51464, x51466;
  wire x51468, x51470, x51472, x51474, x51476, x51478, x51480, x51482;
  wire x51484, x51486, x51488, x51490, x51492, x51494, x51496, x51498;
  wire x51500, x51502, x51504, x51506, x51508, x51510, x51512, x51514;
  wire x51516, x51518, x51520, x51522, x51524, x51526, x51528, x51530;
  wire x51532, x51534, x51536, x51538, x51540, x51542, x51544, x51546;
  wire x51548, x51550, x51552, x51554, x51556, x51558, x51560, x51562;
  wire x51564, x51566, x51568, x51570, x51572, x51574, x51576, x51578;
  wire x51579, x51581, x51583, x51585, x51587, x51589, x51591, x51593;
  wire x51595, x51597, x51599, x51601, x51603, x51605, x51607, x51609;
  wire x51611, x51613, x51615, x51617, x51619, x51621, x51623, x51625;
  wire x51627, x51629, x51631, x51633, x51635, x51637, x51639, x51641;
  wire x51643, x51645, x51647, x51649, x51651, x51653, x51655, x51657;
  wire x51659, x51661, x51663, x51665, x51667, x51669, x51671, x51673;
  wire x51675, x51677, x51679, x51681, x51683, x51685, x51687, x51689;
  wire x51691, x51693, x51695, x51697, x51699, x51701, x51703, x51705;
  wire x51707, x51709, x51711, x51713, x51715, x51717, x51719, x51721;
  wire x51723, x51725, x51727, x51729, x51731, x51733, x51735, x51737;
  wire x51739, x51740, x51742, x51744, x51746, x51748, x51750, x51752;
  wire x51754, x51756, x51758, x51760, x51762, x51764, x51766, x51768;
  wire x51770, x51772, x51774, x51776, x51778, x51780, x51782, x51784;
  wire x51786, x51788, x51790, x51792, x51794, x51796, x51798, x51800;
  wire x51802, x51804, x51806, x51808, x51810, x51812, x51814, x51816;
  wire x51818, x51820, x51822, x51824, x51826, x51828, x51830, x51832;
  wire x51834, x51836, x51838, x51840, x51842, x51844, x51846, x51848;
  wire x51850, x51852, x51854, x51856, x51858, x51860, x51862, x51864;
  wire x51866, x51868, x51870, x51872, x51874, x51876, x51878, x51880;
  wire x51882, x51884, x51886, x51888, x51890, x51892, x51894, x51896;
  wire x51898, x51900, x51902, x51904, x51906, x51908, x51910, x51912;
  wire x51914, x51916, x51918, x51919, x51921, x51923, x51925, x51927;
  wire x51929, x51931, x51933, x51935, x51937, x51939, x51941, x51943;
  wire x51945, x51947, x51949, x51951, x51953, x51955, x51957, x51959;
  wire x51961, x51963, x51965, x51967, x51969, x51971, x51973, x51975;
  wire x51977, x51979, x51981, x51983, x51984, x51985, x51986, x51987;
  wire x51988, x51990, x51991, x51992, x51993, x51994, x51995, x51996;
  wire x51998, x51999, x52000, x52001, x52002, x52003, x52004, x52006;
  wire x52007, x52008, x52009, x52010, x52011, x52012, x52013, x52014;
  wire x52015, x52017, x52018, x52019, x52020, x52021, x52022, x52023;
  wire x52025, x52026, x52027, x52028, x52029, x52030, x52031, x52033;
  wire x52034, x52035, x52036, x52037, x52038, x52039, x52041, x52042;
  wire x52043, x52045, x52046, x52047, x52048, x52050, x52051, x52052;
  wire x52053, x52054, x52055, x52056, x52058, x52059, x52060, x52062;
  wire x52063, x52064, x52065, x52066, x52067, x52068, x52070, x52071;
  wire x52072, x52073, x52074, x52075, x52076, x52078, x52079, x52080;
  wire x52082, x52083, x52084, x52085, x52087, x52088, x52089, x52091;
  wire x52092, x52093, x52094, x52096, x52097, x52098, x52099, x52100;
  wire x52101, x52102, x52104, x52105, x52106, x52108, x52109, x52110;
  wire x52111, x52113, x52114, x52115, x52117, x52118, x52119, x52120;
  wire x52122, x52123, x52124, x52125, x52126, x52127, x52128, x52130;
  wire x52131, x52132, x52134, x52135, x52136, x52137, x52139, x52140;
  wire x52141, x52143, x52144, x52145, x52146, x52147, x52148, x52149;
  wire x52151, x52152, x52153, x52154, x52155, x52156, x52157, x52159;
  wire x52160, x52161, x52163, x52164, x52165, x52166, x52168, x52169;
  wire x52170, x52172, x52173, x52174, x52175, x52177, x52178, x52179;
  wire x52181, x52182, x52183, x52184, x52186, x52187, x52188, x52189;
  wire x52190, x52191, x52192, x52194, x52195, x52196, x52198, x52199;
  wire x52200, x52201, x52203, x52204, x52205, x52207, x52208, x52209;
  wire x52210, x52212, x52213, x52214, x52216, x52217, x52218, x52219;
  wire x52221, x52222, x52223, x52224, x52225, x52226, x52227, x52229;
  wire x52230, x52231, x52233, x52234, x52235, x52236, x52238, x52239;
  wire x52240, x52242, x52243, x52244, x52245, x52247, x52248, x52249;
  wire x52251, x52252, x52253, x52254, x52255, x52256, x52257, x52259;
  wire x52260, x52261, x52262, x52263, x52264, x52265, x52267, x52268;
  wire x52269, x52271, x52272, x52273, x52274, x52276, x52277, x52278;
  wire x52280, x52281, x52282, x52283, x52285, x52286, x52287, x52289;
  wire x52290, x52291, x52292, x52294, x52295, x52296, x52297, x52298;
  wire x52299, x52300, x52302, x52303, x52304, x52305, x52306, x52307;
  wire x52308, x52310, x52311, x52312, x52314, x52315, x52316, x52317;
  wire x52319, x52320, x52321, x52323, x52324, x52325, x52326, x52328;
  wire x52329, x52330, x52332, x52333, x52334, x52335, x52337, x52338;
  wire x52339, x52341, x52342, x52343, x52344, x52346, x52347, x52348;
  wire x52349, x52350, x52351, x52352, x52354, x52355, x52356, x52358;
  wire x52359, x52360, x52361, x52363, x52364, x52365, x52367, x52368;
  wire x52369, x52370, x52372, x52373, x52374, x52376, x52377, x52378;
  wire x52379, x52381, x52382, x52383, x52385, x52386, x52387, x52388;
  wire x52389, x52390, x52391, x52393, x52394, x52395, x52396, x52397;
  wire x52398, x52399, x52401, x52402, x52403, x52405, x52406, x52407;
  wire x52408, x52410, x52411, x52412, x52414, x52415, x52416, x52417;
  wire x52419, x52420, x52421, x52423, x52424, x52425, x52426, x52428;
  wire x52429, x52430, x52432, x52433, x52434, x52435, x52437, x52438;
  wire x52439, x52441, x52442, x52443, x52444, x52446, x52447, x52448;
  wire x52449, x52450, x52451, x52452, x52454, x52455, x52456, x52458;
  wire x52459, x52460, x52461, x52463, x52464, x52465, x52467, x52468;
  wire x52469, x52470, x52472, x52473, x52474, x52476, x52477, x52478;
  wire x52479, x52481, x52482, x52483, x52485, x52486, x52487, x52488;
  wire x52490, x52491, x52492, x52494, x52495, x52496, x52497, x52499;
  wire x52500, x52501, x52502, x52503, x52504, x52505, x52507, x52508;
  wire x52509, x52511, x52512, x52513, x52514, x52516, x52517, x52518;
  wire x52520, x52521, x52522, x52523, x52525, x52526, x52527, x52529;
  wire x52530, x52531, x52532, x52534, x52535, x52536, x52538, x52539;
  wire x52540, x52541, x52543, x52544, x52545, x52547, x52548, x52549;
  wire x52550, x52551, x52552, x52553, x52555, x52556, x52557, x52558;
  wire x52559, x52560, x52561, x52563, x52564, x52565, x52567, x52568;
  wire x52569, x52570, x52572, x52573, x52574, x52576, x52577, x52578;
  wire x52579, x52581, x52582, x52583, x52585, x52586, x52587, x52588;
  wire x52590, x52591, x52592, x52594, x52595, x52596, x52597, x52599;
  wire x52600, x52601, x52603, x52604, x52605, x52606, x52608, x52609;
  wire x52610, x52612, x52613, x52614, x52615, x52617, x52618, x52619;
  wire x52620, x52621, x52622, x52623, x52625, x52626, x52627, x52629;
  wire x52630, x52631, x52632, x52634, x52635, x52636, x52638, x52639;
  wire x52640, x52641, x52643, x52644, x52645, x52647, x52648, x52649;
  wire x52650, x52652, x52653, x52654, x52656, x52657, x52658, x52659;
  wire x52661, x52662, x52663, x52665, x52666, x52667, x52668, x52670;
  wire x52671, x52672, x52674, x52675, x52676, x52677, x52679, x52680;
  wire x52681, x52682, x52683, x52684, x52685, x52687, x52688, x52689;
  wire x52691, x52692, x52693, x52694, x52696, x52697, x52698, x52700;
  wire x52701, x52702, x52703, x52705, x52706, x52707, x52709, x52710;
  wire x52711, x52712, x52714, x52715, x52716, x52718, x52719, x52720;
  wire x52721, x52723, x52724, x52725, x52727, x52728, x52729, x52730;
  wire x52732, x52733, x52734, x52736, x52737, x52738, x52739, x52740;
  wire x52741, x52742, x52744, x52745, x52746, x52747, x52748, x52749;
  wire x52750, x52752, x52753, x52754, x52756, x52757, x52758, x52759;
  wire x52761, x52762, x52763, x52765, x52766, x52767, x52768, x52770;
  wire x52771, x52772, x52774, x52775, x52776, x52777, x52779, x52780;
  wire x52781, x52783, x52784, x52785, x52786, x52788, x52789, x52790;
  wire x52792, x52793, x52794, x52795, x52797, x52798, x52799, x52801;
  wire x52802, x52803, x52804, x52806, x52807, x52808, x52809, x52810;
  wire x52811, x52812, x52814, x52815, x52816, x52817, x52818, x52819;
  wire x52820, x52822, x52823, x52824, x52826, x52827, x52828, x52829;
  wire x52831, x52832, x52833, x52835, x52836, x52837, x52838, x52840;
  wire x52841, x52842, x52844, x52845, x52846, x52847, x52849, x52850;
  wire x52851, x52853, x52854, x52855, x52856, x52858, x52859, x52860;
  wire x52862, x52863, x52864, x52865, x52867, x52868, x52869, x52871;
  wire x52872, x52873, x52874, x52876, x52877, x52878, x52880, x52881;
  wire x52882, x52883, x52885, x52886, x52887, x52888, x52889, x52890;
  wire x52891, x52893, x52894, x52895, x52897, x52898, x52899, x52900;
  wire x52902, x52903, x52904, x52906, x52907, x52908, x52909, x52911;
  wire x52912, x52913, x52915, x52916, x52917, x52918, x52920, x52921;
  wire x52922, x52924, x52925, x52926, x52927, x52929, x52930, x52931;
  wire x52933, x52934, x52935, x52936, x52938, x52939, x52940, x52942;
  wire x52943, x52944, x52945, x52947, x52948, x52949, x52951, x52952;
  wire x52953, x52954, x52955, x52956, x52957, x52959, x52960, x52961;
  wire x52962, x52963, x52964, x52965, x52967, x52968, x52969, x52971;
  wire x52972, x52973, x52974, x52976, x52977, x52978, x52980, x52981;
  wire x52982, x52983, x52985, x52986, x52987, x52989, x52990, x52991;
  wire x52992, x52994, x52995, x52996, x52998, x52999, x53000, x53001;
  wire x53003, x53004, x53005, x53007, x53008, x53009, x53010, x53012;
  wire x53013, x53014, x53016, x53017, x53018, x53019, x53021, x53022;
  wire x53023, x53025, x53026, x53027, x53028, x53030, x53031, x53032;
  wire x53034, x53035, x53036, x53037, x53039, x53040, x53041, x53042;
  wire x53043, x53044, x53045, x53047, x53048, x53049, x53051, x53052;
  wire x53053, x53054, x53056, x53057, x53058, x53060, x53061, x53062;
  wire x53063, x53065, x53066, x53067, x53069, x53070, x53071, x53072;
  wire x53074, x53075, x53076, x53078, x53079, x53080, x53081, x53083;
  wire x53084, x53085, x53087, x53088, x53089, x53090, x53092, x53093;
  wire x53094, x53096, x53097, x53098, x53099, x53101, x53102, x53103;
  wire x53105, x53106, x53107, x53108, x53110, x53111, x53112, x53114;
  wire x53115, x53116, x53117, x53119, x53120, x53121, x53122, x53123;
  wire x53124, x53125, x53127, x53128, x53129, x53131, x53132, x53133;
  wire x53134, x53136, x53137, x53138, x53140, x53141, x53142, x53143;
  wire x53145, x53146, x53147, x53149, x53150, x53151, x53152, x53154;
  wire x53155, x53156, x53158, x53159, x53160, x53161, x53163, x53164;
  wire x53165, x53167, x53168, x53169, x53170, x53172, x53173, x53174;
  wire x53176, x53177, x53178, x53179, x53181, x53182, x53183, x53185;
  wire x53186, x53187, x53188, x53190, x53191, x53192, x53194, x53195;
  wire x53196, x53197, x53198, x53199, x53200, x53202, x53203, x53204;
  wire x53206, x53207, x53208, x53209, x53211, x53212, x53213, x53215;
  wire x53216, x53217, x53218, x53220, x53221, x53222, x53224, x53225;
  wire x53226, x53227, x53229, x53230, x53231, x53233, x53234, x53235;
  wire x53236, x53238, x53239, x53240, x53242, x53243, x53244, x53245;
  wire x53247, x53248, x53249, x53251, x53252, x53253, x53254, x53256;
  wire x53257, x53258, x53260, x53261, x53262, x53263, x53265, x53266;
  wire x53267, x53269, x53270, x53271, x53272, x53274, x53275, x53276;
  wire x53278, x53279, x53280, x53281, x53283, x53284, x53285, x53287;
  wire x53288, x53289, x53290, x53292, x53293, x53294, x53296, x53297;
  wire x53298, x53299, x53301, x53302, x53303, x53305, x53306, x53307;
  wire x53308, x53310, x53311, x53312, x53314, x53315, x53316, x53317;
  wire x53319, x53320, x53321, x53323, x53324, x53325, x53326, x53328;
  wire x53329, x53330, x53332, x53333, x53334, x53335, x53337, x53338;
  wire x53339, x53341, x53342, x53343, x53344, x53346, x53347, x53348;
  wire x53350, x53351, x53352, x53353, x53355, x53356, x53357, x53359;
  wire x53360, x53361, x53362, x53364, x53365, x53366, x53368, x53369;
  wire x53370, x53371, x53373, x53374, x53375, x53377, x53378, x53379;
  wire x53380, x53382, x53383, x53384, x53386, x53387, x53388, x53390;
  wire x53391, x53392, x53394, x53395, x53396, x53398, x53399, x53400;
  wire x53402, x53403, x53404, x53406, x53407, x53408, x53410, x53411;
  wire x53412, x53414, x53415, x53416, x53418, x53419, x53420, x53422;
  wire x53423, x53424, x53426, x53427, x53428, x53430, x53431, x53432;
  wire x53434, x53435, x53436, x53438, x53439, x53440, x53442, x53443;
  wire x53444, x53446, x53447, x53448, x53450, x53451, x53452, x53454;
  wire x53455, x53456, x53458, x53459, x53460, x53464, x53466, x53467;
  wire x53468, x53471, x53472, x53473, x53474, x53475, x53476, x53479;
  wire x53480, x53481, x53482, x53483, x53484, x53487, x53488, x53490;
  wire x53491, x53492, x53493, x53494, x53495, x53496, x53497, x53500;
  wire x53501, x53503, x53505, x53506, x53507, x53508, x53509, x53510;
  wire x53512, x53513, x53514, x53516, x53517, x53520, x53521, x53523;
  wire x53525, x53526, x53527, x53528, x53529, x53530, x53532, x53533;
  wire x53534, x53536, x53537, x53540, x53541, x53543, x53545, x53546;
  wire x53547, x53548, x53549, x53550, x53552, x53553, x53554, x53556;
  wire x53557, x53560, x53561, x53563, x53565, x53566, x53567, x53569;
  wire x53570, x53571, x53573, x53574, x53575, x53577, x53578, x53581;
  wire x53582, x53584, x53586, x53587, x53588, x53590, x53591, x53592;
  wire x53594, x53595, x53596, x53598, x53599, x53602, x53603, x53605;
  wire x53607, x53608, x53609, x53610, x53612, x53613, x53614, x53615;
  wire x53616, x53618, x53619, x53620, x53622, x53623, x53626, x53627;
  wire x53629, x53631, x53632, x53633, x53634, x53637, x53638, x53639;
  wire x53640, x53641, x53643, x53644, x53645, x53647, x53648, x53649;
  wire x53650, x53651, x53654, x53655, x53657, x53659, x53660, x53661;
  wire x53662, x53665, x53666, x53667, x53668, x53669, x53671, x53672;
  wire x53673, x53675, x53676, x53677, x53678, x53679, x53682, x53683;
  wire x53685, x53687, x53688, x53689, x53690, x53693, x53694, x53696;
  wire x53697, x53698, x53700, x53701, x53702, x53703, x53705, x53706;
  wire x53707, x53709, x53710, x53711, x53712, x53713, x53716, x53717;
  wire x53719, x53721, x53722, x53723, x53724, x53727, x53728, x53730;
  wire x53732, x53733, x53735, x53736, x53737, x53738, x53740, x53741;
  wire x53742, x53744, x53745, x53746, x53747, x53749, x53750, x53751;
  wire x53752, x53753, x53756, x53757, x53759, x53761, x53762, x53763;
  wire x53764, x53767, x53768, x53770, x53772, x53773, x53775, x53776;
  wire x53777, x53778, x53780, x53781, x53782, x53784, x53785, x53786;
  wire x53787, x53789, x53790, x53791, x53792, x53793, x53796, x53797;
  wire x53799, x53801, x53802, x53803, x53804, x53807, x53808, x53810;
  wire x53812, x53813, x53815, x53816, x53817, x53818, x53820, x53821;
  wire x53822, x53824, x53825, x53826, x53827, x53829, x53830, x53831;
  wire x53832, x53833, x53836, x53837, x53839, x53841, x53842, x53843;
  wire x53844, x53847, x53848, x53850, x53852, x53853, x53855, x53857;
  wire x53858, x53859, x53861, x53862, x53863, x53865, x53866, x53867;
  wire x53868, x53870, x53871, x53872, x53874, x53875, x53878, x53879;
  wire x53881, x53883, x53884, x53885, x53886, x53889, x53890, x53892;
  wire x53894, x53895, x53897, x53899, x53900, x53901, x53903, x53904;
  wire x53905, x53907, x53908, x53909, x53910, x53912, x53913, x53914;
  wire x53916, x53917, x53920, x53921, x53923, x53925, x53926, x53927;
  wire x53928, x53931, x53932, x53934, x53936, x53937, x53939, x53940;
  wire x53942, x53943, x53944, x53945, x53946, x53948, x53949, x53950;
  wire x53952, x53953, x53954, x53955, x53957, x53958, x53959, x53961;
  wire x53962, x53965, x53966, x53968, x53970, x53971, x53972, x53973;
  wire x53976, x53977, x53979, x53981, x53982, x53984, x53985, x53988;
  wire x53989, x53990, x53991, x53992, x53994, x53995, x53996, x53998;
  wire x53999, x54000, x54001, x54003, x54004, x54005, x54007, x54008;
  wire x54009, x54010, x54011, x54014, x54015, x54017, x54019, x54020;
  wire x54022, x54023, x54026, x54027, x54029, x54031, x54032, x54034;
  wire x54035, x54038, x54039, x54040, x54041, x54042, x54044, x54045;
  wire x54046, x54048, x54049, x54050, x54051, x54053, x54054, x54055;
  wire x54057, x54058, x54059, x54060, x54061, x54064, x54065, x54067;
  wire x54069, x54070, x54072, x54073, x54076, x54077, x54079, x54081;
  wire x54082, x54084, x54085, x54088, x54089, x54091, x54092, x54093;
  wire x54095, x54096, x54097, x54098, x54100, x54101, x54102, x54104;
  wire x54105, x54106, x54107, x54109, x54110, x54111, x54113, x54114;
  wire x54115, x54116, x54117, x54120, x54121, x54123, x54125, x54126;
  wire x54128, x54129, x54132, x54133, x54135, x54137, x54138, x54140;
  wire x54141, x54144, x54145, x54147, x54149, x54150, x54152, x54153;
  wire x54154, x54155, x54157, x54158, x54159, x54161, x54162, x54163;
  wire x54164, x54166, x54167, x54168, x54170, x54171, x54172, x54173;
  wire x54175, x54176, x54177, x54179, x54180, x54183, x54184, x54186;
  wire x54188, x54189, x54191, x54192, x54195, x54196, x54198, x54200;
  wire x54201, x54203, x54204, x54207, x54208, x54210, x54212, x54213;
  wire x54215, x54216, x54217, x54218, x54220, x54221, x54222, x54224;
  wire x54225, x54226, x54227, x54229, x54230, x54231, x54233, x54234;
  wire x54235, x54236, x54238, x54239, x54240, x54242, x54243, x54246;
  wire x54247, x54249, x54251, x54252, x54254, x54255, x54258, x54259;
  wire x54261, x54263, x54264, x54266, x54267, x54270, x54271, x54273;
  wire x54275, x54276, x54278, x54279, x54280, x54281, x54283, x54284;
  wire x54285, x54287, x54288, x54289, x54291, x54292, x54293, x54294;
  wire x54296, x54297, x54298, x54300, x54301, x54302, x54303, x54305;
  wire x54306, x54307, x54309, x54310, x54313, x54314, x54316, x54318;
  wire x54319, x54321, x54322, x54325, x54326, x54328, x54330, x54331;
  wire x54333, x54334, x54337, x54338, x54340, x54342, x54343, x54345;
  wire x54347, x54348, x54349, x54351, x54352, x54353, x54355, x54356;
  wire x54357, x54359, x54360, x54361, x54362, x54364, x54365, x54366;
  wire x54368, x54369, x54370, x54371, x54373, x54374, x54375, x54377;
  wire x54378, x54381, x54382, x54384, x54386, x54387, x54389, x54392;
  wire x54393, x54395, x54397, x54398, x54400, x54403, x54404, x54406;
  wire x54408, x54409, x54412, x54413, x54414, x54416, x54417, x54418;
  wire x54420, x54421, x54422, x54424, x54425, x54426, x54428, x54429;
  wire x54430, x54432, x54433, x54434, x54436, x54437, x54438, x54440;
  wire x54441, x54442, x54444, x54445, x54446, x54448, x54449, x54450;
  wire x54452, x54453, x54454, x54456, x54457, x54458, x54460, x54461;
  wire x54462, x54465, x54466, x54467, x54471, x54472, x54473, x54477;
  wire x54478, x54479, x54481, x54482, x54483, x54487, x54488, x54489;
  wire x54491, x54492, x54493, x54497, x54498, x54499, x54501, x54502;
  wire x54503, x54507, x54508, x54509, x54511, x54512, x54513, x54515;
  wire x54517, x54518, x54520, x54521, x54522, x54524, x54525, x54526;
  wire x54528, x54530, x54531, x54533, x54534, x54535, x54537, x54538;
  wire x54539, x54541, x54542, x54543, x54545, x54547, x54548, x54550;
  wire x54551, x54552, x54554, x54555, x54556, x54558, x54559, x54560;
  wire x54562, x54565, x54566, x54568, x54569, x54570, x54572, x54573;
  wire x54574, x54576, x54577, x54578, x54580, x54583, x54584, x54586;
  wire x54588, x54589, x54591, x54592, x54593, x54595, x54596, x54597;
  wire x54599, x54602, x54603, x54605, x54607, x54608, x54610, x54611;
  wire x54612, x54614, x54615, x54616, x54618, x54619, x54620, x54622;
  wire x54623, x54626, x54627, x54629, x54631, x54632, x54634, x54635;
  wire x54636, x54638, x54639, x54640, x54642, x54643, x54644, x54646;
  wire x54647, x54648, x54649, x54650, x54653, x54654, x54656, x54658;
  wire x54659, x54661, x54662, x54663, x54665, x54666, x54667, x54669;
  wire x54670, x54671, x54673, x54674, x54675, x54676, x54677, x54680;
  wire x54681, x54683, x54685, x54686, x54688, x54689, x54690, x54692;
  wire x54693, x54694, x54696, x54697, x54698, x54700, x54701, x54702;
  wire x54703, x54704, x54707, x54708, x54710, x54711, x54712, x54714;
  wire x54716, x54718, x54719, x54721, x54722, x54723, x54725, x54726;
  wire x54727, x54729, x54730, x54731, x54733, x54734, x54735, x54736;
  wire x54737, x54740, x54741, x54743, x54744, x54745, x54747, x54749;
  wire x54751, x54752, x54754, x54755, x54756, x54758, x54759, x54760;
  wire x54762, x54763, x54764, x54765, x54767, x54768, x54769, x54771;
  wire x54772, x54773, x54774, x54775, x54778, x54779, x54781, x54782;
  wire x54783, x54785, x54787, x54789, x54790, x54792, x54793, x54794;
  wire x54796, x54797, x54798, x54800, x54801, x54802, x54803, x54805;
  wire x54806, x54807, x54809, x54810, x54811, x54812, x54813, x54816;
  wire x54817, x54819, x54821, x54822, x54824, x54826, x54828, x54829;
  wire x54831, x54832, x54833, x54835, x54836, x54837, x54839, x54840;
  wire x54841, x54842, x54844, x54845, x54846, x54848, x54849, x54850;
  wire x54851, x54852, x54855, x54856, x54858, x54860, x54861, x54863;
  wire x54865, x54867, x54868, x54870, x54872, x54873, x54875, x54876;
  wire x54877, x54879, x54880, x54881, x54882, x54884, x54885, x54886;
  wire x54888, x54889, x54890, x54891, x54892, x54895, x54896, x54898;
  wire x54900, x54901, x54903, x54905, x54907, x54908, x54910, x54912;
  wire x54913, x54915, x54916, x54917, x54919, x54920, x54921, x54922;
  wire x54924, x54925, x54926, x54928, x54929, x54930, x54931, x54932;
  wire x54935, x54936, x54938, x54940, x54941, x54943, x54944, x54946;
  wire x54947, x54949, x54951, x54952, x54954, x54955, x54957, x54958;
  wire x54960, x54961, x54962, x54964, x54965, x54966, x54967, x54969;
  wire x54970, x54971, x54973, x54974, x54975, x54976, x54978, x54979;
  wire x54980, x54982, x54983, x54986, x54987, x54989, x54991, x54992;
  wire x54994, x54996, x54997, x54999, x55001, x55002, x55004, x55006;
  wire x55007, x55009, x55010, x55011, x55013, x55014, x55015, x55017;
  wire x55018, x55019, x55021, x55022, x55023, x55025, x55026, x55027;
  wire x55029, x55030, x55031, x55032, x55033, x55034, x55035, x55036;
  wire x55037, x55039, x55040, x55041, x55043, x55044, x55045, x55046;
  wire x55047, x55048, x55050, x55051, x55052, x55053, x55054, x55055;
  wire x55057, x55058, x55059, x55061, x55062, x55063, x55064, x55065;
  wire x55066, x55067, x55069, x55070, x55071, x55073, x55074, x55075;
  wire x55076, x55077, x55078, x55079, x55081, x55082, x55083, x55085;
  wire x55086, x55087, x55088, x55089, x55090, x55091, x55093, x55094;
  wire x55095, x55097, x55098, x55099, x55100, x55101, x55102, x55103;
  wire x55105, x55106, x55107, x55109, x55110, x55111, x55112, x55114;
  wire x55115, x55116, x55118, x55119, x55120, x55122, x55123, x55124;
  wire x55125, x55127, x55128, x55129, x55131, x55132, x55133, x55135;
  wire x55136, x55137, x55138, x55140, x55141, x55142, x55144, x55145;
  wire x55146, x55148, x55149, x55150, x55151, x55153, x55154, x55155;
  wire x55157, x55158, x55159, x55161, x55162, x55163, x55164, x55166;
  wire x55167, x55168, x55170, x55171, x55172, x55174, x55175, x55176;
  wire x55178, x55179, x55180, x55181, x55183, x55184, x55185, x55187;
  wire x55188, x55189, x55190, x55192, x55193, x55194, x55196, x55197;
  wire x55198, x55200, x55201, x55202, x55203, x55205, x55206, x55207;
  wire x55209, x55210, x55211, x55212, x55214, x55215, x55216, x55218;
  wire x55219, x55220, x55222, x55223, x55224, x55225, x55227, x55228;
  wire x55229, x55231, x55232, x55233, x55234, x55236, x55237, x55238;
  wire x55240, x55241, x55242, x55244, x55245, x55246, x55247, x55249;
  wire x55250, x55251, x55253, x55254, x55255, x55256, x55258, x55259;
  wire x55260, x55262, x55263, x55264, x55266, x55267, x55268, x55269;
  wire x55271, x55272, x55273, x55275, x55277, x55278, x55279, x55281;
  wire x55282, x55283, x55285, x55286, x55287, x55289, x55290, x55291;
  wire x55292, x55294, x55295, x55296, x55298, x55299, x55301, x55302;
  wire x55304, x55305, x55306, x55308, x55309, x55310, x55311, x55313;
  wire x55314, x55315, x55317, x55318, x55319, x55320, x55322, x55323;
  wire x55324, x55326, x55327, x55329, x55330, x55332, x55333, x55334;
  wire x55336, x55337, x55338, x55339, x55341, x55342, x55343, x55345;
  wire x55346, x55347, x55348, x55350, x55351, x55352, x55354, x55355;
  wire x55357, x55358, x55360, x55361, x55362, x55364, x55365, x55366;
  wire x55367, x55369, x55370, x55371, x55373, x55374, x55376, x55377;
  wire x55379, x55380, x55381, x55383, x55384, x55386, x55387, x55389;
  wire x55390, x55391, x55393, x55394, x55395, x55396, x55398, x55399;
  wire x55400, x55402, x55403, x55405, x55406, x55408, x55410, x55411;
  wire x55413, x55414, x55416, x55417, x55419, x55420, x55421, x55423;
  wire x55424, x55425, x55426, x55428, x55429, x55430, x55432, x55433;
  wire x55435, x55436, x55438, x55440, x55441, x55443, x55444, x55446;
  wire x55447, x55449, x55450, x55451, x55453, x55454, x55455, x55456;
  wire x55458, x55459, x55460, x55462, x55463, x55465, x55466, x55468;
  wire x55470, x55471, x55473, x55474, x55476, x55477, x55479, x55480;
  wire x55481, x55483, x55484, x55485, x55486, x55488, x55489, x55490;
  wire x55492, x55493, x55495, x55496, x55498, x55500, x55501, x55503;
  wire x55504, x55506, x55507, x55509, x55510, x55511, x55513, x55514;
  wire x55515, x55516, x55518, x55519, x55520, x55522, x55523, x55525;
  wire x55526, x55528, x55530, x55531, x55533, x55534, x55536, x55537;
  wire x55539, x55540, x55541, x55543, x55544, x55545, x55546, x55548;
  wire x55549, x55550, x55552, x55553, x55556, x55557, x55559, x55561;
  wire x55562, x55564, x55567, x55568, x55570, x55571, x55572, x55574;
  wire x55575, x55576, x55578, x55579, x55580, x55582, x55583, x55584;
  wire x55585, x55586, x55587, x55588, x55589, x55590, x55591, x55592;
  wire x55593, x55595, x55596, x55597, x55598, x55600, x55601, x55603;
  wire x55604, x55605, x55606, x55608, x55609, x55611, x55612, x55613;
  wire x55614, x55616, x55617, x55619, x55620, x55621, x55622, x55624;
  wire x55625, x55627, x55628, x55629, x55630, x55632, x55633, x55635;
  wire x55636, x55637, x55639, x55640, x55641, x55643, x55644, x55646;
  wire x55647, x55649, x55650, x55651, x55653, x55654, x55655, x55657;
  wire x55658, x55660, x55661, x55663, x55664, x55665, x55667, x55668;
  wire x55669, x55671, x55672, x55674, x55675, x55677, x55678, x55679;
  wire x55681, x55682, x55683, x55685, x55686, x55688, x55689, x55691;
  wire x55692, x55693, x55695, x55696, x55697, x55699, x55700, x55701;
  wire x55702, x55704, x55706, x55707, x55709, x55710, x55711, x55712;
  wire x55714, x55715, x55716, x55718, x55719, x55721, x55722, x55724;
  wire x55726, x55727, x55729, x55730, x55731, x55732, x55734, x55735;
  wire x55736, x55738, x55739, x55741, x55742, x55744, x55746, x55747;
  wire x55749, x55750, x55751, x55752, x55754, x55755, x55756, x55758;
  wire x55759, x55761, x55762, x55764, x55766, x55767, x55769, x55770;
  wire x55771, x55772, x55774, x55775, x55776, x55778, x55779, x55781;
  wire x55782, x55784, x55786, x55787, x55789, x55790, x55791, x55792;
  wire x55794, x55795, x55796, x55798, x55799, x55801, x55802, x55804;
  wire x55806, x55807, x55809, x55810, x55811, x55812, x55814, x55815;
  wire x55816, x55818, x55819, x55822, x55823, x55825, x55827, x55828;
  wire x55830, x55831, x55832, x55833, x55835, x55836, x55837, x55839;
  wire x55840, x55843, x55844, x55846, x55848, x55849, x55851, x55852;
  wire x55853, x55854, x55856, x55857, x55858, x55860, x55861, x55864;
  wire x55865, x55867, x55869, x55870, x55872, x55873, x55874, x55875;
  wire x55877, x55878, x55879, x55881, x55882, x55885, x55886, x55888;
  wire x55890, x55891, x55893, x55894, x55895, x55896, x55898, x55899;
  wire x55900, x55902, x55903, x55906, x55907, x55909, x55911, x55912;
  wire x55914, x55915, x55916, x55917, x55919, x55920, x55921, x55923;
  wire x55924, x55927, x55928, x55930, x55932, x55933, x55935, x55936;
  wire x55937, x55938, x55940, x55941, x55942, x55944, x55945, x55948;
  wire x55949, x55951, x55953, x55954, x55956, x55957, x55958, x55959;
  wire x55961, x55962, x55963, x55965, x55966, x55969, x55970, x55972;
  wire x55974, x55975, x55977, x55978, x55979, x55980, x55982, x55983;
  wire x55984, x55986, x55987, x55990, x55991, x55993, x55995, x55996;
  wire x55998, x55999, x56000, x56002, x56003, x56004, x56006, x56007;
  wire x56008, x56009, x56010, x56011, x56013, x56014, x56015, x56017;
  wire x56018, x56019, x56021, x56022, x56023, x56025, x56026, x56027;
  wire x56028, x56030, x56031, x56032, x56034, x56035, x56036, x56037;
  wire x56039, x56040, x56041, x56043, x56044, x56045, x56046, x56048;
  wire x56049, x56050, x56052, x56053, x56054, x56055, x56057, x56058;
  wire x56059, x56061, x56062, x56063, x56064, x56067, x56069, x56070;
  wire x56072, x56073, x56074, x56076, x56077, x56078, x56079, x56082;
  wire x56084, x56085, x56087, x56088, x56089, x56091, x56092, x56093;
  wire x56094, x56097, x56099, x56100, x56102, x56103, x56104, x56106;
  wire x56107, x56108, x56109, x56112, x56114, x56115, x56117, x56118;
  wire x56119, x56121, x56122, x56123, x56124, x56127, x56129, x56130;
  wire x56132, x56133, x56134, x56136, x56137, x56138, x56139, x56142;
  wire x56145, x56146, x56148, x56149, x56150, x56152, x56153, x56154;
  wire x56155, x56158, x56161, x56162, x56164, x56165, x56166, x56168;
  wire x56169, x56170, x56171, x56174, x56177, x56178, x56180, x56181;
  wire x56182, x56184, x56185, x56186, x56187, x56190, x56193, x56194;
  wire x56196, x56197, x56198, x56200, x56201, x56202, x56203, x56206;
  wire x56209, x56210, x56212, x56213, x56214, x56216, x56217, x56218;
  wire x56219, x56222, x56225, x56226, x56228, x56229, x56230, x56232;
  wire x56233, x56234, x56235, x56238, x56241, x56242, x56244, x56245;
  wire x56246, x56248, x56249, x56250, x56251, x56254, x56257, x56258;
  wire x56260, x56261, x56262, x56264, x56265, x56266, x56267, x56270;
  wire x56273, x56274, x56276, x56277, x56278, x56280, x56281, x56282;
  wire x56283, x56286, x56289, x56290, x56292, x56293, x56294, x56296;
  wire x56297, x56298, x56299, x56302, x56305, x56306, x56308, x56309;
  wire x56310, x56312, x56313, x56314, x56315, x56318, x56321, x56322;
  wire x56324, x56325, x56326, x56328, x56329, x56330, x56331, x56334;
  wire x56337, x56338, x56340, x56341, x56342, x56344, x56345, x56346;
  wire x56347, x56350, x56353, x56354, x56356, x56357, x56358, x56360;
  wire x56361, x56362, x56364, x56365, x56366, x56367, x56368, x56369;
  wire x56370, x56371, x56372, x56374, x56375, x56376, x56379, x56380;
  wire x56381, x56384, x56385, x56386, x56389, x56390, x56391, x56394;
  wire x56395, x56396, x56398, x56400, x56401, x56403, x56404, x56405;
  wire x56407, x56408, x56410, x56411, x56413, x56414, x56415, x56417;
  wire x56418, x56420, x56421, x56423, x56424, x56425, x56427, x56428;
  wire x56430, x56431, x56433, x56434, x56435, x56437, x56438, x56440;
  wire x56441, x56443, x56444, x56445, x56447, x56448, x56450, x56451;
  wire x56453, x56454, x56455, x56457, x56458, x56460, x56461, x56463;
  wire x56464, x56465, x56467, x56468, x56470, x56471, x56473, x56474;
  wire x56475, x56477, x56478, x56480, x56481, x56483, x56484, x56485;
  wire x56487, x56488, x56490, x56491, x56493, x56494, x56495, x56497;
  wire x56498, x56500, x56501, x56503, x56504, x56505, x56507, x56508;
  wire x56510, x56511, x56513, x56514, x56515, x56517, x56518, x56520;
  wire x56521, x56523, x56524, x56525, x56527, x56528, x56530, x56531;
  wire x56533, x56534, x56535, x56537, x56538, x56540, x56541, x56543;
  wire x56544, x56545, x56547, x56548, x56550, x56551, x56553, x56554;
  wire x56555, x56557, x56558, x56560, x56561, x56563, x56564, x56565;
  wire x56567, x56568, x56570, x56571, x56573, x56574, x56575, x56577;
  wire x56578, x56580, x56581, x56583, x56584, x56585, x56587, x56588;
  wire x56589, x56591, x56592, x56593, x56594, x56595, x56596, x56597;
  wire x56599, x56600, x56601, x56603, x56604, x56605, x56607, x56608;
  wire x56609, x56611, x56612, x56613, x56614, x56616, x56617, x56618;
  wire x56620, x56621, x56622, x56623, x56625, x56626, x56627, x56629;
  wire x56630, x56631, x56632, x56634, x56635, x56636, x56638, x56639;
  wire x56640, x56641, x56643, x56644, x56645, x56647, x56648, x56649;
  wire x56650, x56652, x56653, x56654, x56656, x56657, x56658, x56659;
  wire x56661, x56662, x56663, x56665, x56666, x56668, x56669, x56671;
  wire x56672, x56673, x56675, x56676, x56678, x56679, x56681, x56682;
  wire x56683, x56685, x56686, x56688, x56689, x56691, x56692, x56693;
  wire x56695, x56696, x56698, x56699, x56701, x56702, x56703, x56705;
  wire x56706, x56708, x56709, x56711, x56712, x56713, x56715, x56716;
  wire x56718, x56719, x56721, x56722, x56723, x56725, x56726, x56728;
  wire x56729, x56731, x56732, x56733, x56735, x56736, x56738, x56739;
  wire x56741, x56742, x56743, x56745, x56746, x56748, x56749, x56751;
  wire x56752, x56753, x56755, x56756, x56758, x56759, x56761, x56762;
  wire x56763, x56765, x56766, x56768, x56769, x56771, x56772, x56773;
  wire x56775, x56776, x56778, x56779, x56781, x56782, x56783, x56785;
  wire x56786, x56788, x56789, x56791, x56792, x56793, x56795, x56796;
  wire x56798, x56799, x56801, x56802, x56803, x56805, x56806, x56808;
  wire x56809, x56811, x56812, x56813, x56815, x56816, x56818, x56819;
  wire x56821, x56822, x56823, x56825, x56826, x56828, x56829, x56831;
  wire x56832, x56833, x56835, x56836, x56838, x56839, x56841, x56842;
  wire x56843, x56845, x56847, x56848, x56849, x56850, x56851, x56853;
  wire x56854, x56855, x56857, x56859, x56860, x56862, x56864, x56865;
  wire x56867, x56869, x56870, x56872, x56874, x56875, x56877, x56879;
  wire x56880, x56882, x56884, x56885, x56887, x56889, x56890, x56892;
  wire x56894, x56895, x56897, x56899, x56900, x56902, x56904, x56905;
  wire x56907, x56909, x56910, x56912, x56914, x56915, x56917, x56919;
  wire x56920, x56922, x56924, x56925, x56927, x56929, x56930, x56932;
  wire x56934, x56935, x56937, x56939, x56940, x56942, x56944, x56945;
  wire x56947, x56949, x56950, x56952, x56954, x56955, x56957, x56959;
  wire x56960, x56962, x56964, x56965, x56967, x56969, x56970, x56972;
  wire x56974, x56975, x57002, x57003, x57004, x57005, x57006, x57008;
  wire x57009, x57010, x57012, x57013, x57014, x57016, x57017, x57018;
  wire x57020, x57021, x57022, x57024, x57025, x57026, x57028, x57029;
  wire x57030, x57032, x57033, x57034, x57036, x57037, x57038, x57040;
  wire x57041, x57042, x57044, x57045, x57046, x57048, x57049, x57050;
  wire x57052, x57053, x57054, x57056, x57057, x57058, x57060, x57061;
  wire x57062, x57064, x57065, x57066, x57068, x57069, x57070, x57072;
  wire x57073, x57074, x57076, x57077, x57078, x57080, x57081, x57082;
  wire x57084, x57085, x57086, x57088, x57089, x57090, x57092, x57093;
  wire x57094, x57096, x57097, x57098, x57101, x57103, x57104, x57106;
  wire x57107, x57109, x57110, x57112, x57114, x57115, x57117, x57119;
  wire x57120, x57122, x57124, x57125, x57127, x57129, x57130, x57132;
  wire x57134, x57135, x57137, x57139, x57140, x57142, x57144, x57145;
  wire x57147, x57149, x57150, x57152, x57154, x57155, x57157, x57159;
  wire x57160, x57162, x57164, x57165, x57167, x57169, x57170, x57172;
  wire x57174, x57175, x57177, x57179, x57180, x57182, x57184, x57185;
  wire x57187, x57189, x57190, x57192, x57194, x57195, x57197, x57199;
  wire x57200, x57202, x57204, x57205, x57207, x57209, x57210, x57212;
  wire x57214, x57215, x57219, x57221, x57222, x57224, x57225, x57227;
  wire x57228, x57230, x57231, x57233, x57234, x57236, x57238, x57239;
  wire x57241, x57243, x57244, x57246, x57248, x57249, x57251, x57253;
  wire x57254, x57256, x57258, x57259, x57261, x57263, x57264, x57266;
  wire x57268, x57269, x57271, x57273, x57274, x57276, x57278, x57279;
  wire x57281, x57283, x57284, x57286, x57288, x57289, x57291, x57293;
  wire x57294, x57296, x57298, x57299, x57301, x57303, x57304, x57306;
  wire x57308, x57309, x57311, x57313, x57314, x57316, x57318, x57319;
  wire x57325, x57327, x57328, x57330, x57331, x57333, x57334, x57336;
  wire x57337, x57339, x57340, x57342, x57343, x57345, x57346, x57348;
  wire x57349, x57351, x57352, x57354, x57356, x57357, x57359, x57361;
  wire x57362, x57364, x57366, x57367, x57369, x57371, x57372, x57374;
  wire x57376, x57377, x57379, x57381, x57382, x57384, x57386, x57387;
  wire x57389, x57391, x57392, x57394, x57396, x57397, x57405, x57407;
  wire x57408, x57410, x57411, x57413, x57414, x57416, x57417, x57419;
  wire x57420, x57422, x57423, x57425, x57426, x57428, x57429, x57431;
  wire x57432, x57434, x57435, x57436, x57438, x57439, x57440, x57442;
  wire x57443, x57444, x57446, x57447, x57448, x57450, x57451, x57452;
  wire x57454, x57455, x57456, x57458, x57459, x57460, x57462, x57463;
  wire x57464, x57466, x57468, x57469, x57471, x57473, x57474, x57476;
  wire x57477, x57478, x57480, x57481, x57482, x57484, x57485, x57486;
  wire x57488, x57489, x57490, x57492, x57493, x57494, x57496, x57497;
  wire x57498, x57500, x57502, x57503, x57505, x57507, x57508, x57510;
  wire x57512, x57513, x57515, x57517, x57518, x57520, x57522, x57523;
  wire x57525, x57527, x57528, x57530, x57532, x57533, x57535, x57537;
  wire x57538, x57540, x57542, x57543, x57545, x57547, x57548, x57550;
  wire x57552, x57554, x57556, x57558, x57560, x57562, x57564, x57566;
  wire x57568, x57570, x57572, x57574, x57576, x57578, x57580, x57582;
  wire x57584, x57586, x57588, x57590, x57592, x57594, x57596, x57598;
  wire x57600, x57602, x57604, x57606, x57608, x57610, x57611, x57613;
  wire x57615, x57617, x57619, x57621, x57623, x57625, x57627, x57629;
  wire x57631, x57633, x57635, x57637, x57639, x57641, x57643, x57645;
  wire x57647, x57649, x57651, x57653, x57655, x57657, x57659, x57661;
  wire x57663, x57665, x57667, x57668, x57669, x57670, x57672, x57674;
  wire x57676, x57678, x57680, x57682, x57684, x57686, x57688, x57690;
  wire x57692, x57694, x57696, x57698, x57700, x57702, x57704, x57706;
  wire x57708, x57710, x57712, x57714, x57716, x57718, x57719, x57720;
  wire x57721, x57722, x57723, x57724, x57725, x57726, x57728, x57730;
  wire x57732, x57734, x57736, x57738, x57740, x57742, x57744, x57746;
  wire x57748, x57750, x57752, x57754, x57756, x57757, x57758, x57759;
  wire x57760, x57761, x57762, x57763, x57764, x57765, x57766, x57767;
  wire x57768, x57769, x57770, x57771, x57772, x57774, x57775, x57776;
  wire x57778, x57779, x57780, x57782, x57783, x57784, x57786, x57787;
  wire x57788, x57790, x57791, x57792, x57794, x57795, x57796, x57798;
  wire x57799, x57800, x57802, x57803, x57804, x57806, x57807, x57808;
  wire x57810, x57811, x57812, x57814, x57815, x57816, x57818, x57819;
  wire x57820, x57822, x57823, x57824, x57826, x57827, x57828, x57830;
  wire x57831, x57832, x57834, x57835, x57836, x57838, x57839, x57840;
  wire x57842, x57843, x57844, x57846, x57847, x57848, x57850, x57851;
  wire x57852, x57854, x57855, x57856, x57858, x57859, x57860, x57862;
  wire x57863, x57864, x57866, x57867, x57868, x57870, x57871, x57872;
  wire x57874, x57875, x57876, x57878, x57879, x57880, x57882, x57883;
  wire x57884, x57886, x57887, x57888, x57890, x57891, x57892, x57895;
  wire x57897, x57899, x57901, x57903, x57905, x57907, x57909, x57911;
  wire x57913, x57915, x57917, x57919, x57921, x57923, x57925, x57927;
  wire x57928, x57929, x57930, x57931, x57932, x57933, x57934, x57935;
  wire x57936, x57937, x57938, x57939, x57940, x57941, x57942, x57943;
  wire x57944, x57945, x57946, x57947, x57948, x57949, x57950, x57951;
  wire x57952, x57953, x57954, x57955, x57956, x57957, x57958, x57959;
  wire x57961, x57963, x57965, x57967, x57969, x57971, x57973, x57975;
  wire x57977, x57979, x57981, x57983, x57985, x57987, x57989, x57991;
  wire x57993, x57995, x57997, x57999, x58001, x58003, x58005, x58007;
  wire x58009, x58011, x58013, x58015, x58017, x58019, x58021, x58023;
  wire x58024, x58025, x58026, x58027, x58028, x58029, x58030, x58031;
  wire x58032, x58033, x58034, x58035, x58036, x58037, x58038, x58039;
  wire x58040, x58041, x58042, x58043, x58044, x58045, x58046, x58047;
  wire x58048, x58049, x58050, x58051, x58052, x58053, x58054, x58055;
  wire x58056, x58057, x58058, x58059, x58060, x58061, x58062, x58063;
  wire x58064, x58065, x58066, x58067, x58068, x58069, x58070, x58071;
  wire x58072, x58073, x58074, x58075, x58076, x58077, x58078, x58079;
  wire x58080, x58081, x58082, x58083, x58084, x58085, x58086, x58087;
  wire x58088, x58089, x58090, x58091, x58092, x58093, x58094, x58095;
  wire x58096, x58097, x58098, x58099, x58100, x58101, x58102, x58103;
  wire x58104, x58105, x58106, x58107, x58108, x58109, x58110, x58111;
  wire x58112, x58113, x58114, x58115, x58116, x58117, x58118, x58119;
  wire x58120, x58121, x58122, x58123, x58124, x58125, x58126, x58127;
  wire x58128, x58129, x58130, x58131, x58132, x58133, x58134, x58135;
  wire x58136, x58137, x58138, x58139, x58140, x58141, x58142, x58143;
  wire x58144, x58145, x58146, x58147, x58148, x58149, x58150, x58151;
  wire x58152, x58153, x58154, x58155, x58156, x58157, x58158, x58159;
  wire x58160, x58161, x58162, x58163, x58164, x58165, x58166, x58167;
  wire x58168, x58169, x58170, x58171, x58172, x58173, x58174, x58175;
  wire x58176, x58177, x58178, x58179, x58180, x58181, x58182, x58183;
  wire x58184, x58185, x58186, x58187, x58188, x58189, x58190, x58191;
  wire x58192, x58193, x58194, x58195, x58196, x58197, x58198, x58199;
  wire x58200, x58201, x58202, x58203, x58204, x58205, x58206, x58207;
  wire x58208, x58209, x58210, x58211, x58212, x58213, x58214, x58215;
  wire x58216, x58217, x58218, x58219, x58220, x58221, x58222, x58223;
  wire x58224, x58225, x58226, x58227, x58228, x58229, x58230, x58231;
  wire x58232, x58233, x58234, x58235, x58236, x58237, x58238, x58239;
  wire x58240, x58241, x58242, x58243, x58244, x58245, x58246, x58247;
  wire x58248, x58249, x58250, x58251, x58252, x58253, x58254, x58255;
  wire x58256, x58257, x58258, x58259, x58260, x58261, x58262, x58263;
  wire x58264, x58265, x58266, x58267, x58268, x58269, x58270, x58271;
  wire x58272, x58273, x58274, x58275, x58276, x58277, x58278, x58279;
  wire x58280, x58281, x58282, x58283, x58284, x58285, x58286, x58287;
  wire x58288, x58289, x58290, x58291, x58292, x58293, x58294, x58295;
  wire x58296, x58297, x58298, x58299, x58300, x58301, x58302, x58303;
  wire x58304, x58305, x58306, x58307, x58308, x58309, x58310, x58311;
  wire x58312, x58313, x58314, x58315, x58316, x58317, x58318, x58319;
  wire x58320, x58321, x58322, x58323, x58324, x58325, x58326, x58327;
  wire x58328, x58329, x58330, x58331, x58332, x58333, x58334, x58335;
  wire x58336, x58337, x58338, x58339, x58340, x58341, x58342, x58343;
  wire x58344, x58345, x58346, x58347, x58348, x58349, x58350, x58351;
  wire x58352, x58353, x58354, x58355, x58356, x58357, x58358, x58359;
  wire x58360, x58361, x58362, x58363, x58364, x58365, x58366, x58367;
  wire x58368, x58369, x58370, x58371, x58372, x58373, x58374, x58375;
  wire x58376, x58377, x58378, x58379, x58380, x58381, x58382, x58383;
  wire x58384, x58385, x58386, x58387, x58388, x58389, x58390, x58391;
  wire x58392, x58393, x58394, x58395, x58396, x58397, x58398, x58399;
  wire x58400, x58401, x58402, x58403, x58404, x58405, x58406, x58407;
  wire x58408, x58409, x58410, x58411, x58412, x58413, x58414, x58415;
  wire x58416, x58417, x58418, x58419, x58420, x58421, x58422, x58423;
  wire x58424, x58425, x58426, x58427, x58428, x58429, x58430, x58431;
  wire x58432, x58433, x58434, x58435, x58436, x58437, x58438, x58439;
  wire x58440, x58441, x58442, x58443, x58444, x58445, x58446, x58447;
  wire x58448, x58449, x58450, x58451, x58452, x58453, x58454, x58455;
  wire x58456, x58457, x58458, x58459, x58460, x58461, x58462, x58463;
  wire x58464, x58465, x58466, x58467, x58468, x58469, x58470, x58471;
  wire x58472, x58473, x58474, x58475, x58476, x58477, x58478, x58479;
  wire x58480, x58481, x58482, x58483, x58484, x58485, x58486, x58487;
  wire x58488, x58489, x58490, x58491, x58492, x58493, x58494, x58495;
  wire x58496, x58497, x58498, x58499, x58500, x58501, x58502, x58503;
  wire x58504, x58505, x58506, x58507, x58508, x58509, x58510, x58511;
  wire x58512, x58513, x58514, x58515, x58516, x58517, x58518, x58519;
  wire x58520, x58521, x58522, x58523, x58524, x58525, x58526, x58527;
  wire x58528, x58529, x58530, x58531, x58532, x58533, x58534, x58535;
  wire x58536, x58537, x58538, x58539, x58540, x58541, x58542, x58543;
  wire x58544, x58545, x58546, x58547, x58548, x58549, x58550, x58551;
  wire x58552, x58553, x58554, x58555, x58556, x58557, x58558, x58559;
  wire x58560, x58561, x58562, x58563, x58564, x58565, x58566, x58567;
  wire x58568, x58569, x58570, x58571, x58572, x58573, x58574, x58575;
  wire x58576, x58577, x58578, x58579, x58580, x58581, x58582, x58583;
  wire x58584, x58585, x58586, x58587, x58588, x58589, x58590, x58591;
  wire x58592, x58593, x58594, x58595, x58596, x58597, x58598, x58599;
  wire x58600, x58601, x58602, x58603, x58604, x58605, x58606, x58607;
  wire x58608, x58609, x58610, x58611, x58612, x58613, x58614, x58615;
  wire x58616, x58617, x58618, x58619, x58620, x58621, x58622, x58623;
  wire x58624, x58625, x58626, x58627, x58628, x58629, x58630, x58631;
  wire x58632, x58633, x58634, x58635, x58636, x58637, x58638, x58639;
  wire x58640, x58641, x58642, x58643, x58644, x58645, x58646, x58647;
  wire x58648, x58649, x58650, x58651, x58652, x58653, x58654, x58655;
  wire x58656, x58657, x58658, x58659, x58660, x58661, x58662, x58663;
  wire x58664, x58665, x58666, x58667, x58668, x58669, x58670, x58671;
  wire x58672, x58673, x58674, x58675, x58676, x58677, x58678, x58679;
  wire x58680, x58681, x58682, x58683, x58684, x58685, x58686, x58687;
  wire x58688, x58689, x58690, x58691, x58692, x58693, x58694, x58695;
  wire x58696, x58697, x58698, x58699, x58700, x58701, x58702, x58703;
  wire x58704, x58705, x58706, x58707, x58708, x58709, x58710, x58711;
  wire x58712, x58713, x58714, x58715, x58716, x58717, x58718, x58719;
  wire x58720, x58721, x58722, x58723, x58724, x58725, x58726, x58727;
  wire x58728, x58729, x58730, x58731, x58732, x58733, x58734, x58735;
  wire x58736, x58737, x58738, x58739, x58740, x58741, x58742, x58743;
  wire x58744, x58745, x58746, x58747, x58748, x58749, x58750, x58751;
  wire x58752, x58753, x58754, x58755, x58756, x58757, x58758, x58759;
  wire x58760, x58761, x58762, x58763, x58764, x58765, x58766, x58767;
  wire x58768, x58769, x58770, x58771, x58772, x58773, x58774, x58775;
  wire x58776, x58777, x58778, x58779, x58780, x58781, x58782, x58783;
  wire x58784, x58785, x58786, x58787, x58788, x58789, x58790, x58791;
  wire x58792, x58793, x58794, x58795, x58796, x58797, x58798, x58799;
  wire x58800, x58801, x58802, x58803, x58804, x58805, x58806, x58807;
  wire x58808, x58809, x58810, x58811, x58812, x58813, x58814, x58815;
  wire x58816, x58817, x58818, x58819, x58820, x58821, x58822, x58823;
  wire x58824, x58825, x58826, x58827, x58828, x58829, x58830, x58831;
  wire x58832, x58833, x58834, x58835, x58836, x58837, x58838, x58839;
  wire x58840, x58841, x58842, x58843, x58844, x58845, x58846, x58847;
  wire x58848, x58849, x58850, x58851, x58852, x58853, x58854, x58855;
  wire x58856, x58857, x58858, x58859, x58860, x58861, x58862, x58863;
  wire x58864, x58865, x58866, x58867, x58868, x58869, x58870, x58871;
  wire x58872, x58873, x58874, x58875, x58876, x58877, x58878, x58879;
  wire x58880, x58881, x58882, x58883, x58884, x58885, x58886, x58887;
  wire x58888, x58889, x58890, x58891, x58892, x58893, x58894, x58895;
  wire x58896, x58897, x58898, x58899, x58900, x58901, x58902, x58903;
  wire x58904, x58905, x58906, x58907, x58908, x58909, x58910, x58911;
  wire x58912, x58913, x58914, x58915, x58916, x58917, x58918, x58919;
  wire x58920, x58921, x58922, x58923, x58924, x58925, x58926, x58927;
  wire x58928, x58929, x58930, x58931, x58932, x58933, x58934, x58935;
  wire x58936, x58937, x58938, x58939, x58940, x58941, x58942, x58943;
  wire x58944, x58945, x58946, x58947, x58948, x58949, x58950, x58951;
  wire x58952, x58953, x58954, x58955, x58956, x58957, x58958, x58959;
  wire x58960, x58961, x58962, x58963, x58964, x58965, x58966, x58967;
  wire x58968, x58969, x58970, x58971, x58972, x58973, x58974, x58975;
  wire x58976, x58977, x58978, x58979, x58980, x58981, x58982, x58983;
  wire x58984, x58985, x58986, x58987, x58988, x58989, x58990, x58991;
  wire x58992, x58993, x58994, x58995, x58996, x58997, x58998, x58999;
  wire x59000, x59001, x59002, x59003, x59004, x59005, x59006, x59007;
  wire x59008, x59009, x59010, x59011, x59012, x59013, x59014, x59015;
  wire x59016, x59017, x59018, x59019, x59020, x59021, x59022, x59023;
  wire x59024, x59025, x59026, x59027, x59028, x59029, x59030, x59031;
  wire x59032, x59033, x59034, x59035, x59036, x59037, x59038, x59039;
  wire x59040, x59041, x59042, x59043, x59044, x59045, x59046, x59047;
  wire x59048, x59049, x59050, x59051, x59052, x59053, x59054, x59055;
  wire x59056, x59057, x59058, x59059, x59060, x59061, x59062, x59063;
  wire x59064, x59065, x59066, x59067, x59068, x59069, x59070, x59071;
  wire x59072, x59073, x59074, x59075, x59076, x59077, x59078, x59079;
  wire x59080, x59081, x59082, x59083, x59084, x59085, x59086, x59087;
  wire x59088, x59089, x59090, x59091, x59092, x59093, x59094, x59095;
  wire x59096, x59097, x59098, x59099, x59100, x59101, x59102, x59103;
  wire x59104, x59105, x59106, x59107, x59108, x59109, x59110, x59111;
  wire x59112, x59113, x59114, x59115, x59116, x59117, x59118, x59119;
  wire x59120, x59121, x59122, x59123, x59124, x59125, x59126, x59127;
  wire x59128, x59129, x59130, x59131, x59132, x59133, x59134, x59135;
  wire x59136, x59137, x59138, x59139, x59140, x59141, x59142, x59143;
  wire x59144, x59145, x59146, x59147, x59148, x59149, x59150, x59151;
  wire x59152, x59153, x59154, x59155, x59156, x59157, x59158, x59159;
  wire x59160, x59161, x59162, x59163, x59164, x59165, x59166, x59167;
  wire x59168, x59169, x59170, x59171, x59172, x59173, x59174, x59175;
  wire x59176, x59177, x59178, x59179, x59180, x59181, x59182, x59183;
  wire x59184, x59185, x59186, x59187, x59188, x59189, x59190, x59191;
  wire x59192, x59193, x59194, x59195, x59196, x59197, x59198, x59199;
  wire x59200, x59201, x59202, x59203, x59204, x59205, x59206, x59207;
  wire x59208, x59209, x59210, x59211, x59212, x59213, x59214, x59215;
  wire x59216, x59217, x59218, x59219, x59220, x59221, x59222, x59223;
  wire x59224, x59225, x59226, x59227, x59228, x59229, x59230, x59231;
  wire x59232, x59233, x59234, x59235, x59236, x59237, x59238, x59239;
  wire x59240, x59241, x59242, x59243, x59244, x59245, x59246, x59247;
  wire x59248, x59249, x59250, x59251, x59252, x59253, x59254, x59255;
  wire x59256, x59257, x59258, x59259, x59260, x59261, x59262, x59263;
  wire x59264, x59265, x59266, x59267, x59268, x59269, x59270, x59271;
  wire x59272, x59273, x59274, x59275, x59276, x59277, x59278, x59279;
  wire x59280, x59281, x59282, x59283, x59284, x59285, x59286, x59287;
  wire x59288, x59289, x59290, x59291, x59292, x59293, x59294, x59295;
  wire x59296, x59297, x59298, x59299, x59300, x59301, x59302, x59303;
  wire x59304, x59305, x59306, x59307, x59308, x59309, x59310, x59311;
  wire x59312, x59313, x59314, x59315, x59316, x59317, x59318, x59319;
  wire x59320, x59321, x59322, x59323, x59324, x59325, x59326, x59327;
  wire x59328, x59329, x59330, x59331, x59332, x59333, x59334, x59335;
  wire x59336, x59337, x59338, x59339, x59340, x59341, x59342, x59343;
  wire x59344, x59345, x59346, x59347, x59348, x59349, x59350, x59351;
  wire x59352, x59353, x59354, x59355, x59356, x59357, x59358, x59359;
  wire x59360, x59361, x59362, x59363, x59364, x59365, x59366, x59367;
  wire x59368, x59369, x59370, x59371, x59372, x59373, x59374, x59375;
  wire x59376, x59377, x59378, x59379, x59380, x59381, x59382, x59383;
  wire x59384, x59385, x59386, x59387, x59388, x59389, x59390, x59391;
  wire x59392, x59393, x59394, x59395, x59396, x59397, x59398, x59399;
  wire x59400, x59401, x59402, x59403, x59404, x59405, x59406, x59407;
  wire x59408, x59409, x59410, x59411, x59412, x59413, x59414, x59415;
  wire x59416, x59417, x59418, x59419, x59420, x59421, x59422, x59423;
  wire x59424, x59425, x59426, x59427, x59428, x59429, x59430, x59431;
  wire x59432, x59433, x59434, x59435, x59436, x59437, x59438, x59439;
  wire x59440, x59441, x59442, x59443, x59444, x59445, x59446, x59447;
  wire x59448, x59449, x59450, x59451, x59452, x59453, x59454, x59455;
  wire x59456, x59457, x59458, x59459, x59460, x59461, x59462, x59463;
  wire x59464, x59465, x59466, x59467, x59468, x59469, x59470, x59471;
  wire x59472, x59473, x59474, x59475, x59476, x59477, x59478, x59479;
  wire x59480, x59481, x59482, x59483, x59484, x59485, x59486, x59487;
  wire x59488, x59489, x59490, x59491, x59492, x59493, x59494, x59495;
  wire x59496, x59497, x59498, x59499, x59500, x59501, x59502, x59503;
  wire x59504, x59505, x59506, x59507, x59508, x59509, x59510, x59511;
  wire x59512, x59513, x59514, x59515, x59516, x59517, x59518, x59519;
  wire x59520, x59521, x59522, x59523, x59524, x59525, x59526, x59527;
  wire x59528, x59529, x59530, x59531, x59532, x59533, x59534, x59535;
  wire x59536, x59537, x59538, x59539, x59540, x59541, x59542, x59543;
  wire x59544, x59545, x59546, x59547, x59548, x59549, x59550, x59551;
  wire x59552, x59553, x59554, x59555, x59556, x59557, x59558, x59559;
  wire x59560, x59561, x59562, x59563, x59564, x59565, x59566, x59567;
  wire x59568, x59569, x59570, x59571, x59572, x59573, x59574, x59575;
  wire x59576, x59577, x59578, x59579, x59580, x59581, x59582, x59583;
  wire x59584, x59585, x59586, x59587, x59588, x59589, x59590, x59591;
  wire x59592, x59593, x59594, x59595, x59596, x59597, x59598, x59599;
  wire x59600, x59601, x59602, x59603, x59604, x59605, x59606, x59607;
  wire x59608, x59609, x59610, x59611, x59612, x59613, x59614, x59615;
  wire x59616, x59617, x59618, x59619, x59620, x59621, x59622, x59623;
  wire x59624, x59625, x59626, x59627, x59628, x59629, x59630, x59631;
  wire x59632, x59633, x59634, x59635, x59636, x59637, x59638, x59639;
  wire x59640, x59641, x59642, x59643, x59644, x59645, x59646, x59647;
  wire x59648, x59649, x59650, x59651, x59652, x59653, x59654, x59655;
  wire x59656, x59657, x59658, x59659, x59660, x59661, x59662, x59663;
  wire x59664, x59665, x59666, x59667, x59668, x59669, x59670, x59671;
  wire x59672, x59673, x59674, x59675, x59676, x59677, x59678, x59679;
  wire x59680, x59681, x59682, x59683, x59684, x59685, x59686, x59687;
  wire x59688, x59689, x59690, x59691, x59692, x59693, x59694, x59695;
  wire x59696, x59697, x59698, x59699, x59700, x59701, x59702, x59703;
  wire x59704, x59705, x59706, x59707, x59708, x59709, x59710, x59711;
  wire x59712, x59713, x59714, x59715, x59716, x59717, x59718, x59719;
  wire x59720, x59721, x59722, x59723, x59724, x59725, x59726, x59727;
  wire x59728, x59729, x59730, x59731, x59732, x59733, x59734, x59735;
  wire x59736, x59737, x59738, x59739, x59740, x59741, x59742, x59743;
  wire x59744, x59745, x59746, x59747, x59748, x59749, x59750, x59751;
  wire x59752, x59753, x59754, x59755, x59756, x59757, x59758, x59759;
  wire x59760, x59761, x59762, x59763, x59764, x59765, x59766, x59767;
  wire x59768, x59769, x59770, x59771, x59772, x59773, x59774, x59775;
  wire x59776, x59777, x59778, x59779, x59780, x59781, x59782, x59783;
  wire x59784, x59785, x59786, x59787, x59788, x59789, x59790, x59791;
  wire x59792, x59793, x59794, x59795, x59796, x59797, x59798, x59799;
  wire x59800, x59801, x59802, x59803, x59804, x59805, x59806, x59807;
  wire x59808, x59809, x59810, x59811, x59812, x59813, x59814, x59815;
  wire x59816, x59817, x59818, x59819, x59820, x59821, x59822, x59823;
  wire x59824, x59825, x59826, x59827, x59828, x59829, x59830, x59831;
  wire x59832, x59833, x59834, x59835, x59836, x59837, x59838, x59839;
  wire x59840, x59841, x59842, x59843, x59844, x59845, x59846, x59847;
  wire x59848, x59849, x59850, x59851, x59852, x59853, x59854, x59855;
  wire x59856, x59857, x59858, x59859, x59860, x59861, x59862, x59863;
  wire x59864, x59865, x59866, x59867, x59868, x59869, x59870, x59871;
  wire x59872, x59873, x59874, x59875, x59876, x59877, x59878, x59879;
  wire x59880, x59881, x59882, x59883, x59884, x59885, x59886, x59887;
  wire x59888, x59889, x59890, x59891, x59892, x59893, x59894, x59895;
  wire x59896, x59897, x59898, x59899, x59900, x59901, x59902, x59903;
  wire x59904, x59905, x59906, x59907, x59908, x59909, x59910, x59911;
  wire x59912, x59913, x59914, x59915, x59916, x59917, x59918, x59919;
  wire x59920, x59921, x59922, x59923, x59924, x59925, x59926, x59927;
  wire x59928, x59929, x59930, x59931, x59932, x59933, x59934, x59935;
  wire x59936, x59937, x59938, x59939, x59940, x59941, x59942, x59943;
  wire x59944, x59945, x59946, x59947, x59948, x59949, x59950, x59951;
  wire x59952, x59953, x59954, x59955, x59956, x59957, x59958, x59959;
  wire x59960, x59961, x59962, x59963, x59964, x59965, x59966, x59967;
  wire x59968, x59969, x59970, x59971, x59972, x59973, x59974, x59975;
  wire x59976, x59977, x59978, x59979, x59980, x59981, x59982, x59983;
  wire x59984, x59985, x59986, x59987, x59988, x59989, x59990, x59991;
  wire x59992, x59993, x59994, x59995, x59996, x59997, x59998, x59999;
  wire x60000, x60001, x60002, x60003, x60004, x60005, x60006, x60007;
  wire x60008, x60009, x60010, x60011, x60012, x60013, x60014, x60015;
  wire x60016, x60017, x60018, x60019, x60020, x60021, x60022, x60023;
  wire x60024, x60025, x60026, x60027, x60028, x60029, x60030, x60031;
  wire x60032, x60033, x60034, x60035, x60036, x60037, x60038, x60039;
  wire x60040, x60041, x60042, x60043, x60044, x60045, x60046, x60047;
  wire x60048, x60049, x60050, x60051, x60052, x60053, x60054, x60055;
  wire x60056, x60057, x60058, x60059, x60060, x60061, x60062, x60063;
  wire x60064, x60065, x60066, x60067, x60068, x60069, x60070, x60071;
  wire x60072, x60073, x60074, x60075, x60076, x60077, x60078, x60079;
  wire x60080, x60081, x60082, x60083, x60084, x60085, x60086, x60087;
  wire x60088, x60089, x60090, x60091, x60092, x60093, x60094, x60095;
  wire x60096, x60097, x60098, x60099, x60100, x60101, x60102, x60103;
  wire x60104, x60105, x60106, x60107, x60108, x60109, x60110, x60111;
  wire x60112, x60113, x60114, x60115, x60116, x60117, x60118, x60119;
  wire x60120, x60121, x60122, x60123, x60124, x60125, x60126, x60127;
  wire x60128, x60129, x60130, x60131, x60132, x60133, x60134, x60135;
  wire x60136, x60137, x60138, x60139, x60140, x60141, x60142, x60143;
  wire x60144, x60145, x60146, x60147, x60148, x60149, x60150, x60151;
  wire x60152, x60153, x60154, x60155, x60156, x60157, x60158, x60159;
  wire x60160, x60161, x60162, x60163, x60164, x60165, x60166, x60167;
  wire x60168, x60169, x60170, x60171, x60172, x60173, x60174, x60175;
  wire x60176, x60177, x60178, x60179, x60180, x60181, x60182, x60183;
  wire x60184, x60185, x60186, x60187, x60188, x60189, x60190, x60191;
  wire x60192, x60193, x60194, x60195, x60196, x60197, x60198, x60199;
  wire x60200, x60201, x60202, x60203, x60204, x60205, x60206, x60207;
  wire x60208, x60209, x60210, x60211, x60212, x60213, x60214, x60215;
  wire x60216, x60217, x60218, x60219, x60220, x60221, x60222, x60223;
  wire x60224, x60225, x60226, x60227, x60228, x60229, x60230, x60231;
  wire x60232, x60233, x60234, x60235, x60236, x60237, x60238, x60239;
  wire x60240, x60241, x60242, x60243, x60244, x60245, x60246, x60247;
  wire x60248, x60249, x60250, x60251, x60252, x60253, x60254, x60255;
  wire x60256, x60257, x60258, x60259, x60260, x60261, x60262, x60263;
  wire x60264, x60265, x60266, x60267, x60268, x60269, x60270, x60271;
  wire x60272, x60273, x60274, x60275, x60276, x60277, x60278, x60279;
  wire x60280, x60281, x60282, x60283, x60284, x60285, x60286, x60287;
  wire x60288, x60289, x60290, x60291, x60292, x60293, x60294, x60295;
  wire x60296, x60297, x60298, x60299, x60300, x60301, x60302, x60303;
  wire x60304, x60305, x60306, x60307, x60308, x60309, x60310, x60311;
  wire x60312, x60313, x60314, x60315, x60316, x60317, x60318, x60319;
  wire x60320, x60321, x60322, x60323, x60324, x60325, x60326, x60327;
  wire x60328, x60329, x60330, x60331, x60332, x60333, x60334, x60335;
  wire x60336, x60337, x60338, x60339, x60340, x60341, x60342, x60343;
  wire x60344, x60345, x60346, x60347, x60348, x60349, x60350, x60351;
  wire x60352, x60353, x60354, x60355, x60356, x60357, x60358, x60359;
  wire x60360, x60361, x60362, x60363, x60364, x60365, x60366, x60367;
  wire x60368, x60369, x60370, x60371, x60372, x60373, x60374, x60375;
  wire x60376, x60377, x60378, x60379, x60380, x60381, x60382, x60383;
  wire x60384, x60385, x60386, x60387, x60388, x60389, x60390, x60391;
  wire x60392, x60393, x60394, x60395, x60396, x60397, x60398, x60399;
  wire x60400, x60401, x60402, x60403, x60404, x60405, x60406, x60407;
  wire x60408, x60409, x60410, x60411, x60412, x60413, x60414, x60415;
  wire x60416, x60417, x60418, x60419, x60420, x60421, x60422, x60423;
  wire x60424, x60425, x60426, x60427, x60428, x60429, x60430, x60431;
  wire x60432, x60433, x60434, x60435, x60436, x60437, x60438, x60439;
  wire x60440, x60441, x60442, x60443, x60444, x60445, x60446, x60447;
  wire x60448, x60449, x60450, x60451, x60452, x60453, x60454, x60455;
  wire x60456, x60457, x60458, x60459, x60460, x60461, x60462, x60463;
  wire x60464, x60465, x60466, x60467, x60468, x60469, x60470, x60471;
  wire x60472, x60473, x60474, x60475, x60476, x60477, x60478, x60479;
  wire x60480, x60481, x60482, x60483, x60484, x60485, x60486, x60487;
  wire x60488, x60489, x60490, x60491, x60492, x60493, x60494, x60495;
  wire x60496, x60497, x60498, x60499, x60500, x60501, x60502, x60503;
  wire x60504, x60505, x60506, x60507, x60508, x60509, x60510, x60511;
  wire x60512, x60513, x60514, x60515, x60516, x60517, x60518, x60519;
  wire x60520, x60521, x60522, x60523, x60524, x60525, x60526, x60527;
  wire x60528, x60529, x60530, x60531, x60532, x60533, x60534, x60535;
  wire x60536, x60537, x60538, x60539, x60540, x60541, x60542, x60543;
  wire x60544, x60545, x60546, x60547, x60548, x60549, x60550, x60551;
  wire x60552, x60553, x60554, x60555, x60556, x60557, x60558, x60559;
  wire x60560, x60561, x60562, x60563, x60564, x60565, x60566, x60567;
  wire x60568, x60569, x60570, x60571, x60572, x60573, x60574, x60575;
  wire x60576, x60577, x60578, x60579, x60580, x60581, x60582, x60583;
  wire x60584, x60585, x60586, x60587, x60588, x60589, x60590, x60591;
  wire x60592, x60593, x60594, x60595, x60596, x60597, x60598, x60599;
  wire x60600, x60601, x60602, x60603, x60604, x60605, x60606, x60607;
  wire x60608, x60609, x60610, x60611, x60612, x60613, x60614, x60615;
  wire x60616, x60617, x60618, x60619, x60620, x60621, x60622, x60623;
  wire x60624, x60625, x60626, x60627, x60628, x60629, x60630, x60631;
  wire x60632, x60633, x60634, x60635, x60636, x60637, x60638, x60639;
  wire x60640, x60641, x60642, x60643, x60644, x60645, x60646, x60647;
  wire x60648, x60649, x60650, x60651, x60652, x60653, x60654, x60655;
  wire x60657, x60658, x60659, x60661, x60662, x60663, x60665, x60666;
  wire x60667, x60669, x60670, x60671, x60673, x60674, x60675, x60677;
  wire x60678, x60679, x60681, x60682, x60683, x60685, x60686, x60687;
  wire x60689, x60690, x60691, x60693, x60694, x60695, x60697, x60698;
  wire x60699, x60701, x60702, x60703, x60705, x60706, x60707, x60709;
  wire x60710, x60711, x60713, x60714, x60715, x60717, x60718, x60719;
  wire x60721, x60722, x60723, x60725, x60726, x60727, x60729, x60730;
  wire x60731, x60733, x60734, x60735, x60737, x60738, x60739, x60741;
  wire x60742, x60743, x60745, x60746, x60747, x60749, x60750, x60751;
  wire x60753, x60754, x60755, x60757, x60758, x60759, x60761, x60762;
  wire x60763, x60765, x60766, x60767, x60769, x60770, x60771, x60773;
  wire x60774, x60775, x60777, x60778, x60779, x60781, x60782, x60783;
  wire x60785, x60786, x60787, x60789, x60790, x60791, x60793, x60794;
  wire x60795, x60797, x60798, x60799, x60801, x60802, x60803, x60805;
  wire x60806, x60807, x60809, x60810, x60811, x60813, x60814, x60815;
  wire x60817, x60818, x60819, x60821, x60822, x60823, x60825, x60826;
  wire x60827, x60829, x60830, x60831, x60833, x60834, x60835, x60837;
  wire x60838, x60839, x60841, x60845, x60848, x60851, x60854, x60857;
  wire x60860, x60863, x60866, x60869, x60872, x60875, x60878, x60881;
  wire x60884, x60887, x60890, x60893, x60896, x60899, x60902, x60905;
  wire x60908, x60911, x60914, x60917, x60920, x60923, x60926, x60929;
  wire x60932, x60935, x60936, x60940, x60941, x60945, x60946, x60947;
  wire x60948, x60949, x60950, x60951, x60952, x60953, x60954, x60956;
  wire x60957, x60958, x60959, x60960, x60961, x60963, x60964, x60965;
  wire x60966, x60968, x60969, x60971, x60972, x60973, x60974, x60975;
  wire x60979, x60982, x60985, x60988, x60991, x60994, x60997, x61000;
  wire x61003, x61006, x61009, x61012, x61015, x61018, x61021, x61024;
  wire x61027, x61030, x61033, x61036, x61039, x61042, x61045, x61048;
  wire x61051, x61054, x61057, x61060, x61063, x61066, x61069, x61070;
  wire x61074, x61075, x61078, x61079, x61080, x61081, x61082, x61083;
  wire x61084, x61085, x61086, x61087, x61088, x61089, x61090, x61091;
  wire x61092, x61093, x61094, x61095, x61096, x61097, x61098, x61099;
  wire x61100, x61101, x61102, x61103, x61104, x61108, x61111, x61114;
  wire x61117, x61120, x61123, x61126, x61129, x61132, x61135, x61138;
  wire x61141, x61144, x61147, x61150, x61153, x61156, x61159, x61162;
  wire x61165, x61168, x61171, x61174, x61177, x61180, x61183, x61186;
  wire x61189, x61192, x61195, x61198, x61199, x61203, x61204, x61207;
  wire x61208, x61209, x61210, x61211, x61212, x61213, x61214, x61215;
  wire x61216, x61217, x61218, x61219, x61220, x61221, x61222, x61223;
  wire x61224, x61225, x61226, x61227, x61228, x61229, x61230, x61231;
  wire x61232, x61233, x61237, x61240, x61243, x61246, x61249, x61252;
  wire x61255, x61258, x61261, x61264, x61267, x61270, x61273, x61276;
  wire x61279, x61282, x61285, x61288, x61291, x61294, x61297, x61300;
  wire x61303, x61306, x61309, x61312, x61315, x61318, x61321, x61324;
  wire x61327, x61328, x61332, x61333, x61336, x61337, x61338, x61339;
  wire x61340, x61341, x61342, x61343, x61344, x61345, x61346, x61347;
  wire x61348, x61349, x61350, x61351, x61352, x61353, x61354, x61355;
  wire x61356, x61357, x61358, x61359, x61360, x61361, x61362, x61364;
  wire x61365, x61366, x61368, x61369, x61370, x61372, x61373, x61374;
  wire x61376, x61377, x61378, x61380, x61381, x61382, x61384, x61385;
  wire x61386, x61388, x61389, x61390, x61392, x61393, x61394, x61396;
  wire x61397, x61398, x61400, x61401, x61402, x61404, x61405, x61406;
  wire x61408, x61409, x61410, x61412, x61413, x61414, x61416, x61417;
  wire x61418, x61420, x61421, x61422, x61424, x61426, x61685, x61687;
  wire x61688, x61689, x61690, x61691, x61692, x61693, x61694, x61695;
  wire x61696, x61697, x61698, x61699, x61700, x61701, x61702, x61703;
  wire x61704, x61705, x61706, x61707, x61708, x61709, x61710, x61711;
  wire x61712, x61713, x61714, x61715, x61716, x61717, x61718, x61719;
  wire x61720, x61721, x61722, x61723, x61724, x61725, x61726, x61727;
  wire x61728, x61729, x61730, x61731, x61732, x61733, x61734, x61735;
  wire x61736, x61737, x61738, x61739, x61740, x61741, x61742, x61743;
  wire x61744, x61745, x61746, x61747, x61748, x61749, x61750, x61751;
  wire x61752, x61753, x61754, x61755, x61756, x61757, x61758, x61759;
  wire x61760, x61761, x61762, x61763, x61764, x61765, x61766, x61767;
  wire x61768, x61769, x61770, x61771, x61772, x61773, x61774, x61775;
  wire x61776, x61777, x61778, x61779, x61780, x61781, x61782, x61783;
  wire x61784, x61785, x61786, x61787, x61788, x61789, x61790, x61791;
  wire x61792, x61793, x61794, x61795, x61796, x61797, x61798, x61799;
  wire x61800, x61801, x61802, x61803, x61804, x61805, x61806, x61807;
  wire x61808, x61809, x61810, x61811, x61812, x61813, x61814, x61815;
  wire x61816, x61817, x61818, x61819, x61820, x61821, x61822, x61823;
  wire x61824, x61825, x61826, x61827, x61828, x61829, x61830, x61831;
  wire x61832, x61833, x61834, x61835, x61836, x61837, x61838, x61839;
  wire x61840, x61841, x61842, x61843, x61844, x61845, x61846, x61847;
  wire x61848, x61849, x61850, x61851, x61852, x61853, x61854, x61855;
  wire x61856, x61857, x61858, x61859, x61860, x61861, x61862, x61863;
  wire x61864, x61865, x61866, x61867, x61868, x61869, x61870, x61871;
  wire x61872, x61873, x61874, x61875, x61876, x61877, x61878, x61879;
  wire x61880, x61881, x61882, x61883, x61884, x61885, x61886, x61887;
  wire x61888, x61889, x61890, x61891, x61892, x61893, x61894, x61895;
  wire x61896, x61897, x61898, x61899, x61900, x61901, x61902, x61903;
  wire x61904, x61905, x61906, x61907, x61908, x61909, x61910, x61911;
  wire x61912, x61913, x61914, x61915, x61916, x61917, x61918, x61919;
  wire x61920, x61921, x61922, x61923, x61924, x61925, x61926, x61927;
  wire x61928, x61929, x61930, x61931, x61932, x61933, x61934, x61935;
  wire x61936, x61937, x61938, x61939, x61940, x61941, x61942, x61943;
  wire x61944, x61945, x61946, x61947, x61948, x61949, x61950, x61951;
  wire x61952, x61953, x61954, x61955, x61956, x61957, x61958, x61959;
  wire x61960, x61961, x61962, x61963, x61964, x61965, x61966, x61967;
  wire x61968, x61969, x61970, x61971, x61972, x61973, x61974, x61976;
  wire x61977, x61978, x61979, x61980, x61982, x61983, x61984, x61985;
  wire x61986, x61987, x61989, x61990, x61991, x61992, x61993, x61994;
  wire x61996, x61997, x61998, x61999, x62000, x62001, x62003, x62004;
  wire x62005, x62006, x62007, x62008, x62010, x62011, x62012, x62013;
  wire x62014, x62015, x62017, x62018, x62019, x62020, x62021, x62022;
  wire x62024, x62025, x62026, x62027, x62028, x62029, x62031, x62032;
  wire x62033, x62034, x62035, x62036, x62038, x62039, x62040, x62041;
  wire x62042, x62043, x62045, x62046, x62047, x62048, x62049, x62050;
  wire x62052, x62053, x62054, x62055, x62056, x62057, x62059, x62060;
  wire x62061, x62062, x62063, x62064, x62066, x62067, x62068, x62069;
  wire x62070, x62071, x62073, x62074, x62075, x62076, x62077, x62078;
  wire x62080, x62081, x62082, x62083, x62084, x62085, x62087, x62088;
  wire x62089, x62090, x62091, x62092, x62094, x62095, x62096, x62097;
  wire x62098, x62099, x62101, x62102, x62103, x62104, x62105, x62106;
  wire x62108, x62109, x62110, x62111, x62112, x62113, x62115, x62116;
  wire x62117, x62118, x62119, x62120, x62122, x62123, x62124, x62125;
  wire x62126, x62127, x62129, x62130, x62131, x62132, x62133, x62134;
  wire x62136, x62137, x62138, x62139, x62140, x62141, x62143, x62144;
  wire x62145, x62146, x62147, x62148, x62150, x62151, x62152, x62153;
  wire x62154, x62155, x62157, x62158, x62159, x62160, x62161, x62162;
  wire x62164, x62165, x62166, x62167, x62168, x62169, x62171, x62172;
  wire x62173, x62174, x62175, x62176, x62178, x62179, x62180, x62181;
  wire x62182, x62183, x62185, x62186, x62187, x62188, x62189, x62190;
  wire x62192, x62193, x62194, x62195, x62196, x62197, x62199, x62200;
  wire x62201, x62202, x62203, x62204, x62206, x62207, x62208, x62209;
  wire x62210, x62211, x62213, x62214, x62215, x62216, x62217, x62218;
  wire x62220, x62221, x62222, x62223, x62224, x62225, x62227, x62228;
  wire x62229, x62230, x62231, x62232, x62234, x62235, x62236, x62237;
  wire x62238, x62239, x62241, x62242, x62243, x62244, x62245, x62246;
  wire x62248, x62249, x62250, x62251, x62252, x62253, x62255, x62256;
  wire x62257, x62258, x62259, x62260, x62262, x62263, x62264, x62265;
  wire x62266, x62267, x62269, x62270, x62271, x62272, x62273, x62274;
  wire x62276, x62277, x62278, x62279, x62280, x62281, x62283, x62284;
  wire x62285, x62286, x62287, x62288, x62290, x62291, x62292, x62293;
  wire x62294, x62295, x62297, x62298, x62299, x62300, x62301, x62302;
  wire x62304, x62305, x62306, x62307, x62308, x62309, x62311, x62312;
  wire x62313, x62314, x62315, x62316, x62318, x62319, x62320, x62321;
  wire x62322, x62323, x62325, x62326, x62327, x62328, x62329, x62330;
  wire x62332, x62333, x62334, x62335, x62336, x62337, x62339, x62340;
  wire x62341, x62342, x62343, x62344, x62346, x62347, x62348, x62349;
  wire x62350, x62351, x62353, x62354, x62355, x62356, x62357, x62358;
  wire x62360, x62361, x62362, x62363, x62364, x62365, x62367, x62368;
  wire x62369, x62370, x62371, x62372, x62374, x62375, x62376, x62377;
  wire x62378, x62379, x62381, x62382, x62383, x62384, x62385, x62386;
  wire x62388, x62389, x62390, x62391, x62392, x62393, x62395, x62396;
  wire x62397, x62398, x62399, x62400, x62402, x62403, x62404, x62405;
  wire x62406, x62407, x62409, x62410, x62411, x62412, x62413, x62414;
  wire x62416, x62417, x62418, x62419, x62420, x62421, x62423, x62424;
  wire x62425, x62426, x62427, x62428, x62430, x62431, x62432, x62433;
  wire x62434, x62435, x62437, x62438, x62439, x62440, x62441, x62442;
  wire x62444, x62445, x62446, x62447, x62448, x62449, x62451, x62452;
  wire x62453, x62454, x62455, x62456, x62458, x62459, x62460, x62461;
  wire x62462, x62463, x62465, x62466, x62467, x62468, x62469, x62470;
  wire x62472, x62473, x62474, x62475, x62476, x62477, x62479, x62480;
  wire x62481, x62482, x62483, x62484, x62486, x62487, x62488, x62489;
  wire x62490, x62491, x62493, x62494, x62495, x62496, x62497, x62498;
  wire x62500, x62501, x62502, x62503, x62504, x62505, x62507, x62508;
  wire x62509, x62510, x62511, x62512, x62514, x62515, x62516, x62517;
  wire x62518, x62519, x62521, x62522, x62523, x62524, x62525, x62526;
  wire x62528, x62529, x62530, x62531, x62532, x62533, x62535, x62536;
  wire x62537, x62538, x62539, x62540, x62542, x62543, x62544, x62545;
  wire x62546, x62547, x62549, x62550, x62551, x62552, x62553, x62554;
  wire x62556, x62557, x62558, x62559, x62560, x62561, x62563, x62564;
  wire x62565, x62566, x62567, x62568, x62570, x62571, x62572, x62573;
  wire x62574, x62575, x62577, x62578, x62579, x62580, x62581, x62582;
  wire x62584, x62585, x62586, x62587, x62588, x62589, x62591, x62592;
  wire x62593, x62594, x62595, x62596, x62598, x62599, x62600, x62601;
  wire x62602, x62603, x62605, x62606, x62607, x62608, x62609, x62610;
  wire x62612, x62613, x62614, x62615, x62616, x62617, x62619, x62620;
  wire x62621, x62622, x62623, x62624, x62626, x62627, x62628, x62629;
  wire x62630, x62631, x62633, x62634, x62635, x62636, x62637, x62638;
  wire x62640, x62641, x62642, x62643, x62644, x62645, x62647, x62648;
  wire x62649, x62650, x62651, x62652, x62654, x62655, x62656, x62657;
  wire x62658, x62659, x62661, x62662, x62663, x62664, x62665, x62666;
  wire x62668, x62669, x62670, x62671, x62672, x62673, x62675, x62676;
  wire x62677, x62678, x62679, x62680, x62682, x62683, x62684, x62685;
  wire x62686, x62687, x62689, x62690, x62691, x62692, x62693, x62694;
  wire x62696, x62697, x62698, x62699, x62700, x62701, x62703, x62704;
  wire x62705, x62706, x62707, x62708, x62710, x62711, x62712, x62713;
  wire x62714, x62715, x62717, x62718, x62719, x62720, x62721, x62722;
  wire x62724, x62725, x62726, x62727, x62728, x62729, x62731, x62732;
  wire x62733, x62734, x62735, x62736, x62738, x62739, x62740, x62741;
  wire x62742, x62743, x62745, x62746, x62747, x62748, x62749, x62750;
  wire x62752, x62753, x62754, x62755, x62756, x62757, x62759, x62760;
  wire x62761, x62762, x62763, x62764, x62766, x62767, x62768, x62769;
  wire x62770, x62771, x62773, x62774, x62775, x62776, x62777, x62778;
  wire x62780, x62781, x62782, x62783, x62784, x62785, x62787, x62788;
  wire x62789, x62790, x62791, x62792, x62794, x62795, x62796, x62797;
  wire x62798, x62799, x62801, x62802, x62803, x62804, x62805, x62806;
  wire x62808, x62809, x62810, x62811, x62812, x62813, x62815, x62816;
  wire x62817, x62818, x62819, x62820, x62822, x62823, x62824, x62825;
  wire x62826, x62827, x62829, x62830, x62831, x62832, x62833, x62834;
  wire x62836, x62837, x62838, x62839, x62840, x62841, x62843, x62844;
  wire x62845, x62846, x62847, x62848, x62850, x62851, x62852, x62853;
  wire x62854, x62855, x62857, x62858, x62859, x62860, x62861, x62862;
  wire x62864, x62865, x62866, x62867, x62868, x62869, x62871, x62872;
  wire x62874, x62875, x62876, x62878, x62879, x62880, x62882, x62883;
  wire x62884, x62886, x62887, x62888, x62890, x62891, x62892, x62894;
  wire x62895, x62896, x62898, x62899, x62900, x62902, x62903, x62904;
  wire x62906, x62907, x62908, x62910, x62911, x62912, x62914, x62915;
  wire x62916, x62918, x62919, x62920, x62922, x62923, x62924, x62926;
  wire x62927, x62928, x62930, x62932, x62934, x62935, x62936, x62937;
  wire x62938, x62939, x62940, x62941, x62942, x62943, x62944, x62945;
  wire x62946, x62947, x62948, x62949, x62950, x62951, x62952, x62953;
  wire x62954, x62955, x62956, x62957, x62958, x62959, x62960, x62961;
  wire x62962, x62963, x62964, x62965, x62966, x62967, x62968, x62969;
  wire x62970, x62971, x62972, x62973, x62974, x62975, x62976, x62977;
  wire x62978, x62979, x62980, x62981, x62982, x62983, x62984, x62985;
  wire x62986, x62987, x62988, x62989, x62990, x62991, x62992, x62993;
  wire x62994, x62995, x62996, x62997, x62998, x62999, x63000, x63001;
  wire x63002, x63003, x63004, x63005, x63006, x63007, x63008, x63009;
  wire x63010, x63011, x63012, x63013, x63014, x63015, x63016, x63017;
  wire x63018, x63019, x63020, x63021, x63022, x63023, x63024, x63025;
  wire x63026, x63029, x63030, x63031, x63034, x63035, x63037, x63040;
  wire x63041, x63043, x63046, x63047, x63049, x63052, x63053, x63055;
  wire x63058, x63059, x63061, x63064, x63065, x63067, x63070, x63071;
  wire x63073, x63076, x63077, x63079, x63082, x63083, x63085, x63088;
  wire x63089, x63091, x63094, x63095, x63097, x63100, x63101, x63103;
  wire x63106, x63107, x63109, x63112, x63113, x63115, x63118, x63119;
  wire x63121, x63124, x63125, x63127, x63130, x63131, x63133, x63136;
  wire x63137, x63139, x63142, x63143, x63145, x63148, x63149, x63151;
  wire x63154, x63155, x63157, x63160, x63161, x63163, x63166, x63167;
  wire x63169, x63172, x63173, x63175, x63178, x63179, x63181, x63184;
  wire x63185, x63187, x63190, x63191, x63193, x63196, x63197, x63199;
  wire x63202, x63203, x63205, x63208, x63209, x63240, x63241, x63242;
  wire x63243, x63244, x63246, x63247, x63248, x63250, x63251, x63252;
  wire x63254, x63255, x63256, x63258, x63259, x63260, x63262, x63263;
  wire x63264, x63266, x63267, x63268, x63270, x63271, x63272, x63274;
  wire x63275, x63276, x63278, x63279, x63280, x63282, x63283, x63284;
  wire x63286, x63287, x63288, x63290, x63291, x63292, x63294, x63295;
  wire x63296, x63298, x63299, x63300, x63302, x63303, x63304, x63306;
  wire x63307, x63308, x63310, x63311, x63312, x63314, x63315, x63316;
  wire x63318, x63319, x63320, x63322, x63323, x63324, x63326, x63327;
  wire x63328, x63330, x63331, x63332, x63334, x63335, x63336, x63338;
  wire x63339, x63340, x63342, x63343, x63344, x63346, x63347, x63348;
  wire x63350, x63351, x63352, x63355, x63357, x63358, x63360, x63361;
  wire x63363, x63364, x63366, x63368, x63369, x63371, x63373, x63374;
  wire x63376, x63378, x63379, x63381, x63383, x63384, x63386, x63388;
  wire x63389, x63391, x63393, x63394, x63396, x63398, x63399, x63401;
  wire x63403, x63404, x63406, x63408, x63409, x63411, x63413, x63414;
  wire x63416, x63418, x63419, x63421, x63423, x63424, x63426, x63428;
  wire x63429, x63431, x63433, x63434, x63436, x63438, x63439, x63441;
  wire x63443, x63444, x63446, x63448, x63449, x63451, x63453, x63454;
  wire x63456, x63458, x63459, x63461, x63463, x63464, x63466, x63468;
  wire x63469, x63471, x63473, x63474, x63476, x63478, x63479, x63481;
  wire x63483, x63484, x63486, x63488, x63489, x63492, x63494, x63495;
  wire x63497, x63498, x63500, x63501, x63503, x63504, x63506, x63507;
  wire x63509, x63511, x63512, x63514, x63516, x63517, x63519, x63521;
  wire x63522, x63524, x63526, x63527, x63529, x63531, x63532, x63534;
  wire x63536, x63537, x63539, x63541, x63542, x63544, x63546, x63547;
  wire x63549, x63551, x63552, x63554, x63556, x63557, x63559, x63561;
  wire x63562, x63564, x63566, x63567, x63569, x63571, x63572, x63574;
  wire x63576, x63577, x63579, x63581, x63582, x63584, x63586, x63587;
  wire x63589, x63591, x63592, x63594, x63596, x63597, x63599, x63601;
  wire x63602, x63604, x63606, x63607, x63609, x63611, x63612, x63615;
  wire x63617, x63618, x63620, x63621, x63623, x63624, x63626, x63627;
  wire x63629, x63630, x63632, x63633, x63635, x63636, x63638, x63639;
  wire x63641, x63642, x63644, x63646, x63647, x63649, x63651, x63652;
  wire x63654, x63656, x63657, x63659, x63661, x63662, x63664, x63666;
  wire x63667, x63669, x63671, x63672, x63674, x63676, x63677, x63679;
  wire x63681, x63682, x63684, x63686, x63687, x63689, x63691, x63692;
  wire x63694, x63696, x63697, x63699, x63701, x63702, x63704, x63706;
  wire x63707, x63710, x63712, x63713, x63715, x63716, x63718, x63719;
  wire x63721, x63722, x63724, x63725, x63727, x63728, x63730, x63731;
  wire x63733, x63734, x63736, x63737, x63739, x63740, x63742, x63743;
  wire x63745, x63746, x63748, x63749, x63751, x63752, x63753, x63754;
  wire x63755, x63756, x63758, x63760, x63761, x63763, x63764, x63765;
  wire x63767, x63769, x63770, x63772, x63774, x63775, x63777, x63779;
  wire x63780, x63782, x63783, x63784, x63786, x63788, x63789, x63791;
  wire x63793, x63794, x63795, x63797, x63798, x63799, x63801, x63802;
  wire x63803, x63805, x63806, x63807, x63809, x63810, x63811, x63813;
  wire x63814, x63815, x63816, x63817, x63818, x63820, x63821, x63822;
  wire x63824, x63825, x63826, x63828, x63829, x63830, x63832, x63833;
  wire x63834, x63836, x63837, x63838, x63840, x63841, x63842, x63844;
  wire x63845, x63846, x63848, x63849, x63850, x63852, x63853, x63854;
  wire x63856, x63857, x63858, x63860, x63861, x63862, x63864, x63865;
  wire x63866, x63868, x63869, x63870, x63872, x63873, x63874, x63913;
  wire x63915, x63916, x63917, x63918, x63919, x63920, x63921, x63922;
  wire x63923, x63924, x63925, x63926, x63927, x63928, x63929, x63930;
  wire x63931, x63932, x63933, x63934, x63935, x63936, x63937, x63938;
  wire x63939, x63940, x63941, x63942, x63943, x63944, x63945, x63946;
  wire x63947, x63948, x63949, x63950, x63951, x63952, x63953, x63954;
  wire x63955, x63956, x63957, x63958, x63959, x63960, x63961, x63962;
  wire x63963, x63964, x63965, x63966, x63967, x63968, x63969, x63970;
  wire x63971, x63972, x63973, x63974, x63975, x63976, x63977, x63978;
  wire x63979, x63980, x63981, x63982, x63983, x63984, x63985, x63986;
  wire x63987, x63988, x63989, x63990, x63991, x63992, x63993, x63994;
  wire x63995, x63996, x63997, x63998, x63999, x64000, x64001, x64002;
  wire x64003, x64004, x64005, x64006, x64007, x64008, x64010, x64011;
  wire x64012, x64013, x64014, x64015, x64016, x64017, x64018, x64019;
  wire x64020, x64021, x64022, x64023, x64024, x64025, x64026, x64027;
  wire x64028, x64029, x64030, x64031, x64032, x64033, x64034, x64035;
  wire x64036, x64037, x64038, x64039, x64040, x64041, x64042, x64043;
  wire x64044, x64045, x64046, x64047, x64048, x64049, x64050, x64051;
  wire x64052, x64053, x64054, x64055, x64056, x64057, x64058, x64059;
  wire x64060, x64061, x64062, x64063, x64064, x64065, x64066, x64067;
  wire x64068, x64069, x64070, x64071, x64072, x64073, x64074, x64075;
  wire x64076, x64077, x64078, x64079, x64080, x64081, x64082, x64083;
  wire x64084, x64085, x64086, x64087, x64088, x64089, x64090, x64091;
  wire x64092, x64093, x64094, x64095, x64096, x64097, x64098, x64099;
  wire x64100, x64101, x64103, x64104, x64105, x64106, x64107, x64108;
  wire x64109, x64110, x64111, x64112, x64113, x64114, x64115, x64116;
  wire x64117, x64118, x64119, x64120, x64121, x64122, x64123, x64124;
  wire x64125, x64126, x64127, x64128, x64129, x64130, x64131, x64132;
  wire x64133, x64134, x64135, x64136, x64137, x64138, x64139, x64140;
  wire x64141, x64142, x64143, x64144, x64145, x64146, x64147, x64148;
  wire x64149, x64150, x64151, x64152, x64153, x64154, x64155, x64156;
  wire x64157, x64158, x64159, x64160, x64161, x64162, x64163, x64164;
  wire x64165, x64166, x64167, x64168, x64169, x64170, x64171, x64172;
  wire x64173, x64174, x64175, x64176, x64177, x64178, x64179, x64180;
  wire x64181, x64182, x64183, x64184, x64185, x64186, x64187, x64188;
  wire x64189, x64190, x64192, x64193, x64194, x64195, x64196, x64197;
  wire x64198, x64199, x64200, x64201, x64202, x64203, x64204, x64205;
  wire x64206, x64207, x64208, x64209, x64210, x64211, x64212, x64213;
  wire x64214, x64215, x64216, x64217, x64218, x64219, x64220, x64221;
  wire x64222, x64223, x64224, x64225, x64226, x64227, x64228, x64229;
  wire x64230, x64231, x64232, x64233, x64234, x64235, x64236, x64237;
  wire x64238, x64239, x64240, x64241, x64242, x64243, x64244, x64245;
  wire x64246, x64247, x64248, x64249, x64250, x64251, x64252, x64253;
  wire x64254, x64255, x64256, x64257, x64258, x64259, x64260, x64261;
  wire x64262, x64263, x64264, x64265, x64266, x64267, x64268, x64269;
  wire x64270, x64271, x64273, x64274, x64275, x64276, x64277, x64278;
  wire x64279, x64280, x64281, x64282, x64283, x64284, x64285, x64286;
  wire x64287, x64288, x64289, x64290, x64291, x64292, x64293, x64294;
  wire x64295, x64296, x64297, x64298, x64299, x64300, x64301, x64302;
  wire x64303, x64304, x64305, x64306, x64307, x64308, x64309, x64310;
  wire x64311, x64312, x64313, x64314, x64315, x64316, x64317, x64318;
  wire x64319, x64320, x64321, x64322, x64323, x64324, x64325, x64326;
  wire x64327, x64328, x64329, x64330, x64331, x64332, x64333, x64334;
  wire x64335, x64336, x64338, x64340, x64342, x64344, x64346, x64348;
  wire x64350, x64352, x64354, x64356, x64358, x64360, x64362, x64364;
  wire x64366, x64368, x64370, x64372, x64374, x64376, x64378, x64380;
  wire x64382, x64384, x64386, x64388, x64390, x64392, x64394, x64396;
  wire x64398, x64399, x64400, x64401, x64402, x64403, x64404, x64405;
  wire x64406, x64407, x64408, x64409, x64410, x64411, x64412, x64413;
  wire x64414, x64415, x64416, x64417, x64418, x64419, x64420, x64421;
  wire x64422, x64423, x64424, x64425, x64426, x64427, x64428, x64430;
  wire x64431, x64432, x64434, x64435, x64437, x64439, x64440, x64442;
  wire x64444, x64445, x64447, x64449, x64450, x64452, x64454, x64455;
  wire x64457, x64459, x64460, x64462, x64464, x64465, x64467, x64469;
  wire x64470, x64472, x64474, x64475, x64485, x64486, x64487, x64488;
  wire x64489, x64491, x64492, x64493, x64495, x64496, x64497, x64499;
  wire x64500, x64501, x64503, x64504, x64505, x64507, x64508, x64509;
  wire x64511, x64512, x64513, x64516, x64518, x64519, x64521, x64522;
  wire x64524, x64525, x64527, x64529, x64530, x64532, x64534, x64535;
  wire x64537, x64539, x64540, x64542, x64544, x64545, x64548, x64550;
  wire x64551, x64553, x64554, x64556, x64557, x64559, x64560, x64562;
  wire x64563, x64566, x64568, x64569, x64570, x64571, x64572, x64573;
  wire x64575, x64577, x64578, x64580, x64581, x64582, x64584, x64586;
  wire x64587, x64589, x64591, x64592, x64594, x64596, x64597, x64599;
  wire x64600, x64601, x64603, x64605, x64606, x64645, x64647, x64648;
  wire x64649, x64650, x64651, x64652, x64653, x64654, x64655, x64656;
  wire x64657, x64658, x64659, x64660, x64661, x64662, x64663, x64664;
  wire x64665, x64666, x64667, x64668, x64669, x64670, x64671, x64672;
  wire x64673, x64674, x64675, x64676, x64677, x64678, x64679, x64680;
  wire x64681, x64682, x64683, x64684, x64685, x64686, x64687, x64688;
  wire x64689, x64690, x64691, x64692, x64693, x64694, x64695, x64696;
  wire x64697, x64698, x64699, x64700, x64701, x64702, x64703, x64704;
  wire x64705, x64706, x64707, x64708, x64709, x64710, x64711, x64712;
  wire x64713, x64714, x64715, x64716, x64717, x64718, x64719, x64720;
  wire x64721, x64722, x64723, x64724, x64725, x64726, x64727, x64728;
  wire x64729, x64730, x64731, x64732, x64733, x64734, x64735, x64736;
  wire x64737, x64738, x64739, x64740, x64742, x64743, x64744, x64745;
  wire x64746, x64747, x64748, x64749, x64750, x64751, x64752, x64753;
  wire x64754, x64755, x64756, x64757, x64758, x64759, x64760, x64761;
  wire x64762, x64763, x64764, x64765, x64766, x64767, x64768, x64769;
  wire x64770, x64771, x64772, x64773, x64774, x64775, x64776, x64777;
  wire x64778, x64779, x64780, x64781, x64782, x64783, x64784, x64785;
  wire x64786, x64787, x64788, x64789, x64790, x64791, x64792, x64793;
  wire x64794, x64795, x64796, x64797, x64798, x64799, x64800, x64801;
  wire x64802, x64803, x64804, x64805, x64806, x64807, x64808, x64809;
  wire x64810, x64811, x64812, x64813, x64814, x64815, x64816, x64817;
  wire x64818, x64819, x64820, x64821, x64822, x64823, x64824, x64825;
  wire x64826, x64827, x64828, x64829, x64830, x64831, x64832, x64833;
  wire x64835, x64836, x64837, x64838, x64839, x64840, x64841, x64842;
  wire x64843, x64844, x64845, x64846, x64847, x64848, x64849, x64850;
  wire x64851, x64852, x64853, x64854, x64855, x64856, x64857, x64858;
  wire x64859, x64860, x64861, x64862, x64863, x64864, x64865, x64866;
  wire x64867, x64868, x64869, x64870, x64871, x64872, x64873, x64874;
  wire x64875, x64876, x64877, x64878, x64879, x64880, x64881, x64882;
  wire x64883, x64884, x64885, x64886, x64887, x64888, x64889, x64890;
  wire x64891, x64892, x64893, x64894, x64895, x64896, x64897, x64898;
  wire x64899, x64900, x64901, x64902, x64903, x64904, x64905, x64906;
  wire x64907, x64908, x64909, x64910, x64911, x64912, x64913, x64914;
  wire x64915, x64916, x64917, x64918, x64919, x64920, x64921, x64922;
  wire x64924, x64925, x64926, x64927, x64928, x64929, x64930, x64931;
  wire x64932, x64933, x64934, x64935, x64936, x64937, x64938, x64939;
  wire x64940, x64941, x64942, x64943, x64944, x64945, x64946, x64947;
  wire x64948, x64949, x64950, x64951, x64952, x64953, x64954, x64955;
  wire x64956, x64957, x64958, x64959, x64960, x64961, x64962, x64963;
  wire x64964, x64965, x64966, x64967, x64968, x64969, x64970, x64971;
  wire x64972, x64973, x64974, x64975, x64976, x64977, x64978, x64979;
  wire x64980, x64981, x64982, x64983, x64984, x64985, x64986, x64987;
  wire x64988, x64989, x64990, x64991, x64992, x64993, x64994, x64995;
  wire x64996, x64997, x64998, x64999, x65000, x65001, x65002, x65003;
  wire x65005, x65006, x65007, x65008, x65009, x65010, x65011, x65012;
  wire x65013, x65014, x65015, x65016, x65017, x65018, x65019, x65020;
  wire x65021, x65022, x65023, x65024, x65025, x65026, x65027, x65028;
  wire x65029, x65030, x65031, x65032, x65033, x65034, x65035, x65036;
  wire x65037, x65038, x65039, x65040, x65041, x65042, x65043, x65044;
  wire x65045, x65046, x65047, x65048, x65049, x65050, x65051, x65052;
  wire x65053, x65054, x65055, x65056, x65057, x65058, x65059, x65060;
  wire x65061, x65062, x65063, x65064, x65065, x65066, x65067, x65068;
  wire x65069, x65070, x65071, x65072, x65073, x65074, x65075, x65076;
  wire x65077, x65078, x65079, x65080, x65081, x65082, x65083, x65084;
  wire x65085, x65086, x65087, x65088, x65089, x65090, x65091, x65092;
  wire x65093, x65094, x65095, x65096, x65097, x65098, x65100, x65101;
  wire x65102, x65104, x65105, x65107, x65109, x65110, x65112, x65114;
  wire x65115, x65117, x65119, x65120, x65122, x65124, x65125, x65127;
  wire x65129, x65130, x65132, x65134, x65135, x65137, x65139, x65140;
  wire x65142, x65144, x65145, x65155, x65156, x65157, x65158, x65159;
  wire x65161, x65162, x65163, x65165, x65166, x65167, x65169, x65170;
  wire x65171, x65173, x65174, x65175, x65177, x65178, x65179, x65181;
  wire x65182, x65183, x65186, x65188, x65189, x65191, x65192, x65194;
  wire x65195, x65197, x65199, x65200, x65202, x65204, x65205, x65207;
  wire x65209, x65210, x65212, x65214, x65215, x65218, x65220, x65221;
  wire x65223, x65224, x65226, x65227, x65229, x65230, x65232, x65233;
  wire x65236, x65238, x65239, x65240, x65241, x65242, x65243, x65245;
  wire x65247, x65248, x65250, x65251, x65252, x65254, x65256, x65257;
  wire x65259, x65261, x65262, x65264, x65266, x65267, x65269, x65270;
  wire x65271, x65273, x65275, x65276, x65315, x65317, x65318, x65319;
  wire x65320, x65321, x65322, x65323, x65324, x65325, x65326, x65327;
  wire x65328, x65329, x65330, x65331, x65332, x65333, x65334, x65335;
  wire x65336, x65337, x65338, x65339, x65340, x65341, x65342, x65343;
  wire x65344, x65345, x65346, x65347, x65348, x65349, x65350, x65351;
  wire x65352, x65353, x65354, x65355, x65356, x65357, x65358, x65359;
  wire x65360, x65361, x65362, x65363, x65364, x65365, x65366, x65367;
  wire x65368, x65369, x65370, x65371, x65372, x65373, x65374, x65375;
  wire x65376, x65377, x65378, x65379, x65380, x65381, x65382, x65383;
  wire x65384, x65385, x65386, x65387, x65388, x65389, x65390, x65391;
  wire x65392, x65393, x65394, x65395, x65396, x65397, x65398, x65399;
  wire x65400, x65401, x65402, x65403, x65404, x65405, x65406, x65407;
  wire x65408, x65409, x65410, x65412, x65413, x65414, x65415, x65416;
  wire x65417, x65418, x65419, x65420, x65421, x65422, x65423, x65424;
  wire x65425, x65426, x65427, x65428, x65429, x65430, x65431, x65432;
  wire x65433, x65434, x65435, x65436, x65437, x65438, x65439, x65440;
  wire x65441, x65442, x65443, x65444, x65445, x65446, x65447, x65448;
  wire x65449, x65450, x65451, x65452, x65453, x65454, x65455, x65456;
  wire x65457, x65458, x65459, x65460, x65461, x65462, x65463, x65464;
  wire x65465, x65466, x65467, x65468, x65469, x65470, x65471, x65472;
  wire x65473, x65474, x65475, x65476, x65477, x65478, x65479, x65480;
  wire x65481, x65482, x65483, x65484, x65485, x65486, x65487, x65488;
  wire x65489, x65490, x65491, x65492, x65493, x65494, x65495, x65496;
  wire x65497, x65498, x65499, x65500, x65501, x65502, x65503, x65505;
  wire x65506, x65507, x65508, x65509, x65510, x65511, x65512, x65513;
  wire x65514, x65515, x65516, x65517, x65518, x65519, x65520, x65521;
  wire x65522, x65523, x65524, x65525, x65526, x65527, x65528, x65529;
  wire x65530, x65531, x65532, x65533, x65534, x65535, x65536, x65537;
  wire x65538, x65539, x65540, x65541, x65542, x65543, x65544, x65545;
  wire x65546, x65547, x65548, x65549, x65550, x65551, x65552, x65553;
  wire x65554, x65555, x65556, x65557, x65558, x65559, x65560, x65561;
  wire x65562, x65563, x65564, x65565, x65566, x65567, x65568, x65569;
  wire x65570, x65571, x65572, x65573, x65574, x65575, x65576, x65577;
  wire x65578, x65579, x65580, x65581, x65582, x65583, x65584, x65585;
  wire x65586, x65587, x65588, x65589, x65590, x65591, x65592, x65594;
  wire x65595, x65596, x65597, x65598, x65599, x65600, x65601, x65602;
  wire x65603, x65604, x65605, x65606, x65607, x65608, x65609, x65610;
  wire x65611, x65612, x65613, x65614, x65615, x65616, x65617, x65618;
  wire x65619, x65620, x65621, x65622, x65623, x65624, x65625, x65626;
  wire x65627, x65628, x65629, x65630, x65631, x65632, x65633, x65634;
  wire x65635, x65636, x65637, x65638, x65639, x65640, x65641, x65642;
  wire x65643, x65644, x65645, x65646, x65647, x65648, x65649, x65650;
  wire x65651, x65652, x65653, x65654, x65655, x65656, x65657, x65658;
  wire x65659, x65660, x65661, x65662, x65663, x65664, x65665, x65666;
  wire x65667, x65668, x65669, x65670, x65671, x65672, x65673, x65675;
  wire x65676, x65677, x65678, x65679, x65680, x65681, x65682, x65683;
  wire x65684, x65685, x65686, x65687, x65688, x65689, x65690, x65691;
  wire x65692, x65693, x65694, x65695, x65696, x65697, x65698, x65699;
  wire x65700, x65701, x65702, x65703, x65704, x65705, x65706, x65707;
  wire x65708, x65709, x65710, x65711, x65712, x65713, x65714, x65715;
  wire x65716, x65717, x65718, x65719, x65720, x65721, x65722, x65723;
  wire x65724, x65725, x65726, x65727, x65728, x65729, x65730, x65731;
  wire x65732, x65733, x65734, x65735, x65736, x65737, x65738, x65739;
  wire x65740, x65741, x65742, x65743, x65744, x65745, x65746, x65747;
  wire x65748, x65749, x65750, x65751, x65752, x65753, x65754, x65755;
  wire x65756, x65757, x65758, x65759, x65760, x65761, x65762, x65763;
  wire x65764, x65765, x65766, x65767, x65768, x65770, x65771, x65772;
  wire x65774, x65775, x65777, x65779, x65780, x65782, x65784, x65785;
  wire x65787, x65789, x65790, x65792, x65794, x65795, x65797, x65799;
  wire x65800, x65802, x65804, x65805, x65807, x65809, x65810, x65812;
  wire x65814, x65815, x65825, x65826, x65827, x65828, x65829, x65831;
  wire x65832, x65833, x65835, x65836, x65837, x65839, x65840, x65841;
  wire x65843, x65844, x65845, x65847, x65848, x65849, x65851, x65852;
  wire x65853, x65856, x65858, x65859, x65861, x65862, x65864, x65865;
  wire x65867, x65869, x65870, x65872, x65874, x65875, x65877, x65879;
  wire x65880, x65882, x65884, x65885, x65888, x65890, x65891, x65893;
  wire x65894, x65896, x65897, x65899, x65900, x65902, x65903, x65906;
  wire x65908, x65909, x65910, x65911, x65912, x65913, x65915, x65917;
  wire x65918, x65920, x65921, x65922, x65924, x65926, x65927, x65929;
  wire x65931, x65932, x65934, x65936, x65937, x65939, x65940, x65941;
  wire x65943, x65945, x65946, x65985, x65987, x65988, x65989, x65990;
  wire x65991, x65992, x65993, x65994, x65995, x65996, x65997, x65998;
  wire x65999, x66000, x66001, x66002, x66003, x66004, x66005, x66006;
  wire x66007, x66008, x66009, x66010, x66011, x66012, x66013, x66014;
  wire x66015, x66016, x66017, x66018, x66019, x66020, x66021, x66022;
  wire x66023, x66024, x66025, x66026, x66027, x66028, x66029, x66030;
  wire x66031, x66032, x66033, x66034, x66035, x66036, x66037, x66038;
  wire x66039, x66040, x66041, x66042, x66043, x66044, x66045, x66046;
  wire x66047, x66048, x66049, x66050, x66051, x66052, x66053, x66054;
  wire x66055, x66056, x66057, x66058, x66059, x66060, x66061, x66062;
  wire x66063, x66064, x66065, x66066, x66067, x66068, x66069, x66070;
  wire x66071, x66072, x66073, x66074, x66075, x66076, x66077, x66078;
  wire x66079, x66080, x66082, x66083, x66084, x66085, x66086, x66087;
  wire x66088, x66089, x66090, x66091, x66092, x66093, x66094, x66095;
  wire x66096, x66097, x66098, x66099, x66100, x66101, x66102, x66103;
  wire x66104, x66105, x66106, x66107, x66108, x66109, x66110, x66111;
  wire x66112, x66113, x66114, x66115, x66116, x66117, x66118, x66119;
  wire x66120, x66121, x66122, x66123, x66124, x66125, x66126, x66127;
  wire x66128, x66129, x66130, x66131, x66132, x66133, x66134, x66135;
  wire x66136, x66137, x66138, x66139, x66140, x66141, x66142, x66143;
  wire x66144, x66145, x66146, x66147, x66148, x66149, x66150, x66151;
  wire x66152, x66153, x66154, x66155, x66156, x66157, x66158, x66159;
  wire x66160, x66161, x66162, x66163, x66164, x66165, x66166, x66167;
  wire x66168, x66169, x66170, x66171, x66172, x66173, x66175, x66176;
  wire x66177, x66178, x66179, x66180, x66181, x66182, x66183, x66184;
  wire x66185, x66186, x66187, x66188, x66189, x66190, x66191, x66192;
  wire x66193, x66194, x66195, x66196, x66197, x66198, x66199, x66200;
  wire x66201, x66202, x66203, x66204, x66205, x66206, x66207, x66208;
  wire x66209, x66210, x66211, x66212, x66213, x66214, x66215, x66216;
  wire x66217, x66218, x66219, x66220, x66221, x66222, x66223, x66224;
  wire x66225, x66226, x66227, x66228, x66229, x66230, x66231, x66232;
  wire x66233, x66234, x66235, x66236, x66237, x66238, x66239, x66240;
  wire x66241, x66242, x66243, x66244, x66245, x66246, x66247, x66248;
  wire x66249, x66250, x66251, x66252, x66253, x66254, x66255, x66256;
  wire x66257, x66258, x66259, x66260, x66261, x66262, x66264, x66265;
  wire x66266, x66267, x66268, x66269, x66270, x66271, x66272, x66273;
  wire x66274, x66275, x66276, x66277, x66278, x66279, x66280, x66281;
  wire x66282, x66283, x66284, x66285, x66286, x66287, x66288, x66289;
  wire x66290, x66291, x66292, x66293, x66294, x66295, x66296, x66297;
  wire x66298, x66299, x66300, x66301, x66302, x66303, x66304, x66305;
  wire x66306, x66307, x66308, x66309, x66310, x66311, x66312, x66313;
  wire x66314, x66315, x66316, x66317, x66318, x66319, x66320, x66321;
  wire x66322, x66323, x66324, x66325, x66326, x66327, x66328, x66329;
  wire x66330, x66331, x66332, x66333, x66334, x66335, x66336, x66337;
  wire x66338, x66339, x66340, x66341, x66342, x66343, x66345, x66346;
  wire x66347, x66348, x66349, x66350, x66351, x66352, x66353, x66354;
  wire x66355, x66356, x66357, x66358, x66359, x66360, x66361, x66362;
  wire x66363, x66364, x66365, x66366, x66367, x66368, x66369, x66370;
  wire x66371, x66372, x66373, x66374, x66375, x66376, x66377, x66378;
  wire x66379, x66380, x66381, x66382, x66383, x66384, x66385, x66386;
  wire x66387, x66388, x66389, x66390, x66391, x66392, x66393, x66394;
  wire x66395, x66396, x66397, x66398, x66399, x66400, x66401, x66402;
  wire x66403, x66404, x66405, x66406, x66407, x66408, x66410, x66411;
  wire x66412, x66414, x66415, x66416, x66418, x66419, x66420, x66422;
  wire x66423, x66424, x66426, x66427, x66428, x66430, x66431, x66432;
  wire x66434, x66435, x66436, x66438, x66439, x66440, x66442, x66443;
  wire x66444, x66446, x66447, x66448, x66450, x66451, x66452, x66454;
  wire x66455, x66456, x66458, x66459, x66460, x66462, x66463, x66464;
  wire x66466, x66467, x66468, x66471, x66602, x66604, x66605, x66606;
  wire x66607, x66608, x66609, x66610, x66611, x66612, x66613, x66614;
  wire x66615, x66616, x66617, x66618, x66619, x66620, x66621, x66622;
  wire x66623, x66624, x66625, x66626, x66627, x66628, x66629, x66630;
  wire x66631, x66632, x66633, x66634, x66635, x66636, x66637, x66638;
  wire x66639, x66640, x66641, x66642, x66643, x66644, x66645, x66646;
  wire x66647, x66648, x66649, x66650, x66651, x66652, x66653, x66654;
  wire x66655, x66656, x66657, x66658, x66659, x66660, x66661, x66662;
  wire x66663, x66664, x66665, x66666, x66667, x66668, x66669, x66670;
  wire x66671, x66672, x66673, x66674, x66675, x66676, x66677, x66678;
  wire x66679, x66680, x66681, x66682, x66683, x66684, x66685, x66686;
  wire x66687, x66688, x66689, x66690, x66691, x66692, x66693, x66694;
  wire x66695, x66696, x66697, x66698, x66699, x66700, x66701, x66702;
  wire x66703, x66704, x66705, x66706, x66707, x66708, x66709, x66710;
  wire x66711, x66712, x66713, x66714, x66715, x66716, x66717, x66718;
  wire x66719, x66720, x66721, x66722, x66723, x66724, x66725, x66726;
  wire x66727, x66728, x66729, x66730, x66731, x66732, x66733, x66734;
  wire x66735, x66736, x66737, x66738, x66739, x66740, x66741, x66742;
  wire x66743, x66744, x66745, x66746, x66747, x66748, x66749, x66750;
  wire x66751, x66752, x66753, x66754, x66755, x66756, x66757, x66758;
  wire x66759, x66760, x66761, x66762, x66763, x66764, x66765, x66766;
  wire x66767, x66768, x66769, x66770, x66771, x66772, x66773, x66774;
  wire x66775, x66776, x66777, x66778, x66779, x66780, x66781, x66782;
  wire x66783, x66784, x66785, x66786, x66787, x66788, x66789, x66790;
  wire x66791, x66792, x66793, x66794, x66795, x66796, x66797, x66798;
  wire x66799, x66800, x66801, x66802, x66803, x66804, x66805, x66806;
  wire x66807, x66808, x66809, x66810, x66811, x66812, x66813, x66814;
  wire x66815, x66816, x66817, x66818, x66819, x66820, x66821, x66822;
  wire x66823, x66824, x66825, x66826, x66827, x66828, x66829, x66830;
  wire x66831, x66832, x66833, x66834, x66835, x66836, x66837, x66838;
  wire x66839, x66840, x66841, x66842, x66843, x66844, x66845, x66846;
  wire x66847, x66848, x66849, x66850, x66851, x66852, x66853, x66854;
  wire x66855, x66856, x66857, x66858, x66859, x66860, x66861, x66862;
  wire x66863, x66864, x66865, x66866, x66867, x66868, x66869, x66870;
  wire x66871, x66872, x66873, x66874, x66875, x66876, x66877, x66878;
  wire x66879, x66880, x66881, x66882, x66883, x66884, x66885, x66886;
  wire x66887, x66888, x66889, x66890, x66891, x66892, x66893, x66895;
  wire x66896, x66897, x66899, x66900, x66901, x66903, x66904, x66905;
  wire x66907, x66908, x66909, x66911, x66912, x66913, x66915, x66916;
  wire x66917, x66919, x66920, x66921, x66923, x66924, x66925, x66927;
  wire x66928, x66929, x66931, x66932, x66933, x66935, x66936, x66937;
  wire x66939, x66940, x66941, x66943, x66944, x66945, x66947, x66948;
  wire x66949, x66951, x66952, x66953, x66955, x66956, x66957, x66959;
  wire x66960, x66961, x66963, x66964, x66965, x66967, x66968, x66969;
  wire x66971, x66972, x66973, x66975, x66976, x66977, x66979, x66980;
  wire x66981, x66983, x66984, x66985, x66987, x66988, x66989, x66991;
  wire x66992, x66993, x66995, x66996, x66997, x66999, x67000, x67001;
  wire x67003, x67004, x67005, x67007, x67008, x67009, x67011, x67012;
  wire x67013, x67015, x67016, x67017, x67019, x67020, x67021, x67023;
  wire x67024, x67025, x67027, x67028, x67029, x67031, x67032, x67033;
  wire x67035, x67036, x67037, x67039, x67040, x67041, x67043, x67044;
  wire x67045, x67047, x67048, x67049, x67051, x67052, x67053, x67055;
  wire x67056, x67057, x67059, x67060, x67061, x67063, x67064, x67065;
  wire x67067, x67068, x67069, x67071, x67072, x67073, x67075, x67076;
  wire x67077, x67079, x67080, x67081, x67083, x67084, x67085, x67087;
  wire x67088, x67089, x67091, x67092, x67093, x67095, x67096, x67097;
  wire x67099, x67100, x67101, x67103, x67104, x67105, x67107, x67108;
  wire x67109, x67111, x67112, x67113, x67115, x67116, x67117, x67119;
  wire x67120, x67121, x67123, x67124, x67125, x67127, x67128, x67129;
  wire x67131, x67132, x67133, x67135, x67136, x67137, x67139, x67140;
  wire x67141, x67143, x67144, x67145, x67147, x67148, x67149, x67151;
  wire x67152, x67153, x67155, x67156, x67157, x67159, x67160, x67161;
  wire x67163, x67164, x67165, x67167, x67168, x67169, x67171, x67172;
  wire x67173, x67175, x67176, x67177, x67179, x67180, x67181, x67183;
  wire x67184, x67185, x67187, x67188, x67189, x67191, x67192, x67193;
  wire x67195, x67196, x67197, x67199, x67200, x67201, x67203, x67204;
  wire x67205, x67207, x67208, x67209, x67211, x67212, x67213, x67215;
  wire x67216, x67217, x67219, x67220, x67221, x67223, x67224, x67225;
  wire x67227, x67228, x67229, x67231, x67232, x67233, x67235, x67236;
  wire x67237, x67239, x67240, x67241, x67243, x67244, x67245, x67247;
  wire x67248, x67249, x67251, x67252, x67253, x67255, x67256, x67257;
  wire x67259, x67260, x67261, x67263, x67264, x67265, x67267, x67268;
  wire x67269, x67271, x67272, x67273, x67275, x67276, x67277, x67279;
  wire x67280, x67281, x67283, x67284, x67285, x67287, x67288, x67289;
  wire x67291, x67292, x67293, x67295, x67296, x67297, x67299, x67300;
  wire x67301, x67303, x67304, x67305, x67307, x67308, x67309, x67311;
  wire x67312, x67313, x67315, x67316, x67317, x67319, x67320, x67321;
  wire x67323, x67324, x67325, x67327, x67328, x67329, x67331, x67332;
  wire x67333, x67335, x67336, x67337, x67339, x67340, x67341, x67343;
  wire x67344, x67345, x67347, x67348, x67349, x67351, x67352, x67353;
  wire x67355, x67356, x67357, x67359, x67360, x67361, x67363, x67364;
  wire x67365, x67367, x67368, x67369, x67371, x67372, x67373, x67375;
  wire x67376, x67377, x67379, x67380, x67381, x67383, x67384, x67385;
  wire x67387, x67388, x67389, x67391, x67392, x67393, x67395, x67396;
  wire x67397, x67399, x67400, x67401, x67403, x67404, x67406, x67407;
  wire x67408, x67410, x67411, x67412, x67414, x67415, x67416, x67418;
  wire x67419, x67420, x67422, x67423, x67424, x67426, x67427, x67428;
  wire x67430, x67431, x67432, x67434, x67435, x67436, x67438, x67439;
  wire x67440, x67442, x67443, x67444, x67446, x67447, x67448, x67450;
  wire x67451, x67452, x67454, x67455, x67456, x67458, x67459, x67460;
  wire x67462, x67464, x67595, x67597, x67598, x67599, x67600, x67601;
  wire x67602, x67603, x67604, x67605, x67606, x67607, x67608, x67609;
  wire x67610, x67611, x67612, x67613, x67614, x67615, x67616, x67617;
  wire x67618, x67619, x67620, x67621, x67622, x67623, x67624, x67625;
  wire x67626, x67627, x67628, x67629, x67630, x67631, x67632, x67633;
  wire x67634, x67635, x67636, x67637, x67638, x67639, x67640, x67641;
  wire x67642, x67643, x67644, x67645, x67646, x67647, x67648, x67649;
  wire x67650, x67651, x67652, x67653, x67654, x67655, x67656, x67657;
  wire x67658, x67659, x67660, x67661, x67662, x67663, x67664, x67665;
  wire x67666, x67667, x67668, x67669, x67670, x67671, x67672, x67673;
  wire x67674, x67675, x67676, x67677, x67678, x67679, x67680, x67681;
  wire x67682, x67683, x67684, x67685, x67686, x67687, x67688, x67689;
  wire x67690, x67691, x67692, x67693, x67694, x67695, x67696, x67697;
  wire x67698, x67699, x67700, x67701, x67702, x67703, x67704, x67705;
  wire x67706, x67707, x67708, x67709, x67710, x67711, x67712, x67713;
  wire x67714, x67715, x67716, x67717, x67718, x67719, x67720, x67721;
  wire x67722, x67723, x67724, x67725, x67726, x67727, x67728, x67729;
  wire x67730, x67731, x67732, x67733, x67734, x67735, x67736, x67737;
  wire x67738, x67739, x67740, x67741, x67742, x67743, x67744, x67745;
  wire x67746, x67747, x67748, x67749, x67750, x67751, x67752, x67753;
  wire x67754, x67755, x67756, x67757, x67758, x67759, x67760, x67761;
  wire x67762, x67763, x67764, x67765, x67766, x67767, x67768, x67769;
  wire x67770, x67771, x67772, x67773, x67774, x67775, x67776, x67777;
  wire x67778, x67779, x67780, x67781, x67782, x67783, x67784, x67785;
  wire x67786, x67787, x67788, x67789, x67790, x67791, x67792, x67793;
  wire x67794, x67795, x67796, x67797, x67798, x67799, x67800, x67801;
  wire x67802, x67803, x67804, x67805, x67806, x67807, x67808, x67809;
  wire x67810, x67811, x67812, x67813, x67814, x67815, x67816, x67817;
  wire x67818, x67819, x67820, x67821, x67822, x67823, x67824, x67825;
  wire x67826, x67827, x67828, x67829, x67830, x67831, x67832, x67833;
  wire x67834, x67835, x67836, x67837, x67838, x67839, x67840, x67841;
  wire x67842, x67843, x67844, x67845, x67846, x67847, x67848, x67849;
  wire x67850, x67851, x67852, x67853, x67854, x67855, x67856, x67857;
  wire x67858, x67859, x67860, x67861, x67862, x67863, x67864, x67865;
  wire x67866, x67867, x67868, x67869, x67870, x67871, x67872, x67873;
  wire x67874, x67875, x67876, x67877, x67878, x67879, x67880, x67881;
  wire x67882, x67883, x67884, x67885, x67886, x67888, x67889, x67890;
  wire x67892, x67893, x67894, x67896, x67897, x67898, x67900, x67901;
  wire x67902, x67904, x67905, x67906, x67908, x67909, x67910, x67912;
  wire x67913, x67914, x67916, x67917, x67918, x67920, x67921, x67922;
  wire x67924, x67925, x67926, x67928, x67929, x67930, x67932, x67933;
  wire x67934, x67936, x67937, x67938, x67940, x67941, x67942, x67944;
  wire x67945, x67946, x67948, x67949, x67950, x67952, x67953, x67954;
  wire x67956, x67957, x67958, x67960, x67961, x67962, x67964, x67965;
  wire x67966, x67968, x67969, x67970, x67972, x67973, x67974, x67976;
  wire x67977, x67978, x67980, x67981, x67982, x67984, x67985, x67986;
  wire x67988, x67989, x67990, x67992, x67993, x67994, x67996, x67997;
  wire x67998, x68000, x68001, x68002, x68004, x68005, x68006, x68008;
  wire x68009, x68010, x68012, x68013, x68014, x68016, x68017, x68018;
  wire x68020, x68021, x68022, x68024, x68025, x68026, x68028, x68029;
  wire x68030, x68032, x68033, x68034, x68036, x68037, x68038, x68040;
  wire x68041, x68042, x68044, x68045, x68046, x68048, x68049, x68050;
  wire x68052, x68053, x68054, x68056, x68057, x68058, x68060, x68061;
  wire x68062, x68064, x68065, x68066, x68068, x68069, x68070, x68072;
  wire x68073, x68074, x68076, x68077, x68078, x68080, x68081, x68082;
  wire x68084, x68085, x68086, x68088, x68089, x68090, x68092, x68093;
  wire x68094, x68096, x68097, x68098, x68100, x68101, x68102, x68104;
  wire x68105, x68106, x68108, x68109, x68110, x68112, x68113, x68114;
  wire x68116, x68117, x68118, x68120, x68121, x68122, x68124, x68125;
  wire x68126, x68128, x68129, x68130, x68132, x68133, x68134, x68136;
  wire x68137, x68138, x68140, x68141, x68142, x68144, x68145, x68146;
  wire x68148, x68149, x68150, x68152, x68153, x68154, x68156, x68157;
  wire x68158, x68160, x68161, x68162, x68164, x68165, x68166, x68168;
  wire x68169, x68170, x68172, x68173, x68174, x68176, x68177, x68178;
  wire x68180, x68181, x68182, x68184, x68185, x68186, x68188, x68189;
  wire x68190, x68192, x68193, x68194, x68196, x68197, x68198, x68200;
  wire x68201, x68202, x68204, x68205, x68206, x68208, x68209, x68210;
  wire x68212, x68213, x68214, x68216, x68217, x68218, x68220, x68221;
  wire x68222, x68224, x68225, x68226, x68228, x68229, x68230, x68232;
  wire x68233, x68234, x68236, x68237, x68238, x68240, x68241, x68242;
  wire x68244, x68245, x68246, x68248, x68249, x68250, x68252, x68253;
  wire x68254, x68256, x68257, x68258, x68260, x68261, x68262, x68264;
  wire x68265, x68266, x68268, x68269, x68270, x68272, x68273, x68274;
  wire x68276, x68277, x68278, x68280, x68281, x68282, x68284, x68285;
  wire x68286, x68288, x68289, x68290, x68292, x68293, x68294, x68296;
  wire x68297, x68298, x68300, x68301, x68302, x68304, x68305, x68306;
  wire x68308, x68309, x68310, x68312, x68313, x68314, x68316, x68317;
  wire x68318, x68320, x68321, x68322, x68324, x68325, x68326, x68328;
  wire x68329, x68330, x68332, x68333, x68334, x68336, x68337, x68338;
  wire x68340, x68341, x68342, x68344, x68345, x68346, x68348, x68349;
  wire x68350, x68352, x68353, x68354, x68356, x68357, x68358, x68360;
  wire x68361, x68362, x68364, x68365, x68366, x68368, x68369, x68370;
  wire x68372, x68373, x68374, x68376, x68377, x68378, x68380, x68381;
  wire x68382, x68384, x68385, x68386, x68388, x68389, x68390, x68392;
  wire x68393, x68394, x68396, x68397, x68399, x68400, x68401, x68403;
  wire x68404, x68405, x68407, x68408, x68409, x68411, x68412, x68413;
  wire x68415, x68416, x68417, x68419, x68420, x68421, x68423, x68424;
  wire x68425, x68427, x68428, x68429, x68431, x68432, x68433, x68435;
  wire x68436, x68437, x68439, x68440, x68441, x68443, x68444, x68445;
  wire x68447, x68448, x68449, x68451, x68452, x68453, x68455, x68456;
  wire x68457, x68460, x68462, x68463, x68465, x68466, x68468, x68472;
  wire x68474, x68476, x68477, x68479, x68481, x68482, x68484, x68486;
  wire x68487, x68489, x68490, x68492, x68493, x68495, x68496, x68497;
  wire x68499, x68500, x68503, x68504, x68506, x68507, x68508, x68510;
  wire x68512, x68513, x68515, x68517, x68518, x68520, x68522, x68523;
  wire x68525, x68527, x68528, x68531, x68532, x68534, x68536, x68538;
  wire x68539, x68540, x68542, x68543, x68544, x68546, x68547, x68548;
  wire x68550, x68551, x68552, x68554, x68555, x68556, x68558, x68559;
  wire x68560, x68562, x68564, x68565, x68566, x68567, x68568, x68569;
  wire x68571, x68572, x68573, x68574, x68575, x68576, x68577, x68578;
  wire x68579, x68580, x68581, x68582, x68583, x68584, x68585, x68586;
  wire x68587, x68588, x68589, x68590, x68591, x68592, x68593, x68594;
  wire x68595, x68596, x68597, x68598, x68599, x68600, x68601, x68602;
  wire x68603, x68604, x68605, x68606, x68607, x68608, x68609, x68610;
  wire x68611, x68612, x68613, x68614, x68615, x68616, x68617, x68630;
  wire x68631, x68632, x68633, x68634, x68635, x68636, x68637, x68638;
  wire x68642, x68644, x68645, x68646, x68647, x68648, x68649, x68650;
  wire x68651, x68652, x68653, x68657, x68659, x68664, x68665, x68666;
  wire x68667, x68668, x68669, x68670, x68672, x68673, x68674, x68675;
  wire x68676, x68678, x68680, x68685, x68686, x68687, x68688, x68689;
  wire x68690, x68691, x68693, x68694, x68695, x68696, x68697, x68699;
  wire x68701, x68704, x68705, x68706, x68707, x68708, x68709, x68710;
  wire x68711, x68712, x68713, x68714, x68715, x68716, x68717, x68718;
  wire x68719, x68722, x68723, x68724, x68725, x68726, x68727, x68728;
  wire x68729, x68730, x68731, x68732, x68733, x68734, x68735, x68736;
  wire x68737, x68738, x68739, x68740, x68741, x68742, x68743, x68744;
  wire x68746, x68747, x68748, x68749, x68750, x68751, x68752, x68753;
  wire x68754, x68755, x68756, x68757, x68758, x68759, x68760, x68761;
  wire x68762, x68763, x68764, x68765, x68766, x68767, x68768, x68769;
  wire x68770, x68771, x68772, x68773, x68774, x68775, x68776, x68777;
  wire x68778, x68779, x68780, x68781, x68782, x68783, x68784, x68785;
  wire x68786, x68787, x68788, x68789, x68790, x68791, x68792, x68793;
  wire x68794, x68795, x68796, x68797, x68798, x68799, x68800, x68801;
  wire x68802, x68803, x68804, x68805, x68806, x68807, x68808, x68809;
  wire x68811, x68812, x68813, x68814, x68815, x68816, x68817, x68818;
  wire x68819, x68820, x68821, x68822, x68823, x68824, x68825, x68826;
  wire x68827, x68828, x68829, x68830, x68831, x68832, x68833, x68834;
  wire x68835, x68836, x68837, x68838, x68839, x68840, x68841, x68842;
  wire x68843, x68844, x68845, x68846, x68847, x68848, x68849, x68850;
  wire x68851, x68852, x68853, x68854, x68855, x68856, x68857, x68858;
  wire x68859, x68860, x68861, x68862, x68863, x68864, x68865, x68866;
  wire x68867, x68868, x68869, x68870, x68871, x68872, x68873, x68874;
  wire x68875, x68876, x68877, x68878, x68879, x68880, x68881, x68882;
  wire x68883, x68884, x68885, x68886, x68887, x68888, x68889, x68890;
  wire x68891, x68892, x68893, x68894, x68895, x68896, x68897, x68898;
  wire x68899, x68900, x68901, x68902, x68903, x68904, x68905, x68906;
  wire x68907, x68908, x68909, x68910, x68911, x68912, x68913, x68914;
  wire x68915, x68916, x68917, x68918, x68919, x68920, x68921, x68922;
  wire x68923, x68924, x68925, x68926, x68927, x68928, x68929, x68930;
  wire x68931, x68932, x68933, x68934, x68935, x68936, x68937, x68938;
  wire x68939, x68940, x68941, x68942, x68943, x68944, x68945, x68946;
  wire x68947, x68948, x68949, x68950, x68951, x68952, x68953, x68954;
  wire x68955, x68956, x68957, x68958, x68959, x68960, x68961, x68962;
  wire x68963, x68964, x68965, x68966, x68967, x68968, x68969, x68970;
  wire x68971, x68972, x68973, x68974, x68975, x68976, x68977, x68978;
  wire x68979, x68980, x68981, x68982, x68983, x68984, x68985, x68986;
  wire x68987, x68988, x68989, x68990, x68991, x68992, x68993, x68994;
  wire x68995, x68996, x68997, x68998, x68999, x69000, x69001, x69002;
  wire x69003, x69004, x69005, x69006, x69007, x69008, x69009, x69010;
  wire x69011, x69012, x69013, x69014, x69015, x69016, x69017, x69018;
  wire x69019, x69020, x69021, x69022, x69023, x69024, x69025, x69026;
  wire x69027, x69028, x69029, x69030, x69031, x69032, x69033, x69034;
  wire x69035, x69036, x69037, x69038, x69039, x69040, x69041, x69042;
  wire x69043, x69044, x69045, x69046, x69047, x69048, x69049, x69050;
  wire x69051, x69052, x69053, x69054, x69055, x69056, x69057, x69058;
  wire x69059, x69060, x69061, x69062, x69063, x69064, x69065, x69066;
  wire x69067, x69068, x69069, x69070, x69071, x69072, x69073, x69074;
  wire x69075, x69076, x69077, x69078, x69079, x69080, x69081, x69082;
  wire x69083, x69084, x69085, x69086, x69087, x69088, x69089, x69090;
  wire x69091, x69092, x69093, x69094, x69095, x69096, x69097, x69098;
  wire x69099, x69100, x69101, x69102, x69103, x69104, x69105, x69106;
  wire x69107, x69108, x69109, x69110, x69111, x69112, x69113, x69114;
  wire x69115, x69116, x69117, x69118, x69119, x69120, x69121, x69122;
  wire x69123, x69124, x69125, x69126, x69127, x69128, x69129, x69130;
  wire x69131, x69132, x69133, x69134, x69135, x69136, x69137, x69138;
  wire x69139, x69140, x69141, x69142, x69143, x69144, x69145, x69146;
  wire x69147, x69148, x69149, x69150, x69151, x69152, x69153, x69154;
  wire x69155, x69156, x69157, x69158, x69159, x69160, x69161, x69162;
  wire x69163, x69164, x69165, x69166, x69167, x69168, x69169, x69170;
  wire x69171, x69172, x69173, x69174, x69175, x69176, x69177, x69178;
  wire x69179, x69180, x69181, x69182, x69183, x69184, x69185, x69186;
  wire x69187, x69188, x69189, x69190, x69191, x69192, x69193, x69194;
  wire x69195, x69196, x69197, x69198, x69199, x69200, x69201, x69202;
  wire x69203, x69204, x69205, x69206, x69207, x69208, x69209, x69210;
  wire x69211, x69212, x69213, x69214, x69215, x69216, x69217, x69218;
  wire x69219, x69220, x69221, x69222, x69223, x69224, x69225, x69226;
  wire x69227, x69228, x69229, x69230, x69231, x69232, x69233, x69234;
  wire x69235, x69236, x69237, x69238, x69239, x69240, x69241, x69242;
  wire x69243, x69244, x69245, x69246, x69247, x69248, x69249, x69250;
  wire x69251, x69252, x69253, x69254, x69255, x69256, x69257, x69258;
  wire x69259, x69260, x69261, x69262, x69263, x69264, x69265, x69266;
  wire x69267, x69268, x69269, x69270, x69271, x69272, x69273, x69274;
  wire x69275, x69276, x69277, x69278, x69279, x69280, x69281, x69282;
  wire x69283, x69284, x69285, x69286, x69287, x69288, x69289, x69290;
  wire x69291, x69292, x69293, x69294, x69295, x69296, x69297, x69298;
  wire x69299, x69300, x69301, x69302, x69303, x69304, x69305, x69306;
  wire x69307, x69308, x69309, x69310, x69311, x69312, x69313, x69314;
  wire x69315, x69316, x69317, x69318, x69319, x69320, x69321, x69322;
  wire x69323, x69324, x69325, x69326, x69327, x69328, x69329, x69330;
  wire x69331, x69332, x69333, x69334, x69335, x69336, x69337, x69338;
  wire x69339, x69340, x69341, x69342, x69343, x69344, x69345, x69346;
  wire x69347, x69348, x69349, x69350, x69351, x69352, x69353, x69354;
  wire x69355, x69356, x69357, x69358, x69359, x69360, x69361, x69362;
  wire x69363, x69364, x69365, x69366, x69367, x69368, x69369, x69370;
  wire x69371, x69372, x69373, x69374, x69375, x69376, x69377, x69378;
  wire x69379, x69380, x69381, x69382, x69383, x69384, x69385, x69386;
  wire x69387, x69388, x69389, x69390, x69391, x69392, x69393, x69394;
  wire x69395, x69396, x69397, x69398, x69399, x69400, x69401, x69402;
  wire x69403, x69404, x69405, x69406, x69407, x69408, x69409, x69410;
  wire x69411, x69412, x69413, x69414, x69415, x69416, x69417, x69418;
  wire x69419, x69420, x69421, x69422, x69423, x69424, x69425, x69426;
  wire x69427, x69428, x69429, x69430, x69431, x69432, x69433, x69434;
  wire x69435, x69436, x69437, x69438, x69439, x69440, x69441, x69442;
  wire x69443, x69444, x69445, x69446, x69447, x69448, x69449, x69450;
  wire x69451, x69452, x69453, x69454, x69455, x69456, x69457, x69458;
  wire x69459, x69460, x69461, x69462, x69463, x69464, x69465, x69466;
  wire x69467, x69468, x69469, x69470, x69471, x69472, x69473, x69474;
  wire x69475, x69476, x69477, x69478, x69479, x69480, x69481, x69482;
  wire x69483, x69484, x69485, x69486, x69487, x69488, x69489, x69490;
  wire x69491, x69492, x69493, x69494, x69495, x69496, x69497, x69498;
  wire x69499, x69500, x69501, x69502, x69503, x69504, x69505, x69506;
  wire x69507, x69508, x69509, x69510, x69511, x69512, x69513, x69514;
  wire x69515, x69516, x69517, x69518, x69519, x69520, x69521, x69522;
  wire x69523, x69524, x69525, x69526, x69527, x69528, x69529, x69530;
  wire x69531, x69532, x69533, x69534, x69535, x69536, x69537, x69538;
  wire x69539, x69540, x69541, x69542, x69543, x69544, x69545, x69546;
  wire x69547, x69548, x69549, x69550, x69551, x69552, x69553, x69554;
  wire x69555, x69556, x69557, x69558, x69559, x69560, x69561, x69562;
  wire x69563, x69564, x69565, x69566, x69567, x69568, x69569, x69570;
  wire x69571, x69572, x69573, x69574, x69575, x69576, x69577, x69578;
  wire x69579, x69580, x69581, x69582, x69583, x69584, x69585, x69586;
  wire x69587, x69588, x69589, x69590, x69591, x69592, x69593, x69594;
  wire x69595, x69596, x69597, x69598, x69599, x69600, x69601, x69602;
  wire x69603, x69604, x69605, x69606, x69607, x69608, x69609, x69610;
  wire x69611, x69612, x69613, x69614, x69615, x69616, x69617, x69618;
  wire x69619, x69620, x69621, x69622, x69623, x69624, x69625, x69626;
  wire x69627, x69628, x69629, x69630, x69631, x69632, x69633, x69634;
  wire x69635, x69636, x69637, x69638, x69639, x69640, x69641, x69642;
  wire x69643, x69644, x69645, x69646, x69647, x69648, x69649, x69650;
  wire x69651, x69652, x69653, x69654, x69655, x69656, x69657, x69658;
  wire x69659, x69660, x69661, x69662, x69663, x69664, x69665, x69666;
  wire x69667, x69668, x69669, x69670, x69671, x69672, x69673, x69674;
  wire x69675, x69676, x69677, x69678, x69679, x69680, x69681, x69682;
  wire x69683, x69684, x69685, x69686, x69687, x69688, x69689, x69690;
  wire x69691, x69692, x69693, x69694, x69695, x69696, x69697, x69698;
  wire x69699, x69700, x69701, x69702, x69703, x69704, x69705, x69706;
  wire x69707, x69708, x69709, x69710, x69711, x69712, x69713, x69714;
  wire x69715, x69716, x69717, x69718, x69719, x69720, x69721, x69722;
  wire x69723, x69724, x69725, x69726, x69727, x69728, x69729, x69730;
  wire x69731, x69732, x69733, x69734, x69735, x69736, x69737, x69738;
  wire x69739, x69740, x69741, x69742, x69743, x69744, x69745, x69746;
  wire x69747, x69748, x69749, x69750, x69751, x69752, x69753, x69754;
  wire x69755, x69756, x69757, x69758, x69759, x69760, x69761, x69762;
  wire x69763, x69764, x69765, x69766, x69767, x69768, x69769, x69770;
  wire x69771, x69772, x69773, x69774, x69775, x69776, x69777, x69778;
  wire x69779, x69780, x69781, x69782, x69783, x69784, x69785, x69786;
  wire x69787, x69788, x69789, x69790, x69791, x69792, x69793, x69794;
  wire x69795, x69796, x69797, x69798, x69799, x69800, x69801, x69802;
  wire x69803, x69804, x69805, x69806, x69807, x69808, x69809, x69810;
  wire x69811, x69812, x69813, x69814, x69815, x69816, x69817, x69818;
  wire x69819, x69820, x69821, x69822, x69823, x69824, x69825, x69826;
  wire x69827, x69828, x69829, x69830, x69831, x69832, x69833, x69834;
  wire x69835, x69836, x69837, x69838, x69839, x69840, x69841, x69842;
  wire x69843, x69844, x69845, x69846, x69847, x69848, x69849, x69850;
  wire x69851, x69852, x69853, x69854, x69855, x69856, x69857, x69858;
  wire x69859, x69860, x69861, x69862, x69863, x69864, x69865, x69866;
  wire x69867, x69868, x69869, x69870, x69871, x69872, x69873, x69874;
  wire x69875, x69876, x69877, x69878, x69879, x69880, x69881, x69882;
  wire x69883, x69884, x69885, x69886, x69887, x69888, x69889, x69890;
  wire x69891, x69892, x69893, x69894, x69895, x69896, x69897, x69898;
  wire x69899, x69900, x69901, x69902, x69903, x69904, x69905, x69906;
  wire x69907, x69908, x69909, x69910, x69911, x69912, x69913, x69914;
  wire x69915, x69916, x69917, x69918, x69919, x69920, x69921, x69922;
  wire x69923, x69924, x69925, x69926, x69927, x69928, x69929, x69930;
  wire x69931, x69932, x69933, x69934, x69935, x69936, x69937, x69938;
  wire x69939, x69940, x69941, x69942, x69943, x69944, x69945, x69946;
  wire x69947, x69948, x69949, x69950, x69951, x69952, x69953, x69954;
  wire x69955, x69956, x69957, x69958, x69959, x69960, x69961, x69962;
  wire x69963, x69964, x69965, x69966, x69967, x69968, x69969, x69970;
  wire x69971, x69972, x69973, x69974, x69975, x69976, x69977, x69978;
  wire x69979, x69980, x69981, x69982, x69983, x69984, x69985, x69986;
  wire x69987, x69988, x69989, x69990, x69991, x69992, x69993, x69994;
  wire x69995, x69996, x69997, x69998, x69999, x70000, x70001, x70002;
  wire x70003, x70004, x70005, x70006, x70007, x70008, x70009, x70010;
  wire x70011, x70012, x70013, x70014, x70015, x70016, x70017, x70018;
  wire x70019, x70020, x70021, x70022, x70023, x70024, x70025, x70026;
  wire x70027, x70028, x70029, x70030, x70031, x70032, x70033, x70034;
  wire x70035, x70036, x70037, x70038, x70039, x70040, x70041, x70042;
  wire x70043, x70044, x70045, x70046, x70047, x70048, x70049, x70050;
  wire x70051, x70052, x70053, x70054, x70055, x70056, x70057, x70058;
  wire x70059, x70060, x70061, x70062, x70063, x70064, x70065, x70066;
  wire x70067, x70068, x70069, x70070, x70071, x70072, x70073, x70074;
  wire x70075, x70076, x70077, x70078, x70079, x70080, x70081, x70082;
  wire x70083, x70084, x70085, x70086, x70087, x70088, x70089, x70090;
  wire x70091, x70092, x70093, x70094, x70095, x70096, x70097, x70098;
  wire x70099, x70100, x70101, x70102, x70103, x70104, x70105, x70106;
  wire x70107, x70108, x70109, x70110, x70111, x70112, x70113, x70114;
  wire x70115, x70116, x70117, x70118, x70119, x70120, x70121, x70122;
  wire x70123, x70124, x70125, x70126, x70127, x70128, x70129, x70130;
  wire x70131, x70132, x70133, x70134, x70135, x70136, x70137, x70138;
  wire x70139, x70140, x70141, x70142, x70143, x70144, x70145, x70146;
  wire x70147, x70148, x70149, x70150, x70151, x70152, x70153, x70154;
  wire x70155, x70156, x70157, x70158, x70159, x70160, x70161, x70162;
  wire x70163, x70164, x70165, x70166, x70167, x70168, x70169, x70170;
  wire x70171, x70172, x70173, x70174, x70175, x70176, x70177, x70178;
  wire x70179, x70180, x70181, x70182, x70183, x70184, x70185, x70186;
  wire x70187, x70188, x70189, x70190, x70191, x70192, x70193, x70194;
  wire x70195, x70196, x70197, x70198, x70199, x70200, x70201, x70202;
  wire x70203, x70204, x70205, x70206, x70207, x70208, x70209, x70210;
  wire x70211, x70212, x70213, x70214, x70215, x70216, x70217, x70218;
  wire x70219, x70220, x70221, x70222, x70223, x70224, x70225, x70226;
  wire x70227, x70228, x70229, x70230, x70231, x70232, x70233, x70234;
  wire x70235, x70236, x70237, x70238, x70239, x70240, x70241, x70242;
  wire x70243, x70244, x70245, x70246, x70247, x70248, x70249, x70250;
  wire x70251, x70252, x70253, x70254, x70255, x70256, x70257, x70258;
  wire x70259, x70260, x70261, x70262, x70263, x70264, x70265, x70266;
  wire x70267, x70268, x70269, x70270, x70271, x70272, x70273, x70274;
  wire x70275, x70276, x70277, x70278, x70279, x70280, x70281, x70282;
  wire x70283, x70284, x70285, x70286, x70287, x70288, x70289, x70290;
  wire x70291, x70292, x70293, x70294, x70295, x70296, x70297, x70298;
  wire x70299, x70300, x70301, x70302, x70303, x70304, x70305, x70306;
  wire x70307, x70308, x70309, x70310, x70311, x70312, x70313, x70314;
  wire x70315, x70316, x70317, x70318, x70319, x70320, x70321, x70322;
  wire x70323, x70324, x70325, x70326, x70327, x70328, x70329, x70330;
  wire x70331, x70332, x70333, x70334, x70335, x70336, x70337, x70338;
  wire x70339, x70340, x70341, x70342, x70343, x70344, x70345, x70346;
  wire x70347, x70348, x70349, x70350, x70351, x70352, x70353, x70354;
  wire x70355, x70356, x70357, x70358, x70359, x70360, x70361, x70362;
  wire x70363, x70364, x70365, x70366, x70367, x70368, x70369, x70370;
  wire x70371, x70372, x70373, x70374, x70375, x70376, x70377, x70378;
  wire x70379, x70380, x70381, x70382, x70383, x70384, x70385, x70386;
  wire x70387, x70388, x70389, x70390, x70391, x70392, x70393, x70394;
  wire x70395, x70396, x70397, x70398, x70399, x70400, x70401, x70402;
  wire x70403, x70404, x70405, x70406, x70407, x70408, x70409, x70410;
  wire x70411, x70412, x70413, x70414, x70415, x70416, x70417, x70418;
  wire x70419, x70420, x70421, x70422, x70423, x70424, x70425, x70426;
  wire x70427, x70428, x70429, x70430, x70431, x70432, x70433, x70434;
  wire x70435, x70436, x70437, x70438, x70439, x70440, x70441, x70442;
  wire x70443, x70444, x70445, x70446, x70447, x70448, x70449, x70450;
  wire x70451, x70452, x70453, x70454, x70455, x70456, x70457, x70458;
  wire x70459, x70460, x70461, x70462, x70463, x70464, x70465, x70466;
  wire x70467, x70468, x70469, x70470, x70471, x70472, x70473, x70474;
  wire x70475, x70476, x70477, x70478, x70479, x70480, x70481, x70482;
  wire x70483, x70484, x70485, x70486, x70487, x70488, x70489, x70490;
  wire x70491, x70492, x70493, x70494, x70495, x70496, x70497, x70498;
  wire x70499, x70500, x70501, x70502, x70503, x70504, x70505, x70506;
  wire x70507, x70508, x70509, x70510, x70511, x70512, x70513, x70514;
  wire x70515, x70516, x70517, x70518, x70519, x70520, x70521, x70522;
  wire x70523, x70524, x70525, x70526, x70527, x70528, x70529, x70530;
  wire x70531, x70532, x70533, x70534, x70535, x70536, x70537, x70538;
  wire x70539, x70540, x70541, x70542, x70543, x70544, x70545, x70546;
  wire x70547, x70548, x70549, x70550, x70551, x70552, x70553, x70554;
  wire x70555, x70556, x70557, x70558, x70559, x70560, x70561, x70562;
  wire x70563, x70564, x70565, x70566, x70567, x70568, x70569, x70570;
  wire x70571, x70572, x70573, x70574, x70575, x70576, x70577, x70578;
  wire x70579, x70580, x70581, x70582, x70583, x70584, x70585, x70586;
  wire x70587, x70588, x70589, x70590, x70591, x70592, x70593, x70594;
  wire x70595, x70596, x70597, x70598, x70599, x70600, x70601, x70602;
  wire x70603, x70604, x70605, x70606, x70607, x70608, x70609, x70610;
  wire x70611, x70612, x70613, x70614, x70615, x70616, x70617, x70618;
  wire x70619, x70620, x70621, x70622, x70623, x70624, x70625, x70626;
  wire x70627, x70628, x70629, x70630, x70631, x70632, x70633, x70634;
  wire x70635, x70636, x70637, x70638, x70639, x70640, x70641, x70642;
  wire x70643, x70644, x70645, x70646, x70647, x70648, x70649, x70650;
  wire x70651, x70652, x70653, x70654, x70655, x70656, x70657, x70658;
  wire x70659, x70660, x70661, x70662, x70663, x70664, x70665, x70666;
  wire x70667, x70668, x70669, x70670, x70671, x70672, x70673, x70674;
  wire x70675, x70676, x70677, x70678, x70679, x70680, x70681, x70682;
  wire x70683, x70684, x70685, x70686, x70687, x70688, x70689, x70690;
  wire x70691, x70692, x70693, x70694, x70695, x70696, x70697, x70698;
  wire x70699, x70700, x70701, x70702, x70703, x70704, x70705, x70706;
  wire x70707, x70708, x70709, x70710, x70711, x70712, x70713, x70714;
  wire x70715, x70716, x70717, x70718, x70719, x70720, x70721, x70722;
  wire x70723, x70724, x70725, x70726, x70727, x70728, x70729, x70730;
  wire x70731, x70732, x70733, x70734, x70735, x70736, x70737, x70738;
  wire x70739, x70740, x70741, x70742, x70743, x70744, x70745, x70746;
  wire x70747, x70748, x70749, x70750, x70751, x70752, x70753, x70754;
  wire x70755, x70756, x70757, x70758, x70759, x70760, x70761, x70762;
  wire x70763, x70764, x70765, x70766, x70767, x70768, x70769, x70770;
  wire x70771, x70772, x70773, x70774, x70775, x70776, x70777, x70778;
  wire x70779, x70780, x70781, x70782, x70783, x70784, x70785, x70786;
  wire x70787, x70788, x70789, x70790, x70791, x70792, x70793, x70794;
  wire x70795, x70796, x70797, x70798, x70799, x70800, x70801, x70802;
  wire x70803, x70804, x70805, x70806, x70807, x70808, x70809, x70810;
  wire x70811, x70812, x70813, x70814, x70815, x70816, x70817, x70818;
  wire x70819, x70820, x70821, x70822, x70823, x70824, x70825, x70826;
  wire x70827, x70828, x70829, x70830, x70831, x70832, x70833, x70834;
  wire x70835, x70836, x70837, x70838, x70839, x70840, x70841, x70842;
  wire x70843, x70844, x70845, x70846, x70847, x70848, x70849, x70850;
  wire x70851, x70852, x70853, x70854, x70855, x70856, x70857, x70858;
  wire x70859, x70860, x70861, x70862, x70863, x70864, x70865, x70866;
  wire x70867, x70868, x70869, x70870, x70871, x70872, x70873, x70874;
  wire x70875, x70876, x70877, x70878, x70879, x70880, x70881, x70882;
  wire x70883, x70884, x70885, x70886, x70887, x70888, x70889, x70890;
  wire x70891, x70892, x70893, x70894, x70895, x70896, x70897, x70898;
  wire x70899, x70900, x70901, x70902, x70903, x70904, x70905, x70906;
  wire x70907, x70908, x70909, x70910, x70911, x70912, x70913, x70914;
  wire x70915, x70916, x70917, x70918, x70919, x70920, x70921, x70922;
  wire x70923, x70924, x70925, x70926, x70927, x70928, x70929, x70930;
  wire x70931, x70932, x70933, x70934, x70935, x70936, x70937, x70938;
  wire x70939, x70940, x70941, x70942, x70943, x70944, x70945, x70946;
  wire x70947, x70948, x70949, x70950, x70951, x70952, x70953, x70954;
  wire x70955, x70956, x70957, x70958, x70959, x70960, x70961, x70962;
  wire x70963, x70964, x70965, x70966, x70967, x70968, x70969, x70970;
  wire x70971, x70972, x70973, x70974, x70975, x70976, x70977, x70978;
  wire x70979, x70980, x70981, x70982, x70983, x70984, x70985, x70986;
  wire x70987, x70988, x70989, x70990, x70991, x70992, x70993, x70994;
  wire x70995, x70996, x70997, x70998, x70999, x71000, x71001, x71002;
  wire x71003, x71004, x71005, x71006, x71007, x71008, x71009, x71010;
  wire x71011, x71012, x71013, x71014, x71015, x71016, x71017, x71018;
  wire x71019, x71020, x71021, x71022, x71023, x71024, x71025, x71026;
  wire x71029, x71030, x71031, x71034, x71035, x71036, x71039, x71040;
  wire x71041, x71044, x71045, x71046, x71049, x71050, x71051, x71054;
  wire x71055, x71056, x71058, x71060, x71062, x71064, x71066, x71068;
  wire x71070, x71072, x71074, x71076, x71079, x71080, x71081, x71084;
  wire x71085, x71086, x71089, x71090, x71091, x71094, x71095, x71096;
  wire x71099, x71100, x71101, x71104, x71105, x71106, x71108, x71110;
  wire x71112, x71114, x71116, x71118, x71120, x71122, x71124, x71128;
  wire x71129, x71130, x71131, x71134, x71137, x71140, x71141, x71142;
  wire x71143, x71144, x71145, x71146, x71148, x71149, x71150, x71151;
  wire x71153, x71154, x71155, x71156, x71158, x71159, x71160, x71161;
  wire x71163, x71164, x71165, x71166, x71168, x71169, x71170, x71171;
  wire x71173, x71174, x71175, x71176, x71178, x71179, x71180, x71181;
  wire x71183, x71184, x71186, x71187, x71189, x71190, x71192, x71193;
  wire x71195, x71196, x71198, x71199, x71200, x71201, x71203, x71204;
  wire x71206, x71207, x71208, x71209, x71211, x71212, x71213, x71214;
  wire x71216, x71217, x71218, x71219, x71221, x71222, x71223, x71224;
  wire x71226, x71227, x71228, x71229, x71231, x71232, x71233, x71234;
  wire x71236, x71237, x71238, x71239, x71241, x71242, x71243, x71244;
  wire x71246, x71247, x71248, x71249, x71251, x71252, x71253, x71254;
  wire x71256, x71257, x71258, x71259, x71261, x71262, x71263, x71264;
  wire x71266, x71267, x71268, x71269, x71271, x71272, x71273, x71274;
  wire x71276, x71278, x71280, x71281, x71282, x71283, x71285, x71286;
  wire x71287, x71288, x71290, x71291, x71292, x71293, x71295, x71296;
  wire x71297, x71298, x71300, x71301, x71302, x71303, x71305, x71306;
  wire x71307, x71308, x71310, x71311, x71312, x71313, x71315, x71316;
  wire x71317, x71318, x71320, x71321, x71322, x71323, x71325, x71326;
  wire x71327, x71328, x71330, x71331, x71332, x71333, x71335, x71336;
  wire x71337, x71338, x71340, x71341, x71342, x71343, x71345, x71346;
  wire x71347, x71348, x71350, x71351, x71352, x71353, x71355, x71356;
  wire x71357, x71358, x71360, x71361, x71362, x71363, x71365, x71366;
  wire x71367, x71368, x71370, x71371, x71372, x71373, x71375, x71376;
  wire x71377, x71378, x71380, x71381, x71382, x71383, x71385, x71386;
  wire x71387, x71388, x71390, x71391, x71392, x71393, x71395, x71396;
  wire x71397, x71398, x71400, x71401, x71402, x71403, x71405, x71406;
  wire x71407, x71408, x71410, x71411, x71412, x71413, x71415, x71416;
  wire x71417, x71418, x71420, x71421, x71422, x71423, x71425, x71426;
  wire x71427, x71428, x71430, x71431, x71432, x71433, x71435, x71436;
  wire x71437, x71438, x71440, x71441, x71442, x71443, x71445, x71446;
  wire x71447, x71448, x71450, x71451, x71452, x71453, x71455, x71456;
  wire x71457, x71458, x71460, x71461, x71462, x71463, x71465, x71466;
  wire x71467, x71468, x71470, x71471, x71472, x71473, x71475, x71476;
  wire x71477, x71478, x71480, x71481, x71483, x71484, x71486, x71487;
  wire x71488, x71489, x71491, x71492, x71493, x71494, x71496, x71497;
  wire x71498, x71499, x71501, x71502, x71503, x71504, x71506, x71507;
  wire x71508, x71509, x71511, x71512, x71513, x71514, x71516, x71517;
  wire x71518, x71519, x71521, x71522, x71523, x71524, x71526, x71527;
  wire x71528, x71529, x71531, x71532, x71533, x71534, x71536, x71537;
  wire x71538, x71539, x71541, x71542, x71543, x71544, x71546, x71547;
  wire x71548, x71549, x71551, x71552, x71553, x71554, x71556, x71557;
  wire x71558, x71559, x71561, x71562, x71563, x71564, x71566, x71567;
  wire x71568, x71569, x71571, x71572, x71573, x71574, x71576, x71577;
  wire x71578, x71579, x71581, x71582, x71583, x71584, x71586, x71587;
  wire x71588, x71589, x71591, x71592, x71593, x71594, x71596, x71597;
  wire x71598, x71599, x71601, x71602, x71603, x71604, x71606, x71607;
  wire x71608, x71609, x71611, x71612, x71613, x71614, x71616, x71617;
  wire x71618, x71619, x71621, x71622, x71623, x71624, x71626, x71627;
  wire x71628, x71629, x71631, x71632, x71633, x71634, x71636, x71637;
  wire x71638, x71639, x71640, x71641, x71643, x71644, x71645, x71646;
  wire x71648, x71649, x71650, x71651, x71653, x71654, x71655, x71656;
  wire x71658, x71659, x71660, x71661, x71663, x71664, x71665, x71666;
  wire x71668, x71669, x71670, x71671, x71673, x71674, x71675, x71676;
  wire x71678, x71679, x71680, x71681, x71683, x71684, x71685, x71686;
  wire x71688, x71689, x71690, x71691, x71693, x71694, x71695, x71696;
  wire x71698, x71699, x71700, x71701, x71703, x71704, x71705, x71706;
  wire x71708, x71709, x71710, x71711, x71713, x71714, x71715, x71716;
  wire x71718, x71719, x71720, x71721, x71723, x71724, x71725, x71726;
  wire x71728, x71729, x71730, x71731, x71733, x71734, x71735, x71736;
  wire x71738, x71739, x71740, x71741, x71743, x71744, x71745, x71746;
  wire x71748, x71749, x71750, x71751, x71753, x71754, x71755, x71756;
  wire x71758, x71759, x71760, x71761, x71763, x71764, x71765, x71766;
  wire x71768, x71769, x71770, x71771, x71773, x71774, x71775, x71776;
  wire x71778, x71779, x71780, x71781, x71783, x71784, x71785, x71786;
  wire x71788, x71789, x71790, x71791, x71793, x71794, x71795, x71796;
  wire x71798, x71799, x71800, x71801, x71803, x71804, x71805, x71806;
  wire x71808, x71809, x71810, x71811, x71813, x71814, x71815, x71816;
  wire x71818, x71819, x71820, x71821, x71823, x71824, x71825, x71826;
  wire x71828, x71829, x71830, x71831, x71833, x71834, x71835, x71836;
  wire x71838, x71839, x71840, x71841, x71843, x71844, x71845, x71846;
  wire x71848, x71849, x71850, x71851, x71853, x71854, x71855, x71856;
  wire x71858, x71859, x71860, x71861, x71863, x71864, x71865, x71866;
  wire x71868, x71869, x71870, x71871, x71873, x71874, x71875, x71876;
  wire x71878, x71879, x71880, x71881, x71883, x71884, x71885, x71886;
  wire x71888, x71889, x71890, x71891, x71893, x71894, x71895, x71896;
  wire x71898, x71899, x71900, x71901, x71903, x71904, x71905, x71906;
  wire x71908, x71909, x71911, x71912, x71914, x71915, x71917, x71918;
  wire x71920, x71921, x71923, x71924, x71926, x71927, x71929, x71930;
  wire x71932, x71933, x71935, x71936, x71938, x71939, x71940, x71941;
  wire x71943, x71944, x71945, x71946, x71948, x71949, x71950, x71951;
  wire x71953, x71954, x71955, x71956, x71958, x71959, x71960, x71961;
  wire x71963, x71964, x71965, x71966, x71968, x71969, x71970, x71971;
  wire x71973, x71974, x71975, x71976, x71978, x71979, x71980, x71981;
  wire x71983, x71984, x71985, x71986, x71988, x71989, x71990, x71991;
  wire x71993, x71994, x71995, x71996, x71998, x71999, x72000, x72001;
  wire x72003, x72004, x72005, x72006, x72008, x72009, x72010, x72011;
  wire x72013, x72014, x72015, x72016, x72018, x72019, x72020, x72021;
  wire x72023, x72024, x72025, x72026, x72028, x72029, x72030, x72031;
  wire x72033, x72034, x72035, x72036, x72038, x72039, x72040, x72041;
  wire x72043, x72044, x72045, x72046, x72048, x72049, x72050, x72051;
  wire x72053, x72054, x72055, x72056, x72058, x72059, x72060, x72061;
  wire x72063, x72064, x72065, x72066, x72068, x72069, x72070, x72071;
  wire x72073, x72074, x72075, x72076, x72078, x72079, x72080, x72081;
  wire x72083, x72084, x72085, x72086, x72088, x72089, x72090, x72091;
  wire x72093, x72094, x72095, x72096, x72098, x72099, x72100, x72101;
  wire x72103, x72104, x72105, x72106, x72108, x72109, x72110, x72111;
  wire x72113, x72114, x72115, x72116, x72118, x72119, x72120, x72121;
  wire x72123, x72124, x72125, x72126, x72128, x72129, x72130, x72131;
  wire x72133, x72134, x72135, x72136, x72138, x72139, x72140, x72141;
  wire x72143, x72144, x72145, x72146, x72148, x72149, x72150, x72151;
  wire x72153, x72154, x72155, x72156, x72158, x72159, x72160, x72161;
  wire x72163, x72164, x72165, x72166, x72168, x72169, x72170, x72171;
  wire x72173, x72174, x72175, x72176, x72178, x72179, x72180, x72181;
  wire x72183, x72184, x72185, x72186, x72188, x72189, x72190, x72191;
  wire x72193, x72194, x72195, x72196, x72198, x72199, x72200, x72201;
  wire x72203, x72204, x72205, x72206, x72208, x72209, x72210, x72211;
  wire x72213, x72214, x72215, x72216, x72218, x72219, x72220, x72221;
  wire x72223, x72224, x72225, x72226, x72228, x72229, x72230, x72231;
  wire x72233, x72234, x72235, x72236, x72238, x72239, x72240, x72241;
  wire x72243, x72244, x72245, x72246, x72248, x72249, x72250, x72251;
  wire x72253, x72254, x72255, x72256, x72258, x72259, x72260, x72261;
  wire x72263, x72264, x72265, x72266, x72268, x72269, x72270, x72271;
  wire x72273, x72274, x72275, x72276, x72278, x72279, x72280, x72281;
  wire x72283, x72284, x72285, x72286, x72288, x72289, x72290, x72291;
  wire x72293, x72294, x72295, x72296, x72298, x72299, x72300, x72301;
  wire x72303, x72304, x72305, x72306, x72308, x72309, x72310, x72311;
  wire x72313, x72314, x72315, x72316, x72318, x72319, x72320, x72321;
  wire x72323, x72324, x72325, x72326, x72328, x72329, x72330, x72331;
  wire x72333, x72334, x72335, x72336, x72338, x72339, x72340, x72341;
  wire x72343, x72344, x72345, x72346, x72348, x72349, x72350, x72351;
  wire x72353, x72354, x72355, x72356, x72358, x72359, x72360, x72361;
  wire x72363, x72364, x72365, x72366, x72368, x72369, x72370, x72371;
  wire x72373, x72374, x72375, x72376, x72378, x72379, x72380, x72381;
  wire x72383, x72384, x72385, x72386, x72388, x72389, x72390, x72391;
  wire x72393, x72394, x72395, x72396, x72398, x72399, x72400, x72401;
  wire x72403, x72404, x72405, x72406, x72408, x72409, x72410, x72411;
  wire x72413, x72414, x72415, x72416, x72418, x72419, x72420, x72421;
  wire x72423, x72424, x72425, x72426, x72428, x72429, x72430, x72431;
  wire x72433, x72434, x72435, x72436, x72438, x72439, x72440, x72441;
  wire x72443, x72444, x72445, x72446, x72448, x72449, x72450, x72451;
  wire x72453, x72454, x72455, x72456, x72458, x72459, x72460, x72461;
  wire x72463, x72464, x72465, x72466, x72468, x72469, x72470, x72471;
  wire x72473, x72474, x72475, x72476, x72478, x72479, x72480, x72481;
  wire x72483, x72484, x72485, x72486, x72488, x72489, x72490, x72491;
  wire x72493, x72494, x72495, x72496, x72498, x72499, x72500, x72501;
  wire x72503, x72504, x72505, x72506, x72508, x72509, x72510, x72511;
  wire x72513, x72514, x72515, x72516, x72518, x72519, x72520, x72521;
  wire x72523, x72524, x72525, x72526, x72528, x72529, x72530, x72531;
  wire x72533, x72534, x72535, x72536, x72538, x72539, x72540, x72541;
  wire x72543, x72544, x72545, x72546, x72548, x72549, x72550, x72551;
  wire x72553, x72554, x72555, x72556, x72558, x72559, x72560, x72561;
  wire x72563, x72564, x72565, x72566, x72568, x72569, x72570, x72571;
  wire x72573, x72574, x72575, x72576, x72578, x72579, x72580, x72581;
  wire x72583, x72584, x72585, x72586, x72588, x72589, x72590, x72591;
  wire x72593, x72594, x72595, x72596, x72598, x72599, x72600, x72601;
  wire x72603, x72604, x72605, x72606, x72608, x72609, x72610, x72611;
  wire x72613, x72614, x72615, x72616, x72618, x72619, x72620, x72621;
  wire x72623, x72624, x72625, x72626, x72628, x72629, x72630, x72631;
  wire x72633, x72634, x72635, x72636, x72638, x72639, x72640, x72641;
  wire x72643, x72644, x72645, x72646, x72648, x72649, x72650, x72651;
  wire x72653, x72654, x72655, x72656, x72658, x72659, x72660, x72661;
  wire x72663, x72664, x72665, x72666, x72668, x72669, x72670, x72671;
  wire x72673, x72674, x72675, x72676, x72678, x72679, x72680, x72681;
  wire x72683, x72684, x72685, x72686, x72688, x72689, x72690, x72691;
  wire x72693, x72694, x72695, x72696, x72698, x72699, x72700, x72701;
  wire x72703, x72704, x72705, x72706, x72708, x72709, x72710, x72711;
  wire x72713, x72714, x72715, x72716, x72718, x72719, x72720, x72721;
  wire x72723, x72724, x72725, x72726, x72728, x72729, x72730, x72731;
  wire x72733, x72734, x72735, x72736, x72738, x72739, x72740, x72741;
  wire x72743, x72744, x72745, x72746, x72748, x72749, x72750, x72751;
  wire x72753, x72754, x72755, x72756, x72758, x72759, x72760, x72761;
  wire x72763, x72764, x72765, x72766, x72768, x72769, x72770, x72771;
  wire x72773, x72774, x72775, x72776, x72778, x72779, x72780, x72781;
  wire x72783, x72784, x72785, x72786, x72788, x72789, x72790, x72791;
  wire x72793, x72794, x72795, x72796, x72798, x72799, x72800, x72801;
  wire x72803, x72804, x72805, x72806, x72808, x72809, x72810, x72811;
  wire x72813, x72814, x72815, x72816, x72818, x72819, x72820, x72821;
  wire x72823, x72824, x72825, x72826, x72828, x72829, x72830, x72831;
  wire x72833, x72834, x72835, x72836, x72838, x72839, x72840, x72841;
  wire x72843, x72844, x72845, x72846, x72848, x72849, x72850, x72851;
  wire x72853, x72854, x72855, x72856, x72858, x72859, x72860, x72861;
  wire x72863, x72864, x72865, x72866, x72868, x72869, x72870, x72871;
  wire x72873, x72874, x72875, x72876, x72878, x72879, x72880, x72881;
  wire x72883, x72884, x72885, x72886, x72888, x72889, x72890, x72891;
  wire x72893, x72894, x72895, x72896, x72898, x72899, x72900, x72901;
  wire x72903, x72904, x72905, x72906, x72908, x72909, x72910, x72911;
  wire x72913, x72914, x72915, x72916, x72918, x72919, x72920, x72921;
  wire x72923, x72924, x72925, x72926, x72928, x72929, x72930, x72931;
  wire x72933, x72934, x72935, x72936, x72938, x72939, x72940, x72941;
  wire x72943, x72944, x72945, x72946, x72948, x72949, x72950, x72951;
  wire x72953, x72954, x72955, x72956, x72958, x72959, x72960, x72961;
  wire x72963, x72964, x72965, x72966, x72968, x72969, x72970, x72971;
  wire x72973, x72974, x72975, x72976, x72978, x72979, x72980, x72981;
  wire x72983, x72984, x72985, x72986, x72988, x72989, x72990, x72991;
  wire x72993, x72994, x72995, x72996, x72998, x72999, x73000, x73001;
  wire x73003, x73004, x73005, x73006, x73008, x73009, x73010, x73011;
  wire x73013, x73014, x73015, x73016, x73018, x73019, x73020, x73021;
  wire x73023, x73024, x73025, x73026, x73028, x73029, x73030, x73031;
  wire x73033, x73034, x73035, x73036, x73038, x73039, x73040, x73041;
  wire x73043, x73044, x73045, x73046, x73048, x73049, x73050, x73051;
  wire x73053, x73054, x73055, x73056, x73058, x73059, x73060, x73061;
  wire x73063, x73064, x73065, x73066, x73068, x73069, x73070, x73071;
  wire x73073, x73074, x73075, x73076, x73078, x73079, x73080, x73081;
  wire x73083, x73084, x73085, x73086, x73088, x73089, x73090, x73091;
  wire x73093, x73094, x73095, x73096, x73098, x73099, x73100, x73101;
  wire x73103, x73104, x73105, x73106, x73108, x73109, x73110, x73111;
  wire x73113, x73114, x73115, x73116, x73118, x73119, x73120, x73121;
  wire x73123, x73124, x73125, x73126, x73128, x73129, x73130, x73131;
  wire x73133, x73134, x73135, x73136, x73138, x73139, x73140, x73141;
  wire x73143, x73144, x73145, x73146, x73148, x73149, x73150, x73151;
  wire x73153, x73154, x73155, x73156, x73158, x73159, x73160, x73161;
  wire x73163, x73164, x73165, x73166, x73168, x73169, x73170, x73171;
  wire x73173, x73174, x73175, x73176, x73178, x73179, x73180, x73181;
  wire x73183, x73184, x73185, x73186, x73188, x73189, x73190, x73191;
  wire x73193, x73194, x73195, x73196, x73198, x73199, x73200, x73201;
  wire x73203, x73204, x73205, x73206, x73208, x73209, x73210, x73211;
  wire x73213, x73214, x73215, x73216, x73218, x73219, x73220, x73221;
  wire x73223, x73224, x73225, x73226, x73228, x73229, x73230, x73231;
  wire x73233, x73234, x73235, x73236, x73238, x73239, x73240, x73241;
  wire x73243, x73244, x73245, x73246, x73248, x73249, x73250, x73251;
  wire x73253, x73254, x73255, x73256, x73258, x73259, x73260, x73261;
  wire x73263, x73264, x73265, x73266, x73268, x73269, x73270, x73271;
  wire x73273, x73274, x73275, x73276, x73278, x73279, x73280, x73281;
  wire x73283, x73284, x73285, x73286, x73288, x73289, x73290, x73291;
  wire x73293, x73294, x73295, x73296, x73298, x73299, x73300, x73301;
  wire x73303, x73304, x73305, x73306, x73308, x73309, x73310, x73311;
  wire x73313, x73314, x73315, x73316, x73318, x73319, x73320, x73321;
  wire x73323, x73324, x73325, x73326, x73328, x73329, x73330, x73331;
  wire x73333, x73334, x73335, x73336, x73338, x73339, x73340, x73341;
  wire x73343, x73344, x73345, x73346, x73348, x73349, x73350, x73351;
  wire x73353, x73354, x73355, x73356, x73358, x73359, x73360, x73361;
  wire x73363, x73364, x73365, x73366, x73368, x73369, x73370, x73371;
  wire x73373, x73374, x73375, x73376, x73378, x73379, x73380, x73381;
  wire x73383, x73384, x73385, x73386, x73388, x73389, x73390, x73391;
  wire x73393, x73394, x73395, x73396, x73398, x73399, x73400, x73401;
  wire x73403, x73404, x73405, x73406, x73408, x73409, x73410, x73411;
  wire x73413, x73414, x73415, x73416, x73418, x73419, x73420, x73421;
  wire x73423, x73424, x73425, x73426, x73428, x73429, x73430, x73431;
  wire x73433, x73434, x73435, x73436, x73438, x73439, x73440, x73441;
  wire x73443, x73444, x73445, x73446, x73448, x73449, x73450, x73451;
  wire x73453, x73454, x73455, x73456, x73458, x73459, x73460, x73461;
  wire x73463, x73464, x73465, x73466, x73468, x73469, x73470, x73471;
  wire x73473, x73474, x73475, x73476, x73478, x73479, x73480, x73481;
  wire x73483, x73484, x73485, x73486, x73488, x73489, x73490, x73491;
  wire x73493, x73494, x73495, x73496, x73498, x73499, x73500, x73501;
  wire x73503, x73504, x73505, x73506, x73508, x73509, x73510, x73511;
  wire x73513, x73514, x73515, x73516, x73518, x73519, x73520, x73521;
  wire x73523, x73524, x73525, x73526, x73528, x73529, x73530, x73531;
  wire x73533, x73534, x73535, x73536, x73538, x73539, x73540, x73541;
  wire x73543, x73544, x73545, x73546, x73548, x73549, x73550, x73551;
  wire x73553, x73554, x73555, x73556, x73558, x73559, x73560, x73561;
  wire x73563, x73564, x73565, x73566, x73568, x73569, x73570, x73571;
  wire x73573, x73574, x73575, x73576, x73578, x73579, x73580, x73581;
  wire x73583, x73584, x73585, x73586, x73588, x73589, x73590, x73591;
  wire x73593, x73594, x73595, x73596, x73598, x73599, x73600, x73601;
  wire x73603, x73604, x73605, x73606, x73608, x73609, x73610, x73611;
  wire x73613, x73614, x73615, x73616, x73618, x73619, x73620, x73621;
  wire x73623, x73624, x73625, x73626, x73628, x73629, x73630, x73631;
  wire x73633, x73634, x73635, x73636, x73638, x73639, x73640, x73641;
  wire x73643, x73644, x73645, x73646, x73648, x73649, x73650, x73651;
  wire x73653, x73654, x73655, x73656, x73658, x73659, x73660, x73661;
  wire x73663, x73664, x73665, x73666, x73668, x73669, x73670, x73671;
  wire x73673, x73674, x73675, x73676, x73678, x73679, x73680, x73681;
  wire x73683, x73684, x73685, x73686, x73688, x73689, x73690, x73691;
  wire x73693, x73694, x73695, x73696, x73698, x73699, x73700, x73701;
  wire x73703, x73704, x73705, x73706, x73708, x73709, x73710, x73711;
  wire x73713, x73714, x73715, x73716, x73718, x73719, x73720, x73721;
  wire x73723, x73724, x73725, x73726, x73728, x73729, x73730, x73731;
  wire x73733, x73734, x73735, x73736, x73738, x73739, x73740, x73741;
  wire x73743, x73744, x73745, x73746, x73748, x73749, x73750, x73751;
  wire x73753, x73754, x73755, x73756, x73758, x73759, x73760, x73761;
  wire x73763, x73764, x73765, x73766, x73768, x73769, x73770, x73771;
  wire x73773, x73774, x73775, x73776, x73778, x73779, x73780, x73781;
  wire x73783, x73784, x73785, x73786, x73788, x73789, x73790, x73791;
  wire x73793, x73794, x73795, x73796, x73798, x73799, x73800, x73801;
  wire x73803, x73804, x73805, x73806, x73808, x73809, x73810, x73811;
  wire x73813, x73814, x73815, x73816, x73818, x73819, x73820, x73821;
  wire x73823, x73824, x73825, x73826, x73828, x73829, x73830, x73831;
  wire x73833, x73834, x73835, x73836, x73838, x73839, x73840, x73841;
  wire x73843, x73844, x73845, x73846, x73848, x73849, x73850, x73851;
  wire x73853, x73854, x73855, x73856, x73858, x73859, x73860, x73861;
  wire x73863, x73864, x73865, x73866, x73868, x73869, x73870, x73871;
  wire x73873, x73874, x73875, x73876, x73878, x73879, x73880, x73881;
  wire x73883, x73884, x73885, x73886, x73888, x73889, x73890, x73891;
  wire x73893, x73894, x73895, x73896, x73898, x73899, x73900, x73901;
  wire x73903, x73904, x73905, x73906, x73908, x73909, x73910, x73911;
  wire x73913, x73914, x73915, x73916, x73918, x73919, x73920, x73921;
  wire x73923, x73924, x73925, x73926, x73928, x73929, x73930, x73931;
  wire x73933, x73934, x73935, x73936, x73938, x73939, x73940, x73941;
  wire x73943, x73944, x73945, x73946, x73948, x73949, x73950, x73951;
  wire x73953, x73954, x73955, x73956, x73958, x73959, x73960, x73961;
  wire x73963, x73964, x73965, x73966, x73968, x73969, x73970, x73971;
  wire x73973, x73974, x73975, x73976, x73978, x73979, x73980, x73981;
  wire x73983, x73984, x73985, x73986, x73988, x73989, x73990, x73991;
  wire x73993, x73994, x73995, x73996, x73998, x73999, x74000, x74001;
  wire x74003, x74004, x74006, x74007, x74009, x74010, x74012, x74013;
  wire x74015, x74016, x74018, x74019, x74021, x74022, x74024, x74025;
  wire x74027, x74028, x74030, x74031, x74033, x74034, x74036, x74037;
  wire x74039, x74040, x74042, x74043, x74045, x74046, x74048, x74049;
  wire x74051, x74052, x74054, x74055, x74057, x74058, x74060, x74061;
  wire x74063, x74064, x74066, x74067, x74069, x74070, x74072, x74073;
  wire x74075, x74076, x74078, x74079, x74081, x74082, x74084, x74085;
  wire x74087, x74088, x74090, x74091, x74093, x74094, x74096, x74097;
  wire x74099, x74100, x74102, x74103, x74105, x74106, x74108, x74109;
  wire x74111, x74112, x74114, x74115, x74117, x74118, x74120, x74121;
  wire x74123, x74124, x74126, x74127, x74129, x74130, x74132, x74133;
  wire x74135, x74136, x74138, x74139, x74141, x74142, x74144, x74145;
  wire x74147, x74148, x74150, x74151, x74153, x74154, x74156, x74157;
  wire x74159, x74160, x74162, x74163, x74165, x74166, x74168, x74169;
  wire x74171, x74172, x74174, x74175, x74177, x74178, x74180, x74181;
  wire x74183, x74184, x74186, x74187, x74189, x74190, x74192, x74193;
  wire x74195, x74196, x74198, x74199, x74201, x74202, x74204, x74205;
  wire x74207, x74208, x74210, x74211, x74213, x74214, x74216, x74217;
  wire x74219, x74220, x74222, x74223, x74225, x74226, x74228, x74229;
  wire x74231, x74232, x74234, x74235, x74237, x74238, x74240, x74241;
  wire x74243, x74244, x74246, x74247, x74249, x74250, x74252, x74253;
  wire x74255, x74256, x74258, x74259, x74261, x74262, x74264, x74265;
  wire x74267, x74268, x74270, x74271, x74273, x74274, x74276, x74277;
  wire x74279, x74280, x74282, x74283, x74285, x74286, x74288, x74289;
  wire x74291, x74292, x74294, x74295, x74297, x74298, x74300, x74301;
  wire x74303, x74304, x74306, x74307, x74309, x74310, x74312, x74313;
  wire x74315, x74316, x74318, x74319, x74321, x74322, x74324, x74325;
  wire x74327, x74328, x74330, x74331, x74333, x74334, x74336, x74337;
  wire x74339, x74340, x74342, x74343, x74345, x74346, x74348, x74349;
  wire x74351, x74352, x74354, x74355, x74357, x74358, x74360, x74361;
  wire x74363, x74364, x74366, x74367, x74369, x74370, x74372, x74373;
  wire x74375, x74376, x74378, x74379, x74381, x74382, x74384, x74385;
  wire x74387, x74388, x74390, x74391, x74393, x74394, x74396, x74397;
  wire x74399, x74400, x74402, x74403, x74405, x74406, x74408, x74409;
  wire x74411, x74412, x74414, x74415, x74417, x74418, x74420, x74421;
  wire x74423, x74424, x74426, x74427, x74429, x74430, x74432, x74433;
  wire x74435, x74436, x74438, x74439, x74441, x74442, x74444, x74445;
  wire x74447, x74448, x74450, x74451, x74453, x74454, x74456, x74457;
  wire x74459, x74460, x74462, x74463, x74465, x74466, x74468, x74469;
  wire x74471, x74472, x74474, x74475, x74477, x74478, x74480, x74481;
  wire x74483, x74484, x74486, x74487, x74489, x74490, x74492, x74493;
  wire x74495, x74496, x74498, x74499, x74501, x74502, x74504, x74505;
  wire x74507, x74508, x74510, x74511, x74513, x74514, x74516, x74517;
  wire x74519, x74520, x74522, x74523, x74525, x74526, x74528, x74529;
  wire x74531, x74532, x74534, x74535, x74537, x74538, x74540, x74541;
  wire x74543, x74544, x74546, x74547, x74549, x74550, x74552, x74553;
  wire x74555, x74556, x74558, x74559, x74561, x74562, x74564, x74565;
  wire x74567, x74568, x74570, x74571, x74573, x74574, x74576, x74577;
  wire x74579, x74580, x74582, x74583, x74585, x74586, x74588, x74589;
  wire x74591, x74592, x74594, x74595, x74597, x74598, x74600, x74601;
  wire x74603, x74604, x74606, x74607, x74609, x74610, x74612, x74613;
  wire x74615, x74616, x74618, x74619, x74621, x74622, x74624, x74625;
  wire x74627, x74628, x74630, x74631, x74633, x74634, x74636, x74637;
  wire x74639, x74640, x74642, x74643, x74645, x74646, x74648, x74649;
  wire x74651, x74652, x74654, x74655, x74657, x74658, x74660, x74661;
  wire x74663, x74664, x74666, x74667, x74669, x74670, x74672, x74673;
  wire x74675, x74676, x74678, x74679, x74681, x74682, x74684, x74685;
  wire x74687, x74688, x74690, x74691, x74693, x74694, x74696, x74697;
  wire x74699, x74700, x74702, x74703, x74705, x74706, x74708, x74709;
  wire x74711, x74712, x74714, x74715, x74717, x74718, x74720, x74721;
  wire x74723, x74724, x74726, x74727, x74729, x74730, x74732, x74733;
  wire x74735, x74736, x74738, x74739, x74741, x74742, x74744, x74745;
  wire x74747, x74748, x74750, x74751, x74753, x74754, x74756, x74757;
  wire x74759, x74760, x74762, x74763, x74765, x74766, x74768, x74769;
  wire x74771, x74772, x74774, x74775, x74777, x74778, x74780, x74781;
  wire x74783, x74784, x74786, x74787, x74789, x74790, x74792, x74793;
  wire x74795, x74796, x74798, x74799, x74801, x74802, x74804, x74805;
  wire x74807, x74808, x74810, x74811, x74813, x74814, x74816, x74817;
  wire x74819, x74820, x74822, x74823, x74825, x74826, x74828, x74829;
  wire x74831, x74832, x74834, x74835, x74837, x74838, x74840, x74841;
  wire x74843, x74844, x74846, x74847, x74849, x74850, x74852, x74853;
  wire x74855, x74856, x74858, x74859, x74861, x74862, x74864, x74865;
  wire x74867, x74868, x74870, x74871, x74873, x74874, x74876, x74877;
  wire x74879, x74880, x74882, x74883, x74885, x74886, x74888, x74889;
  wire x74891, x74892, x74894, x74895, x74897, x74898, x74900, x74901;
  wire x74903, x74904, x74906, x74907, x74909, x74910, x74912, x74913;
  wire x74915, x74916, x74918, x74919, x74921, x74922, x74924, x74925;
  wire x74927, x74928, x74930, x74931, x74933, x74934, x74936, x74937;
  wire x74939, x74940, x74942, x74943, x74945, x74946, x74948, x74949;
  wire x74951, x74952, x74954, x74955, x74957, x74958, x74960, x74961;
  wire x74963, x74964, x74966, x74967, x74969, x74970, x74972, x74973;
  wire x74975, x74976, x74978, x74979, x74981, x74982, x74984, x74985;
  wire x74987, x74988, x74990, x74991, x74993, x74994, x74996, x74997;
  wire x74999, x75000, x75002, x75003, x75005, x75006, x75008, x75009;
  wire x75011, x75012, x75014, x75015, x75017, x75018, x75020, x75021;
  wire x75023, x75024, x75026, x75027, x75029, x75030, x75032, x75033;
  wire x75035, x75036, x75038, x75039, x75041, x75042, x75044, x75045;
  wire x75047, x75048, x75050, x75051, x75053, x75054, x75056, x75057;
  wire x75059, x75060, x75062, x75063, x75065, x75066, x75068, x75069;
  wire x75071, x75072, x75074, x75075, x75077, x75078, x75080, x75081;
  wire x75083, x75084, x75086, x75087, x75089, x75090, x75092, x75093;
  wire x75095, x75096, x75098, x75099, x75101, x75102, x75104, x75105;
  wire x75107, x75108, x75110, x75111, x75113, x75114, x75116, x75117;
  wire x75119, x75120, x75122, x75123, x75125, x75126, x75128, x75129;
  wire x75131, x75132, x75134, x75135, x75137, x75138, x75140, x75141;
  wire x75143, x75144, x75146, x75147, x75149, x75150, x75152, x75153;
  wire x75155, x75156, x75158, x75159, x75161, x75162, x75164, x75165;
  wire x75167, x75168, x75170, x75171, x75173, x75174, x75176, x75177;
  wire x75179, x75180, x75182, x75183, x75185, x75186, x75188, x75189;
  wire x75191, x75192, x75194, x75195, x75197, x75198, x75200, x75201;
  wire x75203, x75204, x75206, x75207, x75209, x75210, x75212, x75213;
  wire x75215, x75216, x75218, x75219, x75221, x75222, x75224, x75225;
  wire x75227, x75228, x75230, x75231, x75233, x75234, x75236, x75237;
  wire x75239, x75240, x75242, x75243, x75245, x75246, x75248, x75249;
  wire x75251, x75252, x75254, x75255, x75257, x75258, x75260, x75261;
  wire x75263, x75264, x75266, x75267, x75269, x75270, x75272, x75273;
  wire x75275, x75276, x75278, x75279, x75281, x75282, x75284, x75285;
  wire x75287, x75288, x75290, x75291, x75293, x75294, x75296, x75297;
  wire x75299, x75300, x75302, x75303, x75305, x75306, x75308, x75309;
  wire x75311, x75312, x75314, x75315, x75317, x75318, x75320, x75321;
  wire x75323, x75324, x75326, x75327, x75329, x75330, x75332, x75333;
  wire x75335, x75336, x75338, x75339, x75341, x75342, x75344, x75345;
  wire x75347, x75348, x75350, x75351, x75353, x75354, x75356, x75357;
  wire x75359, x75360, x75362, x75363, x75365, x75366, x75368, x75369;
  wire x75371, x75372, x75374, x75375, x75377, x75378, x75380, x75381;
  wire x75383, x75384, x75386, x75387, x75389, x75390, x75392, x75393;
  wire x75395, x75396, x75398, x75399, x75401, x75402, x75404, x75405;
  wire x75407, x75408, x75410, x75411, x75413, x75414, x75416, x75417;
  wire x75419, x75420, x75422, x75423, x75425, x75426, x75428, x75429;
  wire x75431, x75432, x75434, x75435, x75437, x75438, x75440, x75441;
  wire x75443, x75444, x75446, x75447, x75449, x75450, x75452, x75453;
  wire x75455, x75456, x75458, x75459, x75461, x75462, x75464, x75465;
  wire x75467, x75468, x75470, x75471, x75473, x75474, x75476, x75477;
  wire x75479, x75480, x75482, x75483, x75485, x75486, x75488, x75489;
  wire x75491, x75492, x75494, x75495, x75497, x75498, x75500, x75501;
  wire x75503, x75504, x75506, x75507, x75509, x75510, x75512, x75513;
  wire x75515, x75516, x75518, x75519, x75521, x75522, x75524, x75525;
  wire x75527, x75528, x75530, x75531, x75533, x75534, x75536, x75537;
  wire x75539, x75540, x75542, x75543, x75545, x75546, x75548, x75549;
  wire x75551, x75552, x75554, x75555, x75557, x75558, x75560, x75561;
  wire x75563, x75564, x75566, x75567, x75569, x75570, x75572, x75573;
  wire x75575, x75576, x75578, x75579, x75581, x75582, x75584, x75585;
  wire x75587, x75588, x75590, x75591, x75593, x75594, x75596, x75597;
  wire x75599, x75600, x75602, x75603, x75605, x75606, x75608, x75609;
  wire x75611, x75612, x75614, x75615, x75617, x75618, x75620, x75621;
  wire x75623, x75624, x75626, x75627, x75629, x75630, x75632, x75633;
  wire x75635, x75636, x75638, x75639, x75641, x75642, x75644, x75645;
  wire x75647, x75648, x75650, x75651, x75653, x75654, x75656, x75657;
  wire x75659, x75660, x75662, x75663, x75665, x75666, x75668, x75669;
  wire x75671, x75672, x75674, x75675, x75677, x75678, x75680, x75681;
  wire x75683, x75684, x75686, x75687, x75689, x75690, x75692, x75693;
  wire x75695, x75696, x75698, x75699, x75701, x75702, x75704, x75705;
  wire x75707, x75708, x75710, x75711, x75713, x75714, x75716, x75717;
  wire x75719, x75720, x75722, x75723, x75725, x75726, x75728, x75729;
  wire x75731, x75732, x75734, x75735, x75737, x75738, x75740, x75741;
  wire x75743, x75744, x75746, x75747, x75749, x75750, x75752, x75753;
  wire x75755, x75756, x75758, x75759, x75761, x75762, x75764, x75765;
  wire x75767, x75768, x75770, x75771, x75773, x75774, x75776, x75777;
  wire x75779, x75780, x75782, x75783, x75785, x75786, x75788, x75789;
  wire x75791, x75792, x75794, x75795, x75797, x75798, x75800, x75801;
  wire x75803, x75804, x75806, x75807, x75809, x75810, x75812, x75813;
  wire x75815, x75816, x75818, x75819, x75821, x75822, x75824, x75825;
  wire x75827, x75828, x75830, x75831, x75833, x75834, x75836, x75837;
  wire x75839, x75840, x75842, x75843, x75845, x75846, x75848, x75849;
  wire x75851, x75852, x75854, x75855, x75857, x75858, x75860, x75861;
  wire x75863, x75864, x75866, x75867, x75869, x75870, x75872, x75873;
  wire x75875, x75876, x75878, x75879, x75881, x75882, x75884, x75885;
  wire x75887, x75888, x75890, x75891, x75893, x75894, x75896, x75897;
  wire x75899, x75900, x75902, x75903, x75905, x75906, x75908, x75909;
  wire x75911, x75912, x75914, x75915, x75917, x75918, x75920, x75921;
  wire x75923, x75924, x75926, x75927, x75929, x75930, x75932, x75933;
  wire x75935, x75936, x75938, x75939, x75941, x75942, x75944, x75945;
  wire x75947, x75948, x75950, x75951, x75953, x75954, x75956, x75957;
  wire x75959, x75960, x75962, x75963, x75965, x75966, x75968, x75969;
  wire x75971, x75972, x75974, x75975, x75977, x75978, x75980, x75981;
  wire x75983, x75984, x75986, x75987, x75989, x75990, x75992, x75993;
  wire x75995, x75996, x75998, x75999, x76001, x76002, x76004, x76005;
  wire x76007, x76008, x76010, x76011, x76013, x76014, x76016, x76017;
  wire x76019, x76020, x76022, x76023, x76025, x76026, x76028, x76029;
  wire x76031, x76032, x76034, x76035, x76037, x76038, x76040, x76041;
  wire x76043, x76044, x76046, x76047, x76049, x76050, x76052, x76053;
  wire x76055, x76056, x76058, x76059, x76061, x76062, x76064, x76065;
  wire x76067, x76068, x76070, x76071, x76073, x76074, x76076, x76077;
  wire x76079, x76080, x76082, x76083, x76085, x76086, x76088, x76089;
  wire x76091, x76092, x76094, x76095, x76097, x76098, x76100, x76101;
  wire x76103, x76104, x76106, x76107, x76109, x76110, x76112, x76113;
  wire x76115, x76116, x76118, x76119, x76121, x76122, x76124, x76125;
  wire x76127, x76128, x76130, x76131, x76133, x76134, x76136, x76137;
  wire x76139, x76140, x76142, x76143, x76145, x76146, x76148, x76149;
  wire x76151, x76152, x76154, x76155, x76157, x76158, x76160, x76161;
  wire x76163, x76164, x76166, x76167, x76169, x76170, x76172, x76173;
  wire x76175, x76176, x76178, x76179, x76181, x76182, x76184, x76185;
  wire x76187, x76188, x76190, x76191, x76193, x76194, x76196, x76197;
  wire x76199, x76200, x76202, x76203, x76205, x76206, x76208, x76209;
  wire x76211, x76212, x76214, x76215, x76217, x76218, x76220, x76221;
  wire x76223, x76224, x76226, x76227, x76229, x76230, x76232, x76233;
  wire x76235, x76236, x76238, x76239, x76241, x76242, x76244, x76245;
  wire x76247, x76248, x76250, x76251, x76253, x76254, x76256, x76257;
  wire x76259, x76260, x76262, x76263, x76265, x76266, x76268, x76269;
  wire x76271, x76272, x76274, x76275, x76277, x76278, x76280, x76281;
  wire x76283, x76284, x76286, x76287, x76289, x76290, x76292, x76293;
  wire x76295, x76296, x76298, x76299, x76301, x76302, x76304, x76305;
  wire x76307, x76308, x76310, x76311, x76313, x76314, x76316, x76317;
  wire x76319, x76320, x76322, x76323, x76325, x76326, x76328, x76329;
  wire x76331, x76332, x76334, x76335, x76337, x76338, x76340, x76341;
  wire x76343, x76344, x76346, x76347, x76349, x76350, x76352, x76353;
  wire x76355, x76356, x76358, x76359, x76361, x76362, x76364, x76365;
  wire x76367, x76368, x76370, x76371, x76373, x76374, x76376, x76377;
  wire x76379, x76380, x76382, x76383, x76385, x76386, x76388, x76389;
  wire x76391, x76392, x76394, x76395, x76397, x76398, x76400, x76401;
  wire x76403, x76404, x76406, x76407, x76409, x76410, x76412, x76413;
  wire x76415, x76416, x76418, x76419, x76421, x76422, x76424, x76425;
  wire x76427, x76428, x76430, x76431, x76433, x76434, x76436, x76437;
  wire x76439, x76440, x76442, x76443, x76445, x76446, x76448, x76449;
  wire x76451, x76452, x76454, x76455, x76457, x76458, x76460, x76461;
  wire x76463, x76464, x76466, x76467, x76469, x76470, x76472, x76473;
  wire x76475, x76476, x76478, x76479, x76481, x76482, x76484, x76485;
  wire x76487, x76488, x76490, x76491, x76493, x76494, x76496, x76497;
  wire x76499, x76500, x76502, x76503, x76505, x76506, x76508, x76509;
  wire x76511, x76512, x76514, x76515, x76517, x76518, x76520, x76521;
  wire x76523, x76524, x76526, x76527, x76529, x76530, x76532, x76533;
  wire x76535, x76536, x76538, x76539, x76541, x76542, x76544, x76545;
  wire x76547, x76548, x76550, x76551, x76553, x76554, x76556, x76557;
  wire x76559, x76560, x76562, x76563, x76565, x76566, x76568, x76569;
  wire x76571, x76572, x76574, x76575, x76577, x76578, x76580, x76581;
  wire x76583, x76584, x76586, x76587, x76589, x76590, x76592, x76593;
  wire x76595, x76596, x76598, x76599, x76601, x76602, x76604, x76605;
  wire x76607, x76608, x76610, x76611, x76613, x76614, x76616, x76617;
  wire x76619, x76620, x76622, x76623, x76625, x76626, x76628, x76629;
  wire x76631, x76632, x76634, x76635, x76637, x76638, x76640, x76641;
  wire x76643, x76644, x76646, x76647, x76649, x76650, x76652, x76653;
  wire x76655, x76656, x76658, x76659, x76661, x76662, x76664, x76665;
  wire x76667, x76668, x76670, x76671, x76673, x76674, x76676, x76677;
  wire x76679, x76680, x76682, x76683, x76685, x76686, x76688, x76689;
  wire x76691, x76692, x76694, x76695, x76697, x76698, x76700, x76701;
  wire x76703, x76704, x76706, x76707, x76709, x76710, x76712, x76713;
  wire x76715, x76716, x76718, x76719, x76721, x76722, x76724, x76725;
  wire x76727, x76728, x76730, x76731, x76733, x76734, x76736, x76737;
  wire x76739, x76740, x76742, x76743, x76745, x76746, x76748, x76749;
  wire x76751, x76752, x76754, x76755, x76757, x76758, x76760, x76761;
  wire x76763, x76764, x76766, x76767, x76769, x76770, x76772, x76773;
  wire x76775, x76776, x76778, x76779, x76781, x76782, x76784, x76785;
  wire x76787, x76788, x76790, x76791, x76793, x76794, x76796, x76797;
  wire x76799, x76800, x76802, x76803, x76805, x76806, x76808, x76809;
  wire x76811, x76812, x76814, x76815, x76817, x76818, x76820, x76821;
  wire x76823, x76824, x76826, x76827, x76829, x76830, x76832, x76833;
  wire x76835, x76836, x76838, x76839, x76841, x76842, x76844, x76845;
  wire x76847, x76848, x76850, x76851, x76853, x76854, x76856, x76857;
  wire x76859, x76860, x76862, x76863, x76865, x76866, x76868, x76869;
  wire x76871, x76872, x76874, x76875, x76877, x76878, x76880, x76881;
  wire x76883, x76884, x76886, x76887, x76889, x76890, x76892, x76893;
  wire x76895, x76896, x76898, x76899, x76901, x76902, x76904, x76905;
  wire x76907, x76908, x76910, x76911, x76913, x76914, x76916, x76917;
  wire x76919, x76920, x76922, x76923, x76925, x76926, x76928, x76929;
  wire x76931, x76932, x76934, x76935, x76937, x76938, x76940, x76941;
  wire x76943, x76944, x76946, x76947, x76949, x76950, x76952, x76953;
  wire x76955, x76956, x76958, x76959, x76961, x76962, x76964, x76965;
  wire x76967, x76968, x76970, x76971, x76973, x76974, x76976, x76977;
  wire x76979, x76980, x76982, x76983, x76985, x76986, x76988, x76989;
  wire x76991, x76992, x76994, x76995, x76997, x76998, x77000, x77001;
  wire x77003, x77004, x77006, x77007, x77009, x77010, x77012, x77013;
  wire x77015, x77016, x77018, x77019, x77021, x77022, x77024, x77025;
  wire x77027, x77028, x77030, x77031, x77033, x77034, x77036, x77037;
  wire x77039, x77040, x77042, x77043, x77045, x77046, x77048, x77049;
  wire x77051, x77052, x77054, x77055, x77057, x77058, x77060, x77061;
  wire x77063, x77064, x77066, x77067, x77069, x77070, x77072, x77073;
  wire x77075, x77076, x77078, x77079, x77081, x77082, x77084, x77085;
  wire x77087, x77088, x77090, x77091, x77093, x77094, x77096, x77097;
  wire x77099, x77100, x77102, x77103, x77105, x77106, x77108, x77109;
  wire x77111, x77112, x77114, x77115, x77117, x77118, x77120, x77121;
  wire x77123, x77124, x77126, x77127, x77129, x77130, x77132, x77133;
  wire x77135, x77136, x77138, x77139, x77141, x77142, x77144, x77145;
  wire x77147, x77148, x77150, x77151, x77153, x77154, x77156, x77157;
  wire x77159, x77160, x77162, x77163, x77165, x77166, x77168, x77169;
  wire x77171, x77172, x77174, x77175, x77177, x77178, x77180, x77181;
  wire x77183, x77184, x77186, x77187, x77189, x77190, x77192, x77193;
  wire x77195, x77196, x77198, x77199, x77201, x77202, x77204, x77205;
  wire x77207, x77208, x77210, x77211, x77213, x77214, x77216, x77217;
  wire x77219, x77220, x77222, x77223, x77225, x77226, x77228, x77229;
  wire x77231, x77232, x77234, x77235, x77237, x77238, x77240, x77241;
  wire x77243, x77244, x77246, x77247, x77249, x77250, x77252, x77253;
  wire x77255, x77256, x77258, x77259, x77261, x77262, x77264, x77265;
  wire x77267, x77268, x77270, x77271, x77273, x77274, x77276, x77277;
  wire x77279, x77280, x77282, x77283, x77285, x77286, x77288, x77289;
  wire x77291, x77292, x77294, x77295, x77297, x77298, x77300, x77301;
  wire x77303, x77304, x77306, x77307, x77309, x77310, x77312, x77313;
  wire x77315, x77316, x77318, x77319, x77321, x77322, x77324, x77325;
  wire x77327, x77328, x77330, x77331, x77333, x77334, x77336, x77337;
  wire x77339, x77340, x77342, x77343, x77345, x77346, x77348, x77349;
  wire x77351, x77352, x77354, x77355, x77357, x77358, x77360, x77361;
  wire x77363, x77364, x77366, x77367, x77369, x77370, x77372, x77373;
  wire x77375, x77376, x77378, x77379, x77381, x77382, x77384, x77385;
  wire x77387, x77388, x77390, x77391, x77393, x77394, x77396, x77397;
  wire x77399, x77400, x77402, x77403, x77405, x77406, x77408, x77409;
  wire x77411, x77412, x77414, x77415, x77417, x77418, x77420, x77421;
  wire x77423, x77424, x77426, x77427, x77429, x77430, x77432, x77433;
  wire x77435, x77436, x77438, x77439, x77441, x77442, x77444, x77445;
  wire x77447, x77448, x77450, x77451, x77453, x77454, x77456, x77457;
  wire x77459, x77460, x77462, x77463, x77465, x77466, x77468, x77469;
  wire x77471, x77472, x77474, x77475, x77477, x77478, x77480, x77481;
  wire x77483, x77484, x77486, x77487, x77489, x77490, x77492, x77493;
  wire x77495, x77496, x77498, x77499, x77501, x77502, x77504, x77505;
  wire x77507, x77508, x77510, x77511, x77513, x77514, x77516, x77517;
  wire x77519, x77520, x77522, x77523, x77525, x77526, x77528, x77529;
  wire x77531, x77532, x77534, x77535, x77537, x77538, x77540, x77541;
  wire x77543, x77544, x77546, x77547, x77549, x77550, x77552, x77553;
  wire x77555, x77556, x77558, x77559, x77561, x77562, x77564, x77565;
  wire x77567, x77568, x77570, x77571, x77573, x77574, x77576, x77577;
  wire x77579, x77580, x77582, x77583, x77585, x77586, x77588, x77589;
  wire x77591, x77592, x77594, x77595, x77597, x77598, x77600, x77601;
  wire x77603, x77604, x77606, x77607, x77609, x77610, x77612, x77613;
  wire x77615, x77616, x77618, x77619, x77621, x77622, x77624, x77625;
  wire x77627, x77628, x77630, x77631, x77633, x77634, x77636, x77637;
  wire x77639, x77640, x77642, x77643, x77645, x77646, x77648, x77649;
  wire x77651, x77652, x77654, x77655, x77657, x77658, x77660, x77661;
  wire x77663, x77664, x77666, x77667, x77669, x77670, x77672, x77673;
  wire x77675, x77676, x77678, x77679, x77681, x77682, x77684, x77685;
  wire x77687, x77688, x77690, x77691, x77693, x77694, x77696, x77697;
  wire x77699, x77700, x77702, x77703, x77705, x77706, x77708, x77709;
  wire x77711, x77712, x77714, x77715, x77717, x77718, x77720, x77721;
  wire x77723, x77724, x77726, x77727, x77729, x77730, x77732, x77733;
  wire x77735, x77736, x77738, x77739, x77741, x77742, x77744, x77745;
  wire x77747, x77748, x77750, x77751, x77753, x77754, x77756, x77757;
  wire x77759, x77760, x77762, x77763, x77765, x77766, x77768, x77769;
  wire x77771, x77772, x77774, x77775, x77777, x77778, x77780, x77781;
  wire x77783, x77784, x77786, x77787, x77789, x77790, x77792, x77793;
  wire x77795, x77796, x77798, x77799, x77801, x77802, x77804, x77805;
  wire x77807, x77808, x77810, x77811, x77813, x77814, x77816, x77817;
  wire x77819, x77820, x77822, x77823, x77825, x77826, x77828, x77829;
  wire x77831, x77832, x77834, x77835, x77837, x77838, x77840, x77841;
  wire x77843, x77844, x77846, x77847, x77849, x77850, x77852, x77853;
  wire x77855, x77856, x77858, x77859, x77861, x77862, x77864, x77865;
  wire x77867, x77868, x77870, x77871, x77873, x77874, x77876, x77877;
  wire x77879, x77880, x77882, x77883, x77885, x77886, x77888, x77889;
  wire x77891, x77892, x77894, x77895, x77897, x77898, x77900, x77901;
  wire x77903, x77904, x77906, x77907, x77909, x77910, x77912, x77913;
  wire x77915, x77916, x77918, x77919, x77921, x77922, x77924, x77925;
  wire x77927, x77928, x77930, x77931, x77933, x77934, x77936, x77937;
  wire x77939, x77940, x77942, x77943, x77945, x77946, x77948, x77949;
  wire x77951, x77952, x77954, x77955, x77957, x77958, x77960, x77961;
  wire x77963, x77964, x77966, x77967, x77969, x77970, x77972, x77973;
  wire x77975, x77976, x77978, x77979, x77981, x77982, x77984, x77985;
  wire x77987, x77988, x77990, x77991, x77993, x77994, x77996, x77997;
  wire x77999, x78000, x78002, x78003, x78005, x78006, x78008, x78009;
  wire x78011, x78012, x78014, x78015, x78017, x78018, x78020, x78021;
  wire x78023, x78024, x78026, x78027, x78029, x78030, x78032, x78033;
  wire x78035, x78036, x78038, x78039, x78041, x78042, x78044, x78045;
  wire x78047, x78048, x78050, x78051, x78053, x78054, x78056, x78057;
  wire x78059, x78060, x78062, x78063, x78065, x78066, x78068, x78069;
  wire x78071, x78072, x78074, x78075, x78077, x78078, x78080, x78081;
  wire x78083, x78084, x78086, x78087, x78089, x78090, x78092, x78093;
  wire x78095, x78096, x78098, x78099, x78101, x78102, x78104, x78105;
  wire x78107, x78108, x78110, x78111, x78113, x78114, x78116, x78117;
  wire x78119, x78120, x78122, x78123, x78125, x78126, x78128, x78129;
  wire x78131, x78132, x78134, x78135, x78137, x78138, x78140, x78141;
  wire x78143, x78144, x78146, x78147, x78149, x78150, x78152, x78153;
  wire x78155, x78156, x78158, x78159, x78161, x78162, x78164, x78165;
  wire x78167, x78168, x78170, x78171, x78173, x78174, x78176, x78177;
  wire x78179, x78180, x78182, x78183, x78185, x78186, x78188, x78189;
  wire x78191, x78192, x78194, x78195, x78197, x78198, x78200, x78201;
  wire x78203, x78204, x78206, x78207, x78209, x78210, x78212, x78213;
  wire x78215, x78216, x78218, x78219, x78221, x78222, x78224, x78225;
  wire x78227, x78228, x78230, x78231, x78233, x78234, x78236, x78237;
  wire x78239, x78240, x78242, x78243, x78245, x78246, x78248, x78249;
  wire x78251, x78252, x78254, x78255, x78257, x78258, x78260, x78261;
  wire x78263, x78264, x78266, x78267, x78269, x78270, x78272, x78273;
  wire x78275, x78276, x78278, x78279, x78281, x78282, x78284, x78285;
  wire x78287, x78288, x78290, x78291, x78293, x78294, x78296, x78297;
  wire x78299, x78300, x78302, x78303, x78305, x78306, x78308, x78309;
  wire x78311, x78312, x78314, x78315, x78317, x78318, x78320, x78321;
  wire x78323, x78324, x78326, x78327, x78329, x78330, x78332, x78333;
  wire x78335, x78336, x78338, x78339, x78341, x78342, x78344, x78345;
  wire x78347, x78348, x78350, x78351, x78353, x78354, x78356, x78357;
  wire x78359, x78360, x78362, x78363, x78365, x78366, x78368, x78369;
  wire x78371, x78372, x78374, x78375, x78377, x78378, x78380, x78381;
  wire x78383, x78384, x78386, x78387, x78389, x78390, x78392, x78393;
  wire x78395, x78396, x78398, x78399, x78401, x78402, x78404, x78405;
  wire x78407, x78408, x78410, x78411, x78413, x78414, x78416, x78417;
  wire x78419, x78420, x78422, x78423, x78425, x78426, x78428, x78429;
  wire x78431, x78432, x78434, x78435, x78437, x78438, x78440, x78441;
  wire x78443, x78444, x78446, x78447, x78449, x78450, x78452, x78453;
  wire x78455, x78456, x78458, x78459, x78461, x78462, x78464, x78465;
  wire x78467, x78468, x78470, x78471, x78473, x78474, x78476, x78477;
  wire x78479, x78480, x78482, x78483, x78485, x78486, x78488, x78489;
  wire x78491, x78492, x78494, x78495, x78497, x78498, x78500, x78501;
  wire x78503, x78504, x78506, x78507, x78509, x78510, x78512, x78513;
  wire x78515, x78516, x78518, x78519, x78521, x78522, x78524, x78525;
  wire x78527, x78528, x78530, x78531, x78533, x78534, x78536, x78537;
  wire x78539, x78540, x78542, x78543, x78545, x78546, x78548, x78549;
  wire x78551, x78552, x78554, x78555, x78557, x78558, x78560, x78561;
  wire x78563, x78564, x78566, x78567, x78569, x78570, x78572, x78573;
  wire x78575, x78576, x78578, x78579, x78581, x78582, x78584, x78585;
  wire x78587, x78588, x78590, x78591, x78593, x78594, x78596, x78597;
  wire x78599, x78600, x78602, x78603, x78605, x78606, x78608, x78609;
  wire x78611, x78612, x78614, x78615, x78617, x78618, x78620, x78621;
  wire x78623, x78624, x78626, x78627, x78629, x78630, x78632, x78633;
  wire x78635, x78636, x78638, x78639, x78641, x78642, x78644, x78645;
  wire x78647, x78648, x78650, x78651, x78653, x78654, x78656, x78657;
  wire x78659, x78660, x78662, x78663, x78665, x78666, x78668, x78669;
  wire x78671, x78672, x78674, x78675, x78677, x78678, x78680, x78681;
  wire x78683, x78684, x78686, x78687, x78689, x78690, x78692, x78693;
  wire x78695, x78696, x78698, x78699, x78701, x78702, x78704, x78705;
  wire x78707, x78708, x78710, x78711, x78713, x78714, x78716, x78717;
  wire x78719, x78720, x78722, x78723, x78725, x78726, x78728, x78729;
  wire x78731, x78732, x78734, x78735, x78737, x78738, x78740, x78741;
  wire x78743, x78744, x78746, x78747, x78749, x78750, x78752, x78753;
  wire x78755, x78756, x78758, x78759, x78761, x78762, x78764, x78765;
  wire x78767, x78768, x78770, x78771, x78773, x78774, x78776, x78777;
  wire x78779, x78780, x78782, x78783, x78785, x78786, x78788, x78789;
  wire x78791, x78792, x78794, x78795, x78797, x78798, x78800, x78801;
  wire x78803, x78804, x78806, x78807, x78809, x78810, x78812, x78813;
  wire x78815, x78816, x78818, x78819, x78821, x78822, x78824, x78825;
  wire x78827, x78828, x78830, x78831, x78833, x78834, x78836, x78837;
  wire x78839, x78840, x78842, x78843, x78845, x78846, x78848, x78849;
  wire x78851, x78852, x78854, x78855, x78857, x78858, x78860, x78861;
  wire x78863, x78864, x78866, x78867, x78869, x78870, x78872, x78873;
  wire x78875, x78876, x78878, x78879, x78881, x78882, x78884, x78885;
  wire x78887, x78888, x78890, x78891, x78893, x78894, x78896, x78897;
  wire x78899, x78900, x78902, x78903, x78905, x78906, x78908, x78909;
  wire x78911, x78912, x78914, x78915, x78917, x78918, x78920, x78921;
  wire x78923, x78924, x78926, x78927, x78929, x78930, x78932, x78933;
  wire x78935, x78936, x78938, x78939, x78941, x78942, x78944, x78945;
  wire x78947, x78948, x78950, x78951, x78953, x78954, x78956, x78957;
  wire x78959, x78960, x78962, x78963, x78965, x78966, x78968, x78969;
  wire x78971, x78972, x78974, x78975, x78977, x78978, x78980, x78981;
  wire x78983, x78984, x78986, x78987, x78989, x78990, x78992, x78993;
  wire x78995, x78996, x78998, x78999, x79001, x79002, x79004, x79005;
  wire x79007, x79008, x79010, x79011, x79013, x79014, x79016, x79017;
  wire x79019, x79020, x79022, x79023, x79025, x79026, x79028, x79029;
  wire x79031, x79032, x79034, x79035, x79037, x79038, x79040, x79041;
  wire x79043, x79044, x79046, x79047, x79049, x79050, x79052, x79053;
  wire x79055, x79056, x79058, x79059, x79061, x79062, x79064, x79065;
  wire x79067, x79068, x79070, x79071, x79073, x79074, x79076, x79077;
  wire x79079, x79080, x79082, x79083, x79085, x79086, x79088, x79089;
  wire x79091, x79092, x79094, x79095, x79097, x79098, x79100, x79101;
  wire x79103, x79104, x79106, x79107, x79109, x79110, x79112, x79113;
  wire x79115, x79116, x79118, x79119, x79121, x79122, x79124, x79125;
  wire x79127, x79128, x79130, x79131, x79133, x79134, x79136, x79137;
  wire x79139, x79140, x79142, x79143, x79145, x79146, x79148, x79149;
  wire x79151, x79152, x79154, x79155, x79157, x79158, x79160, x79161;
  wire x79163, x79164, x79166, x79167, x79169, x79170, x79172, x79173;
  wire x79175, x79176, x79178, x79179, x79181, x79182, x79184, x79185;
  wire x79187, x79188, x79190, x79191, x79193, x79194, x79196, x79197;
  wire x79199, x79200, x79202, x79203, x79205, x79206, x79208, x79209;
  wire x79211, x79212, x79214, x79215, x79217, x79218, x79220, x79221;
  wire x79223, x79224, x79226, x79227, x79229, x79230, x79232, x79233;
  wire x79235, x79236, x79238, x79239, x79241, x79242, x79244, x79245;
  wire x79247, x79248, x79250, x79251, x79253, x79254, x79256, x79257;
  wire x79259, x79260, x79262, x79263, x79265, x79266, x79268, x79269;
  wire x79271, x79272, x79274, x79275, x79277, x79278, x79280, x79281;
  wire x79283, x79284, x79286, x79287, x79289, x79290, x79292, x79293;
  wire x79295, x79296, x79298, x79299, x79301, x79302, x79304, x79305;
  wire x79307, x79308, x79310, x79311, x79313, x79314, x79316, x79317;
  wire x79319, x79320, x79322, x79323, x79325, x79326, x79328, x79329;
  wire x79331, x79332, x79334, x79335, x79337, x79338, x79340, x79341;
  wire x79343, x79344, x79346, x79347, x79349, x79350, x79352, x79353;
  wire x79355, x79356, x79358, x79359, x79361, x79362, x79364, x79365;
  wire x79367, x79368, x79370, x79371, x79373, x79374, x79376, x79377;
  wire x79379, x79380, x79382, x79383, x79385, x79386, x79388, x79389;
  wire x79391, x79392, x79394, x79395, x79397, x79398, x79400, x79401;
  wire x79403, x79404, x79406, x79407, x79409, x79410, x79412, x79413;
  wire x79415, x79416, x79418, x79419, x79421, x79422, x79424, x79425;
  wire x79427, x79428, x79430, x79431, x79433, x79434, x79436, x79437;
  wire x79439, x79440, x79442, x79443, x79445, x79446, x79448, x79449;
  wire x79451, x79452, x79454, x79455, x79457, x79458, x79460, x79461;
  wire x79463, x79464, x79466, x79467, x79469, x79470, x79472, x79473;
  wire x79475, x79476, x79478, x79479, x79481, x79482, x79484, x79485;
  wire x79487, x79488, x79490, x79491, x79493, x79494, x79496, x79497;
  wire x79499, x79500, x79502, x79503, x79505, x79506, x79508, x79509;
  wire x79511, x79512, x79514, x79515, x79517, x79518, x79520, x79521;
  wire x79523, x79524, x79526, x79527, x79529, x79530, x79532, x79533;
  wire x79535, x79536, x79538, x79539, x79541, x79542, x79544, x79545;
  wire x79547, x79548, x79550, x79551, x79553, x79554, x79556, x79557;
  wire x79559, x79560, x79562, x79563, x79565, x79566, x79568, x79569;
  wire x79571, x79572, x79574, x79575, x79577, x79578, x79580, x79581;
  wire x79583, x79584, x79586, x79587, x79589, x79590, x79592, x79593;
  wire x79595, x79596, x79598, x79599, x79601, x79602, x79604, x79605;
  wire x79607, x79608, x79610, x79611, x79613, x79614, x79616, x79617;
  wire x79619, x79620, x79622, x79623, x79625, x79626, x79628, x79629;
  wire x79631, x79632, x79634, x79635, x79637, x79638, x79640, x79641;
  wire x79643, x79644, x79646, x79647, x79649, x79650, x79652, x79653;
  wire x79655, x79656, x79658, x79659, x79661, x79662, x79664, x79665;
  wire x79667, x79668, x79670, x79671, x79673, x79674, x79676, x79677;
  wire x79679, x79680, x79682, x79683, x79685, x79686, x79688, x79689;
  wire x79691, x79692, x79694, x79695, x79697, x79698, x79700, x79701;
  wire x79703, x79704, x79706, x79707, x79709, x79710, x79712, x79713;
  wire x79715, x79716, x79718, x79719, x79721, x79722, x79724, x79725;
  wire x79727, x79728, x79730, x79731, x79733, x79734, x79736, x79737;
  wire x79739, x79740, x79742, x79743, x79745, x79746, x79748, x79749;
  wire x79751, x79752, x79754, x79755, x79757, x79758, x79760, x79761;
  wire x79763, x79764, x79766, x79767, x79769, x79770, x79772, x79773;
  wire x79775, x79776, x79778, x79779, x79781, x79782, x79784, x79785;
  wire x79787, x79788, x79790, x79791, x79793, x79794, x79796, x79797;
  wire x79799, x79800, x79802, x79803, x79805, x79806, x79808, x79809;
  wire x79811, x79812, x79814, x79815, x79817, x79818, x79820, x79821;
  wire x79823, x79824, x79826, x79827, x79829, x79830, x79832, x79833;
  wire x79835, x79836, x79838, x79839, x79841, x79842, x79844, x79845;
  wire x79847, x79848, x79850, x79851, x79853, x79854, x79856, x79857;
  wire x79859, x79860, x79862, x79863, x79865, x79866, x79868, x79869;
  wire x79871, x79872, x79874, x79875, x79877, x79878, x79880, x79881;
  wire x79883, x79884, x79886, x79887, x79889, x79890, x79892, x79893;
  wire x79895, x79896, x79898, x79899, x79901, x79902, x79904, x79905;
  wire x79907, x79908, x79910, x79911, x79913, x79914, x79916, x79917;
  wire x79919, x79920, x79922, x79923, x79925, x79926, x79928, x79929;
  wire x79931, x79932, x79934, x79935, x79937, x79938, x79940, x79941;
  wire x79943, x79944, x79946, x79947, x79949, x79950, x79952, x79953;
  wire x79955, x79956, x79958, x79959, x79961, x79962, x79964, x79965;
  wire x79967, x79968, x79970, x79971, x79973, x79974, x79976, x79977;
  wire x79979, x79980, x79982, x79983, x79985, x79986, x79988, x79989;
  wire x79991, x79992, x79994, x79995, x79997, x79998, x80000, x80001;
  wire x80003, x80004, x80006, x80007, x80009, x80010, x80012, x80013;
  wire x80015, x80016, x80018, x80019, x80021, x80022, x80024, x80025;
  wire x80027, x80028, x80030, x80031, x80033, x80034, x80036, x80037;
  wire x80039, x80040, x80042, x80043, x80045, x80046, x80048, x80049;
  wire x80051, x80052, x80054, x80055, x80057, x80058, x80060, x80061;
  wire x80063, x80064, x80066, x80067, x80069, x80070, x80072, x80073;
  wire x80075, x80076, x80078, x80079, x80081, x80082, x80084, x80085;
  wire x80087, x80088, x80090, x80091, x80093, x80094, x80096, x80097;
  wire x80099, x80100, x80102, x80103, x80105, x80106, x80108, x80109;
  wire x80111, x80112, x80114, x80115, x80117, x80118, x80120, x80121;
  wire x80123, x80124, x80126, x80127, x80129, x80130, x80132, x80133;
  wire x80135, x80136, x80138, x80139, x80141, x80142, x80144, x80145;
  wire x80147, x80148, x80150, x80151, x80153, x80154, x80156, x80157;
  wire x80159, x80160, x80162, x80163, x80165, x80166, x80168, x80169;
  wire x80171, x80172, x80174, x80175, x80177, x80178, x80180, x80181;
  wire x80183, x80184, x80186, x80187, x80189, x80190, x80192, x80193;
  wire x80195, x80196, x80198, x80199, x80201, x80202, x80204, x80205;
  wire x80207, x80208, x80210, x80211, x80213, x80214, x80216, x80217;
  wire x80219, x80220, x80222, x80223, x80225, x80226, x80228, x80229;
  wire x80231, x80232, x80234, x80235, x80237, x80238, x80240, x80241;
  wire x80243, x80244, x80246, x80247, x80249, x80250, x80252, x80253;
  wire x80255, x80256, x80258, x80259, x80261, x80262, x80264, x80265;
  wire x80267, x80268, x80270, x80271, x80273, x80274, x80276, x80277;
  wire x80279, x80280, x80282, x80283, x80285, x80286, x80288, x80289;
  wire x80291, x80292, x80294, x80295, x80297, x80298, x80300, x80301;
  wire x80303, x80304, x80306, x80307, x80309, x80310, x80312, x80313;
  wire x80315, x80316, x80318, x80319, x80321, x80322, x80324, x80325;
  wire x80327, x80328, x80330, x80331, x80333, x80334, x80336, x80337;
  wire x80339, x80340, x80342, x80343, x80345, x80346, x80348, x80349;
  wire x80351, x80352, x80354, x80355, x80357, x80358, x80360, x80361;
  wire x80363, x80364, x80366, x80367, x80369, x80370, x80372, x80373;
  wire x80375, x80376, x80378, x80379, x80381, x80382, x80384, x80385;
  wire x80387, x80388, x80390, x80391, x80393, x80394, x80396, x80397;
  wire x80399, x80400, x80402, x80403, x80405, x80406, x80408, x80409;
  wire x80411, x80412, x80414, x80415, x80417, x80418, x80420, x80421;
  wire x80423, x80424, x80426, x80427, x80429, x80430, x80432, x80433;
  wire x80435, x80436, x80438, x80439, x80441, x80442, x80444, x80445;
  wire x80447, x80448, x80450, x80451, x80453, x80454, x80456, x80457;
  wire x80459, x80460, x80462, x80463, x80465, x80466, x80468, x80469;
  wire x80471, x80472, x80474, x80475, x80477, x80478, x80480, x80481;
  wire x80483, x80484, x80486, x80487, x80489, x80490, x80492, x80493;
  wire x80495, x80496, x80498, x80499, x80501, x80502, x80504, x80505;
  wire x80507, x80508, x80510, x80511, x80513, x80514, x80516, x80517;
  wire x80519, x80520, x80522, x80523, x80525, x80526, x80528, x80529;
  wire x80531, x80532, x80534, x80535, x80537, x80538, x80540, x80541;
  wire x80543, x80544, x80546, x80547, x80549, x80550, x80552, x80553;
  wire x80555, x80556, x80558, x80559, x80561, x80562, x80564, x80565;
  wire x80567, x80568, x80570, x80571, x80573, x80574, x80576, x80577;
  wire x80579, x80580, x80582, x80583, x80585, x80586, x80588, x80589;
  wire x80591, x80592, x80594, x80595, x80597, x80598, x80600, x80601;
  wire x80603, x80604, x80606, x80607, x80609, x80610, x80612, x80613;
  wire x80615, x80616, x80618, x80619, x80621, x80622, x80624, x80625;
  wire x80627, x80628, x80630, x80631, x80633, x80634, x80636, x80637;
  wire x80639, x80640, x80642, x80643, x80645, x80646, x80648, x80649;
  wire x80651, x80652, x80654, x80655, x80657, x80658, x80660, x80661;
  wire x80663, x80664, x80666, x80667, x80669, x80670, x80672, x80673;
  wire x80675, x80676, x80678, x80679, x80681, x80682, x80684, x80685;
  wire x80687, x80688, x80690, x80691, x80693, x80694, x80696, x80697;
  wire x80699, x80700, x80702, x80703, x80705, x80706, x80708, x80709;
  wire x80711, x80712, x80714, x80715, x80717, x80718, x80720, x80721;
  wire x80723, x80724, x80726, x80727, x80729, x80730, x80732, x80733;
  wire x80735, x80736, x80738, x80739, x80741, x80742, x80744, x80745;
  wire x80747, x80748, x80750, x80751, x80753, x80754, x80756, x80757;
  wire x80759, x80760, x80762, x80763, x80765, x80766, x80768, x80769;
  wire x80771, x80772, x80774, x80775, x80777, x80778, x80780, x80781;
  wire x80783, x80784, x80786, x80787, x80789, x80790, x80792, x80793;
  wire x80795, x80796, x80798, x80799, x80801, x80802, x80804, x80805;
  wire x80807, x80808, x80810, x80811, x80813, x80814, x80816, x80817;
  wire x80819, x80820, x80822, x80823, x80825, x80826, x80828, x80829;
  wire x80831, x80832, x80834, x80835, x80837, x80838, x80840, x80841;
  wire x80843, x80844, x80846, x80847, x80849, x80850, x80852, x80853;
  wire x80855, x80856, x80858, x80859, x80861, x80862, x80864, x80865;
  wire x80867, x80868, x80870, x80871, x80873, x80874, x80876, x80877;
  wire x80879, x80880, x80882, x80883, x80885, x80886, x80888, x80889;
  wire x80891, x80892, x80894, x80895, x80897, x80898, x80900, x80901;
  wire x80903, x80904, x80906, x80907, x80909, x80910, x80912, x80913;
  wire x80915, x80916, x80918, x80919, x80921, x80922, x80924, x80925;
  wire x80927, x80928, x80930, x80931, x80933, x80934, x80936, x80937;
  wire x80939, x80940, x80942, x80943, x80945, x80946, x80948, x80949;
  wire x80951, x80952, x80954, x80955, x80957, x80958, x80960, x80961;
  wire x80963, x80964, x80966, x80967, x80969, x80970, x80972, x80973;
  wire x80975, x80976, x80978, x80979, x80981, x80982, x80984, x80985;
  wire x80987, x80988, x80990, x80991, x80993, x80994, x80996, x80997;
  wire x80999, x81000, x81002, x81003, x81005, x81006, x81008, x81009;
  wire x81011, x81012, x81014, x81015, x81017, x81018, x81020, x81021;
  wire x81023, x81024, x81026, x81027, x81029, x81030, x81032, x81033;
  wire x81035, x81036, x81038, x81039, x81041, x81042, x81044, x81045;
  wire x81047, x81048, x81050, x81051, x81053, x81054, x81056, x81057;
  wire x81059, x81060, x81062, x81063, x81065, x81066, x81068, x81069;
  wire x81071, x81072, x81074, x81075, x81077, x81078, x81080, x81081;
  wire x81083, x81084, x81086, x81087, x81089, x81090, x81092, x81093;
  wire x81095, x81096, x81098, x81099, x81101, x81102, x81104, x81105;
  wire x81107, x81108, x81110, x81111, x81113, x81114, x81116, x81117;
  wire x81119, x81120, x81122, x81123, x81125, x81126, x81128, x81129;
  wire x81131, x81132, x81134, x81135, x81137, x81138, x81140, x81141;
  wire x81143, x81144, x81146, x81147, x81149, x81150, x81152, x81153;
  wire x81155, x81156, x81158, x81159, x81161, x81162, x81164, x81165;
  wire x81167, x81168, x81170, x81171, x81173, x81174, x81176, x81177;
  wire x81179, x81180, x81182, x81183, x81185, x81186, x81188, x81189;
  wire x81191, x81192, x81194, x81195, x81197, x81198, x81200, x81201;
  wire x81203, x81204, x81206, x81207, x81209, x81210, x81212, x81213;
  wire x81215, x81216, x81218, x81219, x81221, x81222, x81224, x81225;
  wire x81227, x81228, x81230, x81231, x81233, x81234, x81236, x81237;
  wire x81239, x81240, x81242, x81243, x81245, x81246, x81248, x81249;
  wire x81251, x81252, x81254, x81255, x81257, x81258, x81260, x81261;
  wire x81263, x81264, x81266, x81267, x81269, x81270, x81272, x81273;
  wire x81275, x81276, x81278, x81279, x81281, x81282, x81284, x81285;
  wire x81287, x81288, x81290, x81291, x81293, x81294, x81296, x81297;
  wire x81299, x81300, x81302, x81303, x81305, x81306, x81308, x81309;
  wire x81311, x81312, x81314, x81315, x81317, x81318, x81320, x81321;
  wire x81323, x81324, x81326, x81327, x81329, x81330, x81332, x81333;
  wire x81335, x81336, x81338, x81339, x81341, x81342, x81344, x81345;
  wire x81347, x81348, x81350, x81351, x81353, x81354, x81356, x81357;
  wire x81359, x81360, x81362, x81363, x81365, x81366, x81368, x81369;
  wire x81371, x81372, x81374, x81375, x81377, x81378, x81380, x81381;
  wire x81383, x81384, x81386, x81387, x81389, x81390, x81392, x81393;
  wire x81395, x81396, x81398, x81399, x81401, x81402, x81404, x81405;
  wire x81407, x81408, x81410, x81411, x81413, x81414, x81416, x81417;
  wire x81419, x81420, x81422, x81423, x81425, x81426, x81428, x81429;
  wire x81431, x81432, x81434, x81435, x81437, x81438, x81440, x81441;
  wire x81443, x81444, x81446, x81447, x81449, x81450, x81452, x81453;
  wire x81455, x81456, x81458, x81459, x81461, x81462, x81464, x81465;
  wire x81467, x81468, x81470, x81471, x81473, x81474, x81476, x81477;
  wire x81479, x81480, x81482, x81483, x81485, x81486, x81488, x81489;
  wire x81491, x81492, x81494, x81495, x81497, x81498, x81500, x81501;
  wire x81503, x81504, x81506, x81507, x81509, x81510, x81512, x81513;
  wire x81515, x81516, x81518, x81519, x81521, x81522, x81524, x81525;
  wire x81527, x81528, x81530, x81531, x81533, x81534, x81536, x81537;
  wire x81539, x81540, x81542, x81543, x81545, x81546, x81548, x81549;
  wire x81551, x81552, x81554, x81555, x81557, x81558, x81560, x81561;
  wire x81563, x81564, x81566, x81567, x81569, x81570, x81572, x81573;
  wire x81575, x81576, x81578, x81579, x81581, x81582, x81584, x81585;
  wire x81587, x81588, x81590, x81591, x81593, x81594, x81596, x81597;
  wire x81599, x81600, x81602, x81603, x81605, x81606, x81608, x81609;
  wire x81611, x81612, x81614, x81615, x81617, x81618, x81620, x81621;
  wire x81623, x81624, x81626, x81627, x81629, x81630, x81632, x81633;
  wire x81635, x81636, x81638, x81639, x81641, x81642, x81644, x81645;
  wire x81647, x81648, x81650, x81651, x81653, x81654, x81656, x81657;
  wire x81659, x81660, x81662, x81663, x81665, x81666, x81668, x81669;
  wire x81671, x81672, x81674, x81675, x81677, x81678, x81680, x81681;
  wire x81683, x81684, x81686, x81687, x81689, x81690, x81692, x81693;
  wire x81695, x81696, x81698, x81699, x81701, x81702, x81704, x81705;
  wire x81707, x81708, x81710, x81711, x81713, x81714, x81716, x81717;
  wire x81719, x81720, x81722, x81723, x81725, x81726, x81728, x81729;
  wire x81731, x81732, x81734, x81735, x81737, x81738, x81740, x81741;
  wire x81743, x81744, x81746, x81747, x81749, x81750, x81752, x81753;
  wire x81755, x81756, x81758, x81759, x81761, x81762, x81764, x81765;
  wire x81767, x81768, x81770, x81771, x81773, x81774, x81776, x81777;
  wire x81779, x81780, x81782, x81783, x81785, x81786, x81788, x81789;
  wire x81791, x81792, x81794, x81795, x81797, x81798, x81800, x81801;
  wire x81803, x81804, x81806, x81807, x81809, x81810, x81812, x81813;
  wire x81815, x81816, x81818, x81819, x81821, x81822, x81824, x81825;
  wire x81827, x81828, x81830, x81831, x81833, x81834, x81836, x81837;
  wire x81839, x81840, x81842, x81843, x81845, x81846, x81848, x81849;
  wire x81851, x81852, x81854, x81855, x81857, x81858, x81860, x81861;
  wire x81863, x81864, x81866, x81867, x81869, x81870, x81872, x81873;
  wire x81875, x81876, x81878, x81879, x81881, x81882, x81884, x81885;
  wire x81887, x81888, x81890, x81891, x81893, x81894, x81896, x81897;
  wire x81899, x81900, x81902, x81903, x81905, x81906, x81908, x81909;
  wire x81911, x81912, x81914, x81915, x81917, x81918, x81920, x81921;
  wire x81923, x81924, x81926, x81927, x81929, x81930, x81932, x81933;
  wire x81935, x81936, x81938, x81939, x81941, x81942, x81944, x81945;
  wire x81947, x81948, x81950, x81951, x81953, x81954, x81956, x81957;
  wire x81959, x81960, x81962, x81963, x81965, x81966, x81968, x81969;
  wire x81971, x81972, x81974, x81975, x81977, x81978, x81980, x81981;
  wire x81983, x81984, x81986, x81987, x81989, x81990, x81992, x81993;
  wire x81995, x81996, x81998, x81999, x82001, x82002, x82004, x82005;
  wire x82007, x82008, x82010, x82011, x82013, x82014, x82016, x82017;
  wire x82019, x82020, x82022, x82023, x82025, x82026, x82028, x82029;
  wire x82031, x82032, x82034, x82035, x82037, x82038, x82040, x82041;
  wire x82043, x82044, x82046, x82047, x82049, x82050, x82052, x82053;
  wire x82055, x82056, x82058, x82059, x82061, x82062, x82064, x82065;
  wire x82067, x82068, x82070, x82071, x82073, x82074, x82076, x82077;
  wire x82079, x82080, x82082, x82083, x82085, x82086, x82088, x82089;
  wire x82091, x82092, x82094, x82095, x82097, x82098, x82100, x82101;
  wire x82103, x82104, x82106, x82107, x82109, x82110, x82112, x82113;
  wire x82115, x82116, x82118, x82119, x82121, x82122, x82124, x82125;
  wire x82127, x82128, x82130, x82131, x82133, x82134, x82136, x82137;
  wire x82139, x82140, x82142, x82143, x82145, x82146, x82148, x82149;
  wire x82151, x82152, x82154, x82155, x82157, x82158, x82160, x82161;
  wire x82163, x82164, x82166, x82167, x82169, x82170, x82172, x82173;
  wire x82175, x82176, x82178, x82179, x82181, x82182, x82184, x82185;
  wire x82187, x82188, x82190, x82191, x82193, x82194, x82196, x82197;
  wire x82199, x82200, x82202, x82203, x82205, x82206, x82208, x82209;
  wire x82211, x82212, x82214, x82215, x82217, x82218, x82220, x82221;
  wire x82223, x82224, x82226, x82227, x82229, x82230, x82232, x82233;
  wire x82235, x82236, x82238, x82239, x82241, x82242, x82244, x82245;
  wire x82247, x82248, x82250, x82251, x82253, x82254, x82256, x82257;
  wire x82259, x82260, x82262, x82263, x82265, x82266, x82268, x82269;
  wire x82271, x82272, x82274, x82275, x82277, x82278, x82280, x82281;
  wire x82283, x82284, x82286, x82287, x82289, x82290, x82292, x82293;
  wire x82295, x82296, x82298, x82299, x82301, x82302, x82304, x82305;
  wire x82307, x82308, x82310, x82311, x82313, x82314, x82316, x82317;
  wire x82319, x82320, x82322, x82323, x82325, x82326, x82328, x82329;
  wire x82331, x82332, x82334, x82335, x82337, x82338, x82340, x82341;
  wire x82343, x82344, x82346, x82347, x82349, x82350, x82352, x82353;
  wire x82355, x82356, x82358, x82359, x82361, x82362, x82364, x82365;
  wire x82367, x82368, x82370, x82371, x82373, x82374, x82376, x82377;
  wire x82379, x82380, x82382, x82383, x82385, x82386, x82388, x82389;
  wire x82391, x82392, x82394, x82395, x82397, x82398, x82400, x82401;
  wire x82403, x82404, x82406, x82407, x82409, x82410, x82412, x82413;
  wire x82415, x82416, x82418, x82419, x82421, x82422, x82424, x82425;
  wire x82427, x82428, x82430, x82431, x82433, x82434, x82436, x82437;
  wire x82439, x82440, x82442, x82443, x82445, x82446, x82448, x82449;
  wire x82451, x82452, x82454, x82455, x82457, x82458, x82460, x82461;
  wire x82463, x82464, x82466, x82467, x82469, x82470, x82472, x82473;
  wire x82475, x82476, x82478, x82479, x82481, x82482, x82484, x82485;
  wire x82487, x82488, x82490, x82491, x82493, x82494, x82496, x82497;
  wire x82499, x82500, x82502, x82503, x82505, x82506, x82508, x82509;
  wire x82511, x82512, x82514, x82515, x82517, x82518, x82520, x82521;
  wire x82523, x82524, x82526, x82527, x82529, x82530, x82532, x82533;
  wire x82535, x82536, x82538, x82539, x82541, x82542, x82544, x82545;
  wire x82547, x82548, x82550, x82551, x82553, x82554, x82556, x82557;
  wire x82559, x82560, x82562, x82563, x82565, x82566, x82568, x82569;
  wire x82571, x82572, x82574, x82575, x82577, x82578, x82580, x82581;
  wire x82583, x82584, x82586, x82587, x82589, x82590, x82592, x82593;
  wire x82595, x82596, x82598, x82599, x82601, x82602, x82604, x82605;
  wire x82607, x82608, x82610, x82611, x82613, x82614, x82616, x82617;
  wire x82619, x82620, x82622, x82623, x82625, x82626, x82628, x82629;
  wire x82631, x82632, x82634, x82635, x82637, x82638, x82640, x82641;
  wire x82643, x82644, x82646, x82647, x82649, x82650, x82652, x82653;
  wire x82655, x82656, x82658, x82659, x82661, x82662, x82664, x82665;
  wire x82667, x82668, x82670, x82671, x82673, x82674, x82676, x82677;
  wire x82679, x82680, x82682, x82683, x82685, x82686, x82688, x82689;
  wire x82691, x82692, x82694, x82695, x82697, x82698, x82700, x82701;
  wire x82703, x82704, x82706, x82707, x82709, x82710, x82712, x82713;
  wire x82715, x82716, x82718, x82719, x82721, x82722, x82724, x82725;
  wire x82727, x82728, x82730, x82731, x82733, x82734, x82736, x82737;
  wire x82739, x82740, x82742, x82743, x82745, x82746, x82748, x82749;
  wire x82751, x82752, x82754, x82755, x82757, x82758, x82760, x82761;
  wire x82763, x82764, x82766, x82767, x82769, x82770, x82772, x82773;
  wire x82775, x82776, x82778, x82779, x82781, x82782, x82784, x82785;
  wire x82787, x82788, x82790, x82791, x82793, x82794, x82796, x82797;
  wire x82799, x82800, x82802, x82803, x82805, x82806, x82808, x82809;
  wire x82811, x82812, x82814, x82815, x82817, x82818, x82820, x82821;
  wire x82823, x82824, x82826, x82827, x82829, x82830, x82832, x82833;
  wire x82835, x82836, x82838, x82839, x82841, x82842, x82844, x82845;
  wire x82847, x82848, x82850, x82851, x82853, x82854, x82856, x82857;
  wire x82859, x82860, x82862, x82863, x82865, x82866, x82868, x82869;
  wire x82871, x82872, x82874, x82875, x82877, x82878, x82880, x82881;
  wire x82883, x82884, x82886, x82887, x82889, x82890, x82892, x82893;
  wire x82895, x82896, x82898, x82899, x82901, x82902, x82904, x82905;
  wire x82907, x82908, x82910, x82911, x82913, x82914, x82916, x82917;
  wire x82919, x82920, x82922, x82923, x82925, x82926, x82928, x82929;
  wire x82931, x82932, x82934, x82935, x82937, x82938, x82940, x82941;
  wire x82943, x82944, x82946, x82947, x82949, x82950, x82952, x82953;
  wire x82955, x82956, x82958, x82959, x82961, x82962, x82964, x82965;
  wire x82967, x82968, x82970, x82971, x82973, x82974, x82976, x82977;
  wire x82979, x82980, x82982, x82983, x82985, x82986, x82988, x82989;
  wire x82991, x82992, x82994, x82995, x82997, x82998, x83000, x83001;
  wire x83003, x83004, x83006, x83007, x83009, x83010, x83012, x83013;
  wire x83015, x83016, x83018, x83019, x83021, x83022, x83024, x83025;
  wire x83027, x83028, x83030, x83031, x83033, x83034, x83036, x83037;
  wire x83039, x83040, x83042, x83043, x83045, x83046, x83048, x83049;
  wire x83051, x83052, x83054, x83055, x83057, x83058, x83060, x83061;
  wire x83063, x83064, x83066, x83067, x83069, x83070, x83072, x83073;
  wire x83075, x83076, x83078, x83079, x83081, x83082, x83084, x83085;
  wire x83087, x83088, x83090, x83091, x83093, x83094, x83096, x83097;
  wire x83099, x83100, x83102, x83103, x83105, x83106, x83108, x83109;
  wire x83111, x83112, x83114, x83115, x83117, x83118, x83120, x83121;
  wire x83123, x83124, x83126, x83127, x83129, x83130, x83132, x83133;
  wire x83135, x83136, x83138, x83139, x83141, x83142, x83144, x83145;
  wire x83147, x83148, x83150, x83151, x83153, x83154, x83156, x83157;
  wire x83159, x83160, x83162, x83163, x83165, x83166, x83168, x83169;
  wire x83171, x83172, x83174, x83175, x83177, x83178, x83180, x83181;
  wire x83183, x83184, x83186, x83187, x83189, x83190, x83192, x83193;
  wire x83195, x83196, x83198, x83199, x83201, x83202, x83204, x83205;
  wire x83207, x83208, x83210, x83211, x83213, x83214, x83216, x83217;
  wire x83219, x83220, x83222, x83223, x83225, x83226, x83228, x83229;
  wire x83231, x83232, x83234, x83235, x83237, x83238, x83240, x83241;
  wire x83243, x83244, x83246, x83247, x83249, x83250, x83252, x83253;
  wire x83255, x83256, x83258, x83259, x83261, x83262, x83264, x83265;
  wire x83267, x83268, x83270, x83271, x83273, x83274, x83276, x83277;
  wire x83279, x83280, x83282, x83283, x83285, x83286, x83288, x83289;
  wire x83291, x83292, x83294, x83295, x83297, x83298, x83300, x83301;
  wire x83303, x83304, x83306, x83307, x83309, x83310, x83312, x83313;
  wire x83315, x83316, x83318, x83319, x83321, x83322, x83324, x83325;
  wire x83327, x83328, x83330, x83331, x83333, x83334, x83336, x83337;
  wire x83339, x83340, x83342, x83343, x83345, x83346, x83348, x83349;
  wire x83350, x83351, x83353, x83354, x83355, x83356, x83358, x83359;
  wire x83360, x83361, x83363, x83364, x83365, x83366, x83368, x83369;
  wire x83370, x83371, x83373, x83374, x83375, x83376, x83378, x83379;
  wire x83380, x83381;

  wire x0, x1, x3, x4, x5, x6, x7, x8;
  wire x11, x13, x15, x19, x23, x27, x31, x35;
  wire x39, x64, x65, x66, x67, x68, x69, x70;
  wire x71, x72, x73, x74, x75, x76, x77, x78;
  wire x79, x80, x81, x82, x83, x84, x85, x86;
  wire x87, x88, x89, x90, x91, x92, x93, x96;
  wire x98, x100, x102, x104, x106, x108, x110, x112;
  wire x114, x116, x118, x120, x122, x124, x126, x128;
  wire x130, x132, x134, x136, x138, x140, x142, x144;
  wire x146, x148, x152, x154, x156, x158, x160, x162;
  wire x164, x166, x168, x170, x172, x174, x176, x178;
  wire x180, x182, x184, x186, x188, x190, x192, x194;
  wire x196, x198, x200, x206, x208, x210, x212, x214;
  wire x216, x218, x220, x222, x224, x226, x228, x230;
  wire x232, x234, x236, x238, x240, x242, x244, x246;
  wire x256, x258, x260, x262, x264, x266, x268, x270;
  wire x272, x274, x276, x278, x280, x296, x300, x304;
  wire x308, x312, x316, x320, x324, x328, x332, x336;
  wire x340, x344, x348, x352, x356, x360, x364, x368;
  wire x372, x376, x380, x384, x388, x392, x396, x400;
  wire x404, x408, x410, x634, x635, x636, x637, x640;
  wire x644, x648, x652, x654, x656, x678, x1000, x1001;
  wire x1003, x1005, x1007, x1009, x1011, x1012, x1014, x1016;
  wire x1018, x1020, x1022, x1024, x1026, x1028, x1031, x1033;
  wire x1035, x1038, x1040, x1042, x1046, x1048, x1050, x1052;
  wire x1059, x1062, x1068, x1075, x1077, x1079, x1081, x1083;
  wire x1085, x1087, x1089, x1091, x1093, x1095, x1097, x1101;
  wire x1103, x1106, x1110, x1116, x1125, x1127, x1129, x1131;
  wire x1133, x1135, x1137, x1139, x1141, x1145, x1148, x1152;
  wire x1159, x1161, x1162, x1163, x1164, x1168, x1169, x1170;
  wire x1172, x1175, x1177, x1179, x1180, x1181, x1183, x1186;
  wire x1188, x1190, x1193, x1194, x1196, x1198, x1200, x1201;
  wire x1203, x1205, x1207, x1209, x1210, x1212, x1214, x1216;
  wire x1218, x1220, x1222, x1224, x1226, x1228, x1234, x1240;
  wire x1246, x1252, x1258, x1264, x1270, x1276, x1280, x1282;
  wire x1284, x1290, x1296, x1302, x1308, x1314, x1320, x1326;
  wire x1332, x1338, x1344, x1350, x1356, x1362, x1368, x1374;
  wire x1378, x1380, x1382, x1388, x1394, x1400, x1406, x1412;
  wire x1418, x1424, x1437, x1444, x1448, x1461, x1468, x1472;
  wire x1485, x1492, x1684, x1686, x1688, x1690, x1693, x1695;
  wire x1697, x1699, x1701, x1703, x1705, x1707, x1709, x1711;
  wire x1714, x1717, x1724, x1725, x1727, x1729, x1731, x1732;
  wire x1734, x1736, x1738, x1740, x1741, x1751, x1754, x1757;
  wire x1759, x1761, x1764, x1767, x1769, x1771, x1774, x1777;
  wire x1779, x1781, x1784, x1787, x1789, x1791, x1794, x1797;
  wire x1799, x1801, x1804, x1807, x1809, x1811, x1814, x1817;
  wire x1819, x1821, x1824, x1827, x1829, x1893, x1896, x1897;
  wire x1899, x1901, x1902, x1903, x1904, x1905, x1906, x1907;
  wire x1908, x1910, x1936, x1962, x1988, x2014, x2040, x2066;
  wire x2092, x2244, x2247, x2250, x2253, x2256, x2267, x2278;
  wire x2279, x2281, x2283, x2285, x2286, x2288, x2290, x2292;
  wire x2294, x2295, x2297, x2299, x2301, x2303, x2305, x2307;
  wire x2309, x2311, x2313, x2443, x2573, x2703, x2833, x2963;
  wire x3093, x3223, x3353, x3357, x3359, x3485, x3615, x3745;
  wire x3875, x4005, x4135, x4265, x4395, x4403, x4405, x4527;
  wire x4657, x4787, x4917, x5047, x5177, x5307, x5437, x5441;
  wire x5443, x5447, x5449, x5571, x5701, x5831, x5961, x6091;
  wire x6221, x6351, x6481, x6494, x6501, x7156, x7169, x7176;
  wire x14555, x14557, x14560, x14567, x14568, x14571, x14573, x14575;
  wire x14577, x14579, x14581, x14591, x14594, x14597, x14599, x14601;
  wire x14604, x14607, x14609, x14611, x14614, x14617, x14619, x14621;
  wire x14624, x14627, x14629, x14631, x14634, x14637, x14639, x14641;
  wire x14644, x14647, x14649, x14651, x14654, x14657, x14659, x14661;
  wire x14664, x14667, x14669, x14733, x14735, x14737, x14739, x14741;
  wire x14743, x14746, x14748, x14751, x14752, x14754, x14755, x14756;
  wire x14757, x14758, x14759, x14760, x14761, x14763, x14789, x14815;
  wire x14841, x14867, x14893, x14919, x14945, x15096, x15152, x15217;
  wire x15219, x15222, x15224, x15227, x15229, x15231, x15232, x15236;
  wire x15237, x15240, x15242, x15243, x15246, x15248, x15249, x15252;
  wire x15254, x15255, x15258, x15260, x15261, x15264, x15266, x15267;
  wire x15270, x15272, x15273, x15276, x15278, x15279, x15282, x15284;
  wire x15285, x15288, x15290, x15291, x15294, x15296, x15297, x15300;
  wire x15302, x15303, x15306, x15308, x15309, x15312, x15314, x15315;
  wire x15318, x15320, x15321, x15324, x15326, x15327, x15330, x15332;
  wire x15333, x15336, x15338, x15339, x15342, x15344, x15345, x15348;
  wire x15350, x15351, x15354, x15356, x15357, x15360, x15362, x15365;
  wire x15367, x15370, x15372, x15375, x15377, x15380, x15382, x15385;
  wire x15387, x15390, x15392, x15395, x15397, x15400, x15402, x15405;
  wire x15407, x15410, x15411, x15412, x15413, x15414, x15415, x15416;
  wire x15417, x15418, x15419, x15420, x15421, x15422, x15423, x15424;
  wire x15425, x15426, x15427, x15428, x15429, x15430, x15431, x15432;
  wire x15433, x15434, x15435, x15436, x15437, x15438, x15439, x15440;
  wire x15446, x15450, x15454, x15458, x15462, x15466, x15470, x15474;
  wire x15478, x15482, x15486, x15490, x15494, x15498, x15502, x15506;
  wire x15510, x15514, x15518, x15522, x15526, x15530, x15534, x15538;
  wire x15542, x15546, x15550, x15554, x15558, x15559, x15561, x15564;
  wire x15567, x15570, x15572, x15575, x15577, x15580, x15582, x15585;
  wire x15587, x15590, x15592, x15595, x15597, x15600, x15602, x15605;
  wire x15607, x15610, x15612, x15615, x15617, x15620, x15622, x15625;
  wire x15627, x15630, x15632, x15635, x15637, x15640, x15642, x15645;
  wire x15647, x15650, x15652, x15655, x15657, x15660, x15662, x15665;
  wire x15667, x15670, x15672, x15675, x15677, x15680, x15682, x15685;
  wire x15687, x15690, x15692, x15695, x15697, x15700, x15701, x15703;
  wire x15706, x15709, x15712, x15715, x15718, x15720, x15723, x15725;
  wire x15728, x15730, x15733, x15735, x15738, x15740, x15743, x15745;
  wire x15748, x15750, x15753, x15755, x15758, x15760, x15763, x15765;
  wire x15768, x15770, x15773, x15775, x15778, x15780, x15783, x15785;
  wire x15788, x15790, x15793, x15795, x15798, x15800, x15803, x15805;
  wire x15808, x15810, x15813, x15815, x15818, x15820, x15823, x15825;
  wire x15828, x15829, x15831, x15834, x15837, x15840, x15843, x15846;
  wire x15849, x15852, x15855, x15858, x15860, x15863, x15865, x15868;
  wire x15870, x15873, x15875, x15878, x15880, x15883, x15885, x15888;
  wire x15890, x15893, x15895, x15898, x15900, x15903, x15905, x15908;
  wire x15910, x15913, x15915, x15918, x15920, x15923, x15925, x15928;
  wire x15929, x15931, x15934, x15937, x15940, x15943, x15946, x15949;
  wire x15952, x15955, x15958, x15961, x15964, x15967, x15970, x15973;
  wire x15980, x15982, x15989, x15993, x15997, x16004, x16008, x16012;
  wire x16016, x16020, x16024, x16028, x16035, x16039, x16043, x16047;
  wire x16051, x16055, x16059, x16063, x16067, x16071, x16075, x16079;
  wire x16083, x16087, x16091, x16096, x16098, x16100, x16102, x16104;
  wire x16106, x16108, x16110, x16112, x16114, x16116, x16118, x16120;
  wire x16122, x16124, x16126, x16128, x16130, x16132, x16134, x16136;
  wire x16138, x16140, x16142, x16144, x16146, x16148, x16152, x16154;
  wire x16156, x16158, x16160, x16162, x16164, x16166, x16168, x16170;
  wire x16172, x16174, x16176, x16178, x16180, x16182, x16184, x16186;
  wire x16188, x16190, x16192, x16194, x16196, x16198, x16200, x16206;
  wire x16208, x16210, x16212, x16214, x16216, x16218, x16220, x16222;
  wire x16224, x16226, x16228, x16230, x16232, x16234, x16236, x16238;
  wire x16240, x16242, x16244, x16246, x16256, x16258, x16260, x16262;
  wire x16264, x16266, x16268, x16270, x16272, x16274, x16276, x16278;
  wire x16280, x16296, x16300, x16304, x16308, x16312, x16316, x16320;
  wire x16324, x16328, x16332, x16336, x16340, x16344, x16348, x16352;
  wire x16356, x16360, x16364, x16368, x16372, x16376, x16380, x16384;
  wire x16388, x16392, x16396, x16400, x16404, x16408, x16410, x16508;
  wire x16509, x16512, x16514, x16516, x16518, x16520, x16522, x16524;
  wire x16526, x16528, x16530, x16532, x16534, x16536, x16538, x16540;
  wire x16542, x16544, x16546, x16548, x16550, x16552, x16554, x16556;
  wire x16558, x16560, x16562, x16564, x16566, x16568, x16570, x16572;
  wire x16574, x16576, x16578, x16580, x16582, x16584, x16586, x16588;
  wire x16590, x16592, x16594, x16596, x16598, x16600, x16602, x16604;
  wire x16606, x16608, x16610, x16612, x16658, x16659, x16661, x16662;
  wire x16664, x16665, x16667, x16679, x16680, x16682, x16683, x16685;
  wire x16686, x16688, x16689, x16691, x16692, x16694, x16695, x16697;
  wire x16698, x16700, x16702, x16703, x16705, x16706, x16709, x16713;
  wire x16714, x16716, x16718, x16719, x16722, x16725, x16726, x16729;
  wire x16732, x16735, x16736, x16738, x16741, x16744, x16745, x16747;
  wire x16843, x16844, x16845, x16846, x16847, x16848, x16849, x16850;
  wire x16851, x16852, x16853, x16854, x16855, x16856, x16857, x16858;
  wire x16859, x16860, x16861, x16862, x16863, x16864, x16865, x16866;
  wire x16867, x16868, x16869, x16870, x16871, x16872, x16873, x16874;
  wire x16876, x16973, x16974, x16977, x16979, x16980, x16983, x16985;
  wire x16986, x16989, x16991, x16992, x16995, x16997, x16998, x17001;
  wire x17003, x17004, x17007, x17009, x17010, x17013, x17015, x17016;
  wire x17019, x17021, x17022, x17025, x17027, x17028, x17031, x17033;
  wire x17034, x17037, x17039, x17040, x17043, x17045, x17046, x17049;
  wire x17051, x17052, x17055, x17057, x17058, x17061, x17063, x17064;
  wire x17067, x17069, x17070, x17073, x17075, x17076, x17079, x17081;
  wire x17082, x17085, x17087, x17088, x17091, x17093, x17094, x17097;
  wire x17099, x17100, x17103, x17105, x17106, x17109, x17111, x17112;
  wire x17115, x17117, x17118, x17121, x17123, x17124, x17127, x17129;
  wire x17130, x17133, x17135, x17136, x17139, x17141, x17142, x17145;
  wire x17147, x17148, x17151, x17153, x17154, x17157, x17159, x17160;
  wire x17163, x17164, x17165, x17166, x17167, x17168, x17169, x17170;
  wire x17171, x17172, x17173, x17174, x17175, x17176, x17177, x17178;
  wire x17179, x17180, x17181, x17182, x17183, x17184, x17185, x17186;
  wire x17187, x17188, x17189, x17190, x17191, x17192, x17193, x17199;
  wire x17203, x17207, x17211, x17215, x17219, x17223, x17227, x17231;
  wire x17235, x17239, x17243, x17247, x17251, x17255, x17259, x17263;
  wire x17267, x17271, x17275, x17279, x17283, x17287, x17291, x17295;
  wire x17299, x17303, x17307, x17311, x17315, x17317, x17320, x17323;
  wire x17326, x17328, x17331, x17333, x17336, x17338, x17341, x17343;
  wire x17346, x17348, x17351, x17353, x17356, x17358, x17361, x17363;
  wire x17366, x17368, x17371, x17373, x17376, x17378, x17381, x17383;
  wire x17386, x17388, x17391, x17393, x17396, x17398, x17401, x17403;
  wire x17406, x17408, x17411, x17413, x17416, x17418, x17421, x17423;
  wire x17426, x17428, x17431, x17433, x17436, x17438, x17441, x17443;
  wire x17446, x17448, x17451, x17453, x17456, x17458, x17461, x17463;
  wire x17466, x17469, x17472, x17475, x17478, x17480, x17483, x17485;
  wire x17488, x17490, x17493, x17495, x17498, x17500, x17503, x17505;
  wire x17508, x17510, x17513, x17515, x17518, x17520, x17523, x17525;
  wire x17528, x17530, x17533, x17535, x17538, x17540, x17543, x17545;
  wire x17548, x17550, x17553, x17555, x17558, x17560, x17563, x17565;
  wire x17568, x17570, x17573, x17575, x17578, x17580, x17583, x17585;
  wire x17588, x17590, x17593, x17595, x17598, x17601, x17604, x17607;
  wire x17610, x17613, x17616, x17619, x17622, x17624, x17627, x17629;
  wire x17632, x17634, x17637, x17639, x17642, x17644, x17647, x17649;
  wire x17652, x17654, x17657, x17659, x17662, x17664, x17667, x17669;
  wire x17672, x17674, x17677, x17679, x17682, x17684, x17687, x17689;
  wire x17692, x17694, x17697, x17699, x17702, x17705, x17708, x17711;
  wire x17714, x17717, x17720, x17723, x17726, x17729, x17732, x17735;
  wire x17738, x17741, x17744, x17748, x17750, x17753, x17755, x17758;
  wire x17760, x17763, x17765, x17768, x17770, x17773, x17775, x17778;
  wire x17780, x17783, x17785, x17788, x17790, x17793, x17795, x17798;
  wire x17800, x17803, x17805, x17808, x17810, x17813, x17815, x17818;
  wire x17820, x17823, x17825, x17828, x17830, x17833, x17835, x17838;
  wire x17840, x17843, x17845, x17848, x17850, x17853, x17855, x17858;
  wire x17860, x17863, x17865, x17868, x17870, x17873, x17875, x17878;
  wire x17880, x17883, x17885, x17888, x17890, x17893, x17895, x17898;
  wire x17900, x17903, x17906, x17908, x17910, x17912, x17914, x17916;
  wire x17918, x17920, x17923, x17925, x17927, x17929, x17931, x17933;
  wire x17935, x17937, x17939, x17941, x17943, x17945, x17947, x17949;
  wire x17951, x17953, x17955, x17958, x17960, x17962, x17964, x17966;
  wire x17968, x17970, x17972, x17974, x17976, x17978, x17980, x17982;
  wire x17984, x17986, x17988, x17990, x17992, x17994, x17996, x17998;
  wire x18000, x18002, x18004, x18006, x18008, x18011, x18013, x18015;
  wire x18017, x18019, x18021, x18023, x18025, x18027, x18029, x18031;
  wire x18033, x18035, x18037, x18039, x18041, x18043, x18045, x18047;
  wire x18049, x18051, x18053, x18055, x18057, x18059, x18061, x18063;
  wire x18065, x18067, x18069, x18071, x18073, x18075, x18077, x18079;
  wire x18082, x18084, x18086, x18088, x18090, x18092, x18094, x18096;
  wire x18098, x18100, x18102, x18104, x18106, x18108, x18110, x18112;
  wire x18114, x18116, x18118, x18120, x18122, x18124, x18126, x18128;
  wire x18130, x18132, x18134, x18136, x18138, x18140, x18142, x18144;
  wire x18146, x18148, x18150, x18152, x18154, x18156, x18158, x18160;
  wire x18162, x18164, x18166, x18168, x18171, x18173, x18175, x18177;
  wire x18179, x18181, x18183, x18185, x18187, x18189, x18191, x18193;
  wire x18195, x18197, x18199, x18201, x18203, x18205, x18207, x18209;
  wire x18211, x18213, x18215, x18217, x18219, x18221, x18223, x18225;
  wire x18227, x18229, x18231, x18233, x18235, x18237, x18239, x18241;
  wire x18243, x18245, x18247, x18249, x18251, x18253, x18255, x18257;
  wire x18259, x18261, x18263, x18265, x18267, x18269, x18271, x18273;
  wire x18275, x18278, x18280, x18282, x18284, x18286, x18288, x18290;
  wire x18292, x18294, x18296, x18298, x18300, x18302, x18304, x18306;
  wire x18308, x18310, x18312, x18314, x18316, x18318, x18320, x18322;
  wire x18324, x18326, x18328, x18330, x18332, x18334, x18336, x18338;
  wire x18340, x18342, x18344, x18346, x18348, x18350, x18352, x18354;
  wire x18356, x18358, x18360, x18362, x18364, x18366, x18368, x18370;
  wire x18372, x18374, x18376, x18378, x18380, x18382, x18384, x18386;
  wire x18388, x18390, x18392, x18394, x18396, x18398, x18400, x18403;
  wire x18405, x18407, x18409, x18411, x18413, x18415, x18417, x18419;
  wire x18421, x18423, x18425, x18427, x18429, x18431, x18433, x18435;
  wire x18437, x18439, x18441, x18443, x18445, x18447, x18449, x18451;
  wire x18453, x18455, x18457, x18459, x18461, x18463, x18465, x18467;
  wire x18469, x18471, x18473, x18475, x18477, x18479, x18481, x18483;
  wire x18485, x18487, x18489, x18491, x18493, x18495, x18497, x18499;
  wire x18501, x18503, x18505, x18507, x18509, x18511, x18513, x18515;
  wire x18517, x18519, x18521, x18523, x18525, x18527, x18529, x18531;
  wire x18533, x18535, x18537, x18539, x18541, x18543, x18546, x18548;
  wire x18550, x18552, x18554, x18556, x18558, x18560, x18562, x18564;
  wire x18566, x18568, x18570, x18572, x18574, x18576, x18578, x18580;
  wire x18582, x18584, x18586, x18588, x18590, x18592, x18594, x18596;
  wire x18598, x18600, x18602, x18604, x18606, x18608, x18610, x18612;
  wire x18614, x18616, x18618, x18620, x18622, x18624, x18626, x18628;
  wire x18630, x18632, x18634, x18636, x18638, x18640, x18642, x18644;
  wire x18646, x18648, x18650, x18652, x18654, x18656, x18658, x18660;
  wire x18662, x18664, x18666, x18668, x18670, x18672, x18674, x18676;
  wire x18678, x18680, x18682, x18684, x18686, x18688, x18690, x18692;
  wire x18694, x18696, x18698, x18700, x18702, x18704, x18707, x18709;
  wire x18711, x18713, x18715, x18717, x18719, x18721, x18723, x18725;
  wire x18727, x18729, x18731, x18733, x18735, x18737, x18739, x18741;
  wire x18743, x18745, x18747, x18749, x18751, x18753, x18755, x18757;
  wire x18759, x18761, x18763, x18765, x18767, x18769, x18771, x18773;
  wire x18775, x18777, x18779, x18781, x18783, x18785, x18787, x18789;
  wire x18791, x18793, x18795, x18797, x18799, x18801, x18803, x18805;
  wire x18807, x18809, x18811, x18813, x18815, x18817, x18819, x18821;
  wire x18823, x18825, x18827, x18829, x18831, x18833, x18835, x18837;
  wire x18839, x18841, x18843, x18845, x18847, x18849, x18851, x18853;
  wire x18855, x18857, x18859, x18861, x18863, x18865, x18867, x18869;
  wire x18871, x18873, x18875, x18877, x18879, x18881, x18883, x18886;
  wire x18888, x18890, x18892, x18894, x18896, x18898, x18900, x18902;
  wire x18904, x18906, x18908, x18910, x18912, x18914, x18916, x18918;
  wire x18920, x18922, x18924, x18926, x18928, x18930, x18932, x18934;
  wire x18936, x18938, x18940, x18942, x18944, x18946, x18948, x18955;
  wire x18963, x18971, x18982, x18990, x18998, x19006, x19010, x19015;
  wire x19023, x19027, x19035, x19043, x19047, x19052, x19056, x19061;
  wire x19069, x19073, x19078, x19082, x19087, x19095, x19099, x19104;
  wire x19108, x19116, x19124, x19128, x19133, x19137, x19142, x19146;
  wire x19151, x19159, x19163, x19168, x19172, x19177, x19181, x19186;
  wire x19194, x19198, x19203, x19207, x19212, x19216, x19224, x19232;
  wire x19236, x19241, x19245, x19250, x19254, x19259, x19267, x19275;
  wire x19279, x19284, x19288, x19293, x19297, x19302, x19306, x19311;
  wire x19319, x19323, x19328, x19332, x19337, x19341, x19346, x19350;
  wire x19358, x19366, x19370, x19375, x19379, x19384, x19388, x19393;
  wire x19397, x19402, x19406, x19411, x19419, x19423, x19428, x19432;
  wire x19437, x19441, x19446, x19450, x19455, x19459, x19464, x19472;
  wire x19476, x19481, x19485, x19490, x19494, x19499, x19503, x19508;
  wire x19512, x19520, x19528, x19532, x19537, x19541, x19546, x19550;
  wire x19555, x19559, x19564, x19568, x19573, x19577, x19582, x19590;
  wire x19594, x19599, x19603, x19608, x19612, x19617, x19621, x19626;
  wire x19630, x19635, x19639, x19644, x19652, x19656, x19661, x19665;
  wire x19670, x19674, x19679, x19683, x19688, x19692, x19697, x19701;
  wire x19709, x19717, x19721, x19726, x19730, x19735, x19739, x19744;
  wire x19748, x19753, x19757, x19762, x19766, x19771, x19779, x19787;
  wire x19791, x19796, x19800, x19805, x19809, x19814, x19818, x19823;
  wire x19827, x19832, x19836, x19841, x19845, x19850, x19858, x19862;
  wire x19867, x19871, x19876, x19880, x19885, x19889, x19894, x19898;
  wire x19903, x19907, x19912, x19916, x19924, x19932, x19936, x19941;
  wire x19945, x19950, x19954, x19959, x19963, x19968, x19972, x19977;
  wire x19981, x19986, x19990, x19995, x19999, x20004, x20012, x20016;
  wire x20021, x20025, x20030, x20034, x20039, x20043, x20048, x20052;
  wire x20057, x20061, x20066, x20070, x20075, x20079, x20084, x20092;
  wire x20096, x20101, x20105, x20110, x20114, x20119, x20123, x20128;
  wire x20132, x20137, x20141, x20146, x20150, x20155, x20159, x20167;
  wire x20171, x20176, x20180, x20185, x20189, x20194, x20198, x20203;
  wire x20207, x20212, x20216, x20221, x20225, x20230, x20234, x20239;
  wire x20243, x20248, x20252, x20257, x20261, x20266, x20270, x20275;
  wire x20279, x20284, x20288, x20293, x20297, x20302, x20306, x20311;
  wire x20315, x20320, x20324, x20329, x20333, x20338, x20342, x20347;
  wire x20351, x20355, x20359, x20363, x20367, x20371, x20375, x20379;
  wire x20383, x20387, x20391, x20395, x20399, x20403, x20407, x20411;
  wire x20415, x20419, x20423, x20427, x20428, x20429, x20431, x20435;
  wire x20436, x20443, x20444, x20451, x20452, x20455, x20464, x20465;
  wire x20468, x20470, x20477, x20481, x20484, x20485, x20488, x20490;
  wire x20497, x20501, x20504, x20505, x20508, x20510, x20517, x20521;
  wire x20524, x20525, x20528, x20530, x20534, x20538, x20542, x20545;
  wire x20546, x20549, x20551, x20555, x20559, x20563, x20566, x20567;
  wire x20570, x20572, x20577, x20583, x20587, x20590, x20591, x20594;
  wire x20596, x20601, x20602, x20608, x20612, x20618, x20619, x20622;
  wire x20624, x20629, x20630, x20636, x20640, x20646, x20647, x20650;
  wire x20652, x20657, x20658, x20661, x20665, x20670, x20674, x20680;
  wire x20681, x20684, x20686, x20691, x20692, x20695, x20697, x20700;
  wire x20705, x20709, x20714, x20720, x20721, x20724, x20726, x20731;
  wire x20732, x20735, x20737, x20740, x20745, x20749, x20754, x20760;
  wire x20761, x20764, x20766, x20771, x20772, x20775, x20777, x20780;
  wire x20785, x20789, x20794, x20800, x20801, x20804, x20806, x20811;
  wire x20812, x20815, x20817, x20820, x20822, x20826, x20830, x20835;
  wire x20839, x20842, x20843, x20846, x20848, x20853, x20854, x20857;
  wire x20859, x20862, x20864, x20868, x20872, x20877, x20881, x20884;
  wire x20885, x20888, x20890, x20895, x20896, x20899, x20901, x20904;
  wire x20907, x20913, x20917, x20922, x20926, x20929, x20930, x20933;
  wire x20935, x20940, x20941, x20944, x20946, x20949, x20952, x20953;
  wire x20959, x20963, x20968, x20972, x20978, x20979, x20982, x20984;
  wire x20987, x20990, x20991, x20994, x20996, x20999, x21002, x21003;
  wire x21009, x21013, x21018, x21022, x21028, x21029, x21032, x21034;
  wire x21037, x21040, x21041, x21044, x21046, x21049, x21052, x21053;
  wire x21056, x21060, x21065, x21069, x21074, x21078, x21084, x21085;
  wire x21088, x21090, x21093, x21096, x21097, x21100, x21102, x21105;
  wire x21108, x21109, x21112, x21114, x21117, x21122, x21126, x21131;
  wire x21135, x21140, x21144, x21147, x21148, x21151, x21153, x21156;
  wire x21159, x21160, x21163, x21165, x21168, x21171, x21172, x21175;
  wire x21177, x21180, x21185, x21189, x21194, x21198, x21203, x21207;
  wire x21210, x21211, x21214, x21216, x21219, x21222, x21223, x21226;
  wire x21228, x21231, x21234, x21235, x21238, x21240, x21243, x21248;
  wire x21252, x21256, x21261, x21265, x21270, x21274, x21277, x21278;
  wire x21281, x21283, x21286, x21289, x21290, x21293, x21295, x21298;
  wire x21301, x21302, x21305, x21307, x21310, x21312, x21316, x21320;
  wire x21324, x21329, x21333, x21338, x21342, x21345, x21346, x21349;
  wire x21351, x21354, x21356, x21357, x21360, x21362, x21365, x21367;
  wire x21368, x21371, x21373, x21376, x21377, x21381, x21385, x21389;
  wire x21393, x21397, x21401, x21405, x21409, x21413, x21417, x21421;
  wire x21425, x21429, x21430, x21434, x21435, x21436, x21440, x21441;
  wire x21442, x21446, x21450, x21451, x21452, x21456, x21460, x21461;
  wire x21462, x21466, x21470, x21471, x21472, x21476, x21480, x21482;
  wire x21485, x21489, x21493, x21495, x21498, x21502, x21506, x21510;
  wire x21512, x21515, x21519, x21523, x21527, x21529, x21530, x21533;
  wire x21537, x21541, x21545, x21547, x21548, x21551, x21553, x21556;
  wire x21560, x21564, x21566, x21567, x21570, x21572, x21575, x21579;
  wire x21583, x21587, x21590, x21591, x21594, x21596, x21599, x21603;
  wire x21607, x21611, x21617, x21618, x21621, x21623, x21626, x21630;
  wire x21634, x21638, x21644, x21645, x21648, x21650, x21653, x21657;
  wire x21661, x21665, x21671, x21672, x21675, x21679, x21681, x21683;
  wire x21686, x21690, x21694, x21698, x21704, x21705, x21708, x21712;
  wire x21714, x21716, x21719, x21723, x21727, x21732, x21736, x21742;
  wire x21743, x21746, x21750, x21752, x21754, x21757, x21761, x21765;
  wire x21770, x21774, x21780, x21781, x21784, x21786, x21789, x21791;
  wire x21793, x21796, x21800, x21804, x21809, x21813, x21819, x21820;
  wire x21823, x21825, x21828, x21830, x21832, x21835, x21837, x21840;
  wire x21844, x21849, x21853, x21859, x21860, x21863, x21865, x21868;
  wire x21870, x21872, x21875, x21877, x21880, x21884, x21889, x21893;
  wire x21899, x21900, x21903, x21905, x21908, x21911, x21914, x21916;
  wire x21919, x21922, x21925, x21929, x21934, x21938, x21943, x21947;
  wire x21950, x21951, x21954, x21956, x21959, x21961, x21964, x21966;
  wire x21969, x21971, x21974, x21978, x21982, x21986, x21990, x21994;
  wire x22004, x22008, x22015, x22022, x22026, x22034, x22038, x22046;
  wire x22050, x22058, x22062, x22070, x22074, x22079, x22083, x22087;
  wire x22092, x22096, x22100, x22105, x22109, x22113, x22118, x22122;
  wire x22126, x22131, x22135, x22139, x22143, x22148, x22152, x22157;
  wire x22161, x22165, x22170, x22174, x22179, x22183, x22187, x22192;
  wire x22196, x22201, x22205, x22209, x22214, x22218, x22223, x22227;
  wire x22231, x22236, x22240, x22242, x22246, x22250, x22254, x22259;
  wire x22263, x22266, x22269, x22273, x22278, x22282, x22287, x22291;
  wire x22294, x22297, x22301, x22306, x22310, x22315, x22319, x22322;
  wire x22325, x22329, x22334, x22338, x22341, x22344, x22348, x22351;
  wire x22354, x22358, x22363, x22367, x22370, x22373, x22375, x22378;
  wire x22381, x22384, x22388, x22393, x22397, x22400, x22403, x22405;
  wire x22408, x22411, x22414, x22418, x22423, x22427, x22430, x22433;
  wire x22435, x22438, x22441, x22444, x22448, x22453, x22457, x22460;
  wire x22463, x22465, x22468, x22471, x22474, x22478, x22483, x22487;
  wire x22490, x22493, x22495, x22498, x22501, x22504, x22508, x22513;
  wire x22517, x22520, x22521, x22524, x22526, x22529, x22531, x22532;
  wire x22535, x22539, x22543, x22547, x22560, x22565, x22568, x22573;
  wire x22576, x22581, x22584, x22589, x22592, x22597, x22600, x22604;
  wire x22608, x22611, x22614, x22618, x22622, x22625, x22628, x22632;
  wire x22636, x22639, x22642, x22646, x22650, x22653, x22656, x22660;
  wire x22664, x22669, x22671, x22674, x22679, x22683, x22686, x22689;
  wire x22691, x22694, x22699, x22703, x22706, x22709, x22711, x22714;
  wire x22719, x22723, x22726, x22729, x22731, x22734, x22739, x22743;
  wire x22746, x22749, x22751, x22754, x22759, x22763, x22766, x22769;
  wire x22771, x22774, x22779, x22783, x22786, x22787, x22790, x22792;
  wire x22795, x22800, x22804, x22807, x22808, x22811, x22813, x22816;
  wire x22821, x22825, x22828, x22829, x22832, x22834, x22837, x22842;
  wire x22846, x22849, x22850, x22853, x22855, x22858, x22863, x22867;
  wire x22870, x22871, x22874, x22876, x22879, x22884, x22888, x22891;
  wire x22892, x22895, x22897, x22900, x22905, x22909, x22912, x22913;
  wire x22916, x22918, x22921, x22926, x22930, x22933, x22934, x22937;
  wire x22939, x22942, x22947, x22951, x22954, x22955, x22958, x22960;
  wire x22963, x22967, x22971, x22978, x22982, x22986, x22990, x22995;
  wire x22999, x23004, x23008, x23013, x23017, x23022, x23026, x23031;
  wire x23032, x23034, x23037, x23041, x23046, x23047, x23049, x23052;
  wire x23056, x23061, x23062, x23064, x23067, x23071, x23076, x23077;
  wire x23079, x23082, x23086, x23091, x23092, x23094, x23097, x23101;
  wire x23106, x23107, x23109, x23110, x23113, x23117, x23122, x23123;
  wire x23125, x23126, x23129, x23133, x23138, x23139, x23141, x23142;
  wire x23145, x23149, x23154, x23155, x23157, x23158, x23161, x23165;
  wire x23170, x23171, x23173, x23174, x23177, x23181, x23186, x23187;
  wire x23189, x23190, x23193, x23197, x23202, x23203, x23205, x23206;
  wire x23209, x23213, x23218, x23219, x23221, x23222, x23225, x23229;
  wire x23234, x23235, x23237, x23238, x23241, x23245, x23250, x23251;
  wire x23253, x23254, x23257, x23261, x23266, x23267, x23269, x23270;
  wire x23273, x23277, x23282, x23283, x23285, x23286, x23289, x23293;
  wire x23298, x23299, x23301, x23302, x23305, x23309, x23314, x23315;
  wire x23317, x23318, x23321, x23325, x23329, x23339, x23343, x23344;
  wire x23348, x23349, x23353, x23354, x23358, x23359, x23363, x23365;
  wire x23368, x23372, x23375, x23378, x23382, x23385, x23388, x23392;
  wire x23395, x23398, x23402, x23405, x23408, x23412, x23415, x23418;
  wire x23422, x23425, x23428, x23432, x23435, x23438, x23442, x23445;
  wire x23448, x23452, x23455, x23458, x23462, x23465, x23468, x23472;
  wire x23475, x23478, x23482, x23485, x23488, x23492, x23495, x23498;
  wire x23502, x23505, x23508, x23512, x23515, x23518, x23522, x23525;
  wire x23528, x23532, x23535, x23538, x23542, x23545, x23548, x23552;
  wire x23556, x23564, x23568, x23572, x23576, x23581, x23585, x23590;
  wire x23594, x23599, x23603, x23608, x23612, x23617, x23621, x23626;
  wire x23630, x23633, x23636, x23640, x23643, x23646, x23650, x23653;
  wire x23656, x23660, x23663, x23666, x23670, x23673, x23676, x23680;
  wire x23683, x23686, x23690, x23693, x23696, x23700, x23703, x23706;
  wire x23710, x23713, x23716, x23720, x23723, x23726, x23730, x23733;
  wire x23736, x23740, x23743, x23746, x23750, x23753, x23756, x23760;
  wire x23763, x23766, x23770, x23773, x23776, x23780, x23783, x23786;
  wire x23790, x23793, x23796, x23800, x23803, x23806, x23810, x23812;
  wire x23818, x23822, x23824, x23827, x23829, x23832, x23834, x23837;
  wire x23839, x23842, x23844, x23847, x23849, x23852, x23854, x23857;
  wire x23859, x23862, x23864, x23867, x23869, x23872, x23874, x23877;
  wire x23879, x23882, x23884, x23887, x23889, x23892, x23894, x23897;
  wire x23899, x23902, x23904, x23907, x23909, x23912, x23914, x23917;
  wire x23919, x23922, x23924, x23927, x23929, x23932, x23934, x23937;
  wire x23939, x23942, x23943, x23944, x23945, x23946, x23947, x23948;
  wire x23949, x23950, x23951, x23952, x23953, x23954, x23955, x23956;
  wire x23957, x23958, x23959, x23960, x23961, x23962, x23963, x23964;
  wire x23965, x23966, x23967, x23973, x23977, x23981, x23985, x23989;
  wire x23993, x23997, x24001, x24005, x24009, x24013, x24017, x24021;
  wire x24025, x24029, x24033, x24037, x24041, x24045, x24049, x24053;
  wire x24057, x24061, x24065, x24066, x24068, x24071, x24074, x24077;
  wire x24079, x24082, x24084, x24087, x24089, x24092, x24094, x24097;
  wire x24099, x24102, x24104, x24107, x24109, x24112, x24114, x24117;
  wire x24119, x24122, x24124, x24127, x24129, x24132, x24134, x24137;
  wire x24139, x24142, x24144, x24147, x24149, x24152, x24154, x24157;
  wire x24159, x24162, x24164, x24167, x24169, x24172, x24174, x24177;
  wire x24179, x24182, x24183, x24184, x24186, x24189, x24192, x24195;
  wire x24198, x24201, x24203, x24206, x24208, x24211, x24213, x24216;
  wire x24218, x24221, x24223, x24226, x24228, x24231, x24233, x24236;
  wire x24238, x24241, x24243, x24246, x24248, x24251, x24253, x24256;
  wire x24258, x24261, x24263, x24266, x24268, x24271, x24273, x24276;
  wire x24278, x24281, x24283, x24286, x24287, x24288, x24289, x24290;
  wire x24292, x24295, x24298, x24301, x24304, x24307, x24310, x24313;
  wire x24316, x24319, x24321, x24324, x24326, x24329, x24331, x24334;
  wire x24336, x24339, x24341, x24344, x24346, x24349, x24351, x24354;
  wire x24356, x24359, x24361, x24364, x24365, x24366, x24367, x24368;
  wire x24369, x24370, x24372, x24375, x24378, x24381, x24384, x24387;
  wire x24390, x24393, x24396, x24399, x24403, x24407, x24411, x24415;
  wire x24419, x24423, x24427, x24431, x24433, x24436, x24438, x24441;
  wire x24445, x24449, x24453, x24457, x24461, x24465, x24467, x24470;
  wire x24472, x24475, x24477, x24480, x24482, x24485, x24487, x24490;
  wire x24492, x24495, x24497, x24500, x24502, x24505, x24507, x24510;
  wire x24512, x24515, x24517, x24519, x24521, x24523, x24525, x24527;
  wire x24529, x24531, x24533, x24535, x24537, x24539, x24541, x24543;
  wire x24545, x24547, x24549, x24551, x24553, x24555, x24557, x24559;
  wire x24561, x24563, x24565, x24567, x24569, x24571, x24573, x24575;
  wire x24578, x24580, x24582, x24584, x24586, x24588, x24590, x24592;
  wire x24594, x24596, x24598, x24600, x24602, x24604, x24606, x24608;
  wire x24610, x24612, x24614, x24616, x24618, x24620, x24622, x24624;
  wire x24626, x24628, x24630, x24632, x24637, x24639, x24641, x24643;
  wire x24645, x24647, x24649, x24651, x24653, x24655, x24657, x24659;
  wire x24661, x24663, x24665, x24667, x24669, x24671, x24673, x24675;
  wire x24677, x24679, x24681, x24683, x24693, x24695, x24697, x24699;
  wire x24701, x24703, x24705, x24707, x24709, x24711, x24713, x24715;
  wire x24717, x24719, x24721, x24739, x24743, x24747, x24751, x24755;
  wire x24759, x24763, x24767, x24771, x24775, x24779, x24783, x24787;
  wire x24791, x24795, x24799, x24803, x24807, x24811, x24815, x24819;
  wire x24823, x24827, x24831, x24835, x24839, x24843, x24847, x24851;
  wire x24855, x24859, x24860, x24862, x24864, x24866, x24868, x24870;
  wire x24872, x24874, x24876, x24878, x24880, x24882, x24884, x24886;
  wire x24888, x24890, x24892, x24926, x24928, x24930, x24932, x24934;
  wire x24936, x24938, x24940, x24942, x24944, x24946, x24948, x24950;
  wire x24952, x24954, x24956, x24958, x24960, x24962, x24964, x24966;
  wire x24968, x24970, x24972, x24974, x24976, x24978, x24980, x24982;
  wire x24984, x24986, x24988, x25749, x25772, x25782, x25790, x25796;
  wire x27944, x27945, x27946, x27947, x27948, x27949, x27950, x27951;
  wire x27952, x27953, x27954, x27955, x27956, x27957, x27958, x27959;
  wire x27960, x27961, x27962, x27963, x27964, x27965, x27966, x27967;
  wire x27968, x27969, x27970, x27971, x27972, x27973, x27974, x27975;
  wire x28073, x28074, x28077, x28079, x28080, x28083, x28085, x28086;
  wire x28089, x28091, x28092, x28095, x28097, x28098, x28101, x28103;
  wire x28104, x28107, x28109, x28110, x28113, x28115, x28116, x28119;
  wire x28121, x28122, x28125, x28127, x28128, x28131, x28133, x28134;
  wire x28137, x28139, x28140, x28143, x28145, x28146, x28149, x28151;
  wire x28152, x28155, x28157, x28158, x28161, x28163, x28164, x28167;
  wire x28169, x28170, x28173, x28175, x28176, x28179, x28181, x28182;
  wire x28185, x28187, x28188, x28191, x28193, x28194, x28197, x28199;
  wire x28200, x28203, x28205, x28206, x28209, x28211, x28212, x28215;
  wire x28217, x28218, x28221, x28223, x28224, x28227, x28229, x28230;
  wire x28233, x28235, x28236, x28239, x28241, x28242, x28245, x28247;
  wire x28248, x28251, x28253, x28254, x28257, x28259, x28260, x28263;
  wire x28264, x28265, x28266, x28267, x28268, x28269, x28270, x28271;
  wire x28272, x28273, x28274, x28275, x28276, x28277, x28278, x28279;
  wire x28280, x28281, x28282, x28283, x28284, x28285, x28286, x28287;
  wire x28288, x28289, x28290, x28291, x28292, x28293, x28299, x28303;
  wire x28307, x28311, x28315, x28319, x28323, x28327, x28331, x28335;
  wire x28339, x28343, x28347, x28351, x28355, x28359, x28363, x28367;
  wire x28371, x28375, x28379, x28383, x28387, x28391, x28395, x28399;
  wire x28403, x28407, x28411, x28415, x28417, x28420, x28423, x28426;
  wire x28428, x28431, x28433, x28436, x28438, x28441, x28443, x28446;
  wire x28448, x28451, x28453, x28456, x28458, x28461, x28463, x28466;
  wire x28468, x28471, x28473, x28476, x28478, x28481, x28483, x28486;
  wire x28488, x28491, x28493, x28496, x28498, x28501, x28503, x28506;
  wire x28508, x28511, x28513, x28516, x28518, x28521, x28523, x28526;
  wire x28528, x28531, x28533, x28536, x28538, x28541, x28543, x28546;
  wire x28548, x28551, x28553, x28556, x28558, x28561, x28563, x28566;
  wire x28569, x28572, x28575, x28578, x28580, x28583, x28585, x28588;
  wire x28590, x28593, x28595, x28598, x28600, x28603, x28605, x28608;
  wire x28610, x28613, x28615, x28618, x28620, x28623, x28625, x28628;
  wire x28630, x28633, x28635, x28638, x28640, x28643, x28645, x28648;
  wire x28650, x28653, x28655, x28658, x28660, x28663, x28665, x28668;
  wire x28670, x28673, x28675, x28678, x28680, x28683, x28685, x28688;
  wire x28690, x28693, x28695, x28698, x28701, x28704, x28707, x28710;
  wire x28713, x28716, x28719, x28722, x28724, x28727, x28729, x28732;
  wire x28734, x28737, x28739, x28742, x28744, x28747, x28749, x28752;
  wire x28754, x28757, x28759, x28762, x28764, x28767, x28769, x28772;
  wire x28774, x28777, x28779, x28782, x28784, x28787, x28789, x28792;
  wire x28794, x28797, x28799, x28802, x28805, x28808, x28811, x28814;
  wire x28817, x28820, x28823, x28826, x28829, x28832, x28835, x28838;
  wire x28841, x28844, x28848, x28850, x28853, x28855, x28858, x28860;
  wire x28863, x28865, x28868, x28870, x28873, x28875, x28878, x28880;
  wire x28883, x28885, x28888, x28890, x28893, x28895, x28898, x28900;
  wire x28903, x28905, x28908, x28910, x28913, x28915, x28918, x28920;
  wire x28923, x28925, x28928, x28930, x28933, x28935, x28938, x28940;
  wire x28943, x28945, x28948, x28950, x28953, x28955, x28958, x28960;
  wire x28963, x28965, x28968, x28970, x28973, x28975, x28978, x28980;
  wire x28983, x28985, x28988, x28990, x28993, x28995, x28998, x29000;
  wire x29003, x29006, x29008, x29010, x29012, x29014, x29016, x29018;
  wire x29020, x29023, x29025, x29027, x29029, x29031, x29033, x29035;
  wire x29037, x29039, x29041, x29043, x29045, x29047, x29049, x29051;
  wire x29053, x29055, x29058, x29060, x29062, x29064, x29066, x29068;
  wire x29070, x29072, x29074, x29076, x29078, x29080, x29082, x29084;
  wire x29086, x29088, x29090, x29092, x29094, x29096, x29098, x29100;
  wire x29102, x29104, x29106, x29108, x29111, x29113, x29115, x29117;
  wire x29119, x29121, x29123, x29125, x29127, x29129, x29131, x29133;
  wire x29135, x29137, x29139, x29141, x29143, x29145, x29147, x29149;
  wire x29151, x29153, x29155, x29157, x29159, x29161, x29163, x29165;
  wire x29167, x29169, x29171, x29173, x29175, x29177, x29179, x29182;
  wire x29184, x29186, x29188, x29190, x29192, x29194, x29196, x29198;
  wire x29200, x29202, x29204, x29206, x29208, x29210, x29212, x29214;
  wire x29216, x29218, x29220, x29222, x29224, x29226, x29228, x29230;
  wire x29232, x29234, x29236, x29238, x29240, x29242, x29244, x29246;
  wire x29248, x29250, x29252, x29254, x29256, x29258, x29260, x29262;
  wire x29264, x29266, x29268, x29271, x29273, x29275, x29277, x29279;
  wire x29281, x29283, x29285, x29287, x29289, x29291, x29293, x29295;
  wire x29297, x29299, x29301, x29303, x29305, x29307, x29309, x29311;
  wire x29313, x29315, x29317, x29319, x29321, x29323, x29325, x29327;
  wire x29329, x29331, x29333, x29335, x29337, x29339, x29341, x29343;
  wire x29345, x29347, x29349, x29351, x29353, x29355, x29357, x29359;
  wire x29361, x29363, x29365, x29367, x29369, x29371, x29373, x29375;
  wire x29378, x29380, x29382, x29384, x29386, x29388, x29390, x29392;
  wire x29394, x29396, x29398, x29400, x29402, x29404, x29406, x29408;
  wire x29410, x29412, x29414, x29416, x29418, x29420, x29422, x29424;
  wire x29426, x29428, x29430, x29432, x29434, x29436, x29438, x29440;
  wire x29442, x29444, x29446, x29448, x29450, x29452, x29454, x29456;
  wire x29458, x29460, x29462, x29464, x29466, x29468, x29470, x29472;
  wire x29474, x29476, x29478, x29480, x29482, x29484, x29486, x29488;
  wire x29490, x29492, x29494, x29496, x29498, x29500, x29503, x29505;
  wire x29507, x29509, x29511, x29513, x29515, x29517, x29519, x29521;
  wire x29523, x29525, x29527, x29529, x29531, x29533, x29535, x29537;
  wire x29539, x29541, x29543, x29545, x29547, x29549, x29551, x29553;
  wire x29555, x29557, x29559, x29561, x29563, x29565, x29567, x29569;
  wire x29571, x29573, x29575, x29577, x29579, x29581, x29583, x29585;
  wire x29587, x29589, x29591, x29593, x29595, x29597, x29599, x29601;
  wire x29603, x29605, x29607, x29609, x29611, x29613, x29615, x29617;
  wire x29619, x29621, x29623, x29625, x29627, x29629, x29631, x29633;
  wire x29635, x29637, x29639, x29641, x29643, x29646, x29648, x29650;
  wire x29652, x29654, x29656, x29658, x29660, x29662, x29664, x29666;
  wire x29668, x29670, x29672, x29674, x29676, x29678, x29680, x29682;
  wire x29684, x29686, x29688, x29690, x29692, x29694, x29696, x29698;
  wire x29700, x29702, x29704, x29706, x29708, x29710, x29712, x29714;
  wire x29716, x29718, x29720, x29722, x29724, x29726, x29728, x29730;
  wire x29732, x29734, x29736, x29738, x29740, x29742, x29744, x29746;
  wire x29748, x29750, x29752, x29754, x29756, x29758, x29760, x29762;
  wire x29764, x29766, x29768, x29770, x29772, x29774, x29776, x29778;
  wire x29780, x29782, x29784, x29786, x29788, x29790, x29792, x29794;
  wire x29796, x29798, x29800, x29802, x29804, x29807, x29809, x29811;
  wire x29813, x29815, x29817, x29819, x29821, x29823, x29825, x29827;
  wire x29829, x29831, x29833, x29835, x29837, x29839, x29841, x29843;
  wire x29845, x29847, x29849, x29851, x29853, x29855, x29857, x29859;
  wire x29861, x29863, x29865, x29867, x29869, x29871, x29873, x29875;
  wire x29877, x29879, x29881, x29883, x29885, x29887, x29889, x29891;
  wire x29893, x29895, x29897, x29899, x29901, x29903, x29905, x29907;
  wire x29909, x29911, x29913, x29915, x29917, x29919, x29921, x29923;
  wire x29925, x29927, x29929, x29931, x29933, x29935, x29937, x29939;
  wire x29941, x29943, x29945, x29947, x29949, x29951, x29953, x29955;
  wire x29957, x29959, x29961, x29963, x29965, x29967, x29969, x29971;
  wire x29973, x29975, x29977, x29979, x29981, x29983, x29986, x29988;
  wire x29990, x29992, x29994, x29996, x29998, x30000, x30002, x30004;
  wire x30006, x30008, x30010, x30012, x30014, x30016, x30018, x30020;
  wire x30022, x30024, x30026, x30028, x30030, x30032, x30034, x30036;
  wire x30038, x30040, x30042, x30044, x30046, x30048, x30055, x30063;
  wire x30071, x30082, x30090, x30098, x30106, x30110, x30115, x30123;
  wire x30127, x30135, x30143, x30147, x30152, x30156, x30161, x30169;
  wire x30173, x30178, x30182, x30187, x30195, x30199, x30204, x30208;
  wire x30216, x30224, x30228, x30233, x30237, x30242, x30246, x30251;
  wire x30259, x30263, x30268, x30272, x30277, x30281, x30286, x30294;
  wire x30298, x30303, x30307, x30312, x30316, x30324, x30332, x30336;
  wire x30341, x30345, x30350, x30354, x30359, x30367, x30375, x30379;
  wire x30384, x30388, x30393, x30397, x30402, x30406, x30411, x30419;
  wire x30423, x30428, x30432, x30437, x30441, x30446, x30450, x30458;
  wire x30466, x30470, x30475, x30479, x30484, x30488, x30493, x30497;
  wire x30502, x30506, x30511, x30519, x30523, x30528, x30532, x30537;
  wire x30541, x30546, x30550, x30555, x30559, x30564, x30572, x30576;
  wire x30581, x30585, x30590, x30594, x30599, x30603, x30608, x30612;
  wire x30620, x30628, x30632, x30637, x30641, x30646, x30650, x30655;
  wire x30659, x30664, x30668, x30673, x30677, x30682, x30690, x30694;
  wire x30699, x30703, x30708, x30712, x30717, x30721, x30726, x30730;
  wire x30735, x30739, x30744, x30752, x30756, x30761, x30765, x30770;
  wire x30774, x30779, x30783, x30788, x30792, x30797, x30801, x30809;
  wire x30817, x30821, x30826, x30830, x30835, x30839, x30844, x30848;
  wire x30853, x30857, x30862, x30866, x30871, x30879, x30887, x30891;
  wire x30896, x30900, x30905, x30909, x30914, x30918, x30923, x30927;
  wire x30932, x30936, x30941, x30945, x30950, x30958, x30962, x30967;
  wire x30971, x30976, x30980, x30985, x30989, x30994, x30998, x31003;
  wire x31007, x31012, x31016, x31024, x31032, x31036, x31041, x31045;
  wire x31050, x31054, x31059, x31063, x31068, x31072, x31077, x31081;
  wire x31086, x31090, x31095, x31099, x31104, x31112, x31116, x31121;
  wire x31125, x31130, x31134, x31139, x31143, x31148, x31152, x31157;
  wire x31161, x31166, x31170, x31175, x31179, x31184, x31192, x31196;
  wire x31201, x31205, x31210, x31214, x31219, x31223, x31228, x31232;
  wire x31237, x31241, x31246, x31250, x31255, x31259, x31267, x31271;
  wire x31276, x31280, x31285, x31289, x31294, x31298, x31303, x31307;
  wire x31312, x31316, x31321, x31325, x31330, x31334, x31339, x31343;
  wire x31348, x31352, x31357, x31361, x31366, x31370, x31375, x31379;
  wire x31384, x31388, x31393, x31397, x31402, x31406, x31411, x31415;
  wire x31420, x31424, x31429, x31433, x31438, x31442, x31447, x31451;
  wire x31455, x31459, x31463, x31467, x31471, x31475, x31479, x31483;
  wire x31487, x31491, x31495, x31499, x31503, x31507, x31511, x31515;
  wire x31519, x31523, x31527, x31528, x31529, x31531, x31535, x31536;
  wire x31543, x31544, x31551, x31552, x31555, x31564, x31565, x31568;
  wire x31570, x31577, x31581, x31584, x31585, x31588, x31590, x31597;
  wire x31601, x31604, x31605, x31608, x31610, x31617, x31621, x31624;
  wire x31625, x31628, x31630, x31634, x31638, x31642, x31645, x31646;
  wire x31649, x31651, x31655, x31659, x31663, x31666, x31667, x31670;
  wire x31672, x31677, x31683, x31687, x31690, x31691, x31694, x31696;
  wire x31701, x31702, x31708, x31712, x31718, x31719, x31722, x31724;
  wire x31729, x31730, x31736, x31740, x31746, x31747, x31750, x31752;
  wire x31757, x31758, x31761, x31765, x31770, x31774, x31780, x31781;
  wire x31784, x31786, x31791, x31792, x31795, x31797, x31800, x31805;
  wire x31809, x31814, x31820, x31821, x31824, x31826, x31831, x31832;
  wire x31835, x31837, x31840, x31845, x31849, x31854, x31860, x31861;
  wire x31864, x31866, x31871, x31872, x31875, x31877, x31880, x31885;
  wire x31889, x31894, x31900, x31901, x31904, x31906, x31911, x31912;
  wire x31915, x31917, x31920, x31922, x31926, x31930, x31935, x31939;
  wire x31942, x31943, x31946, x31948, x31953, x31954, x31957, x31959;
  wire x31962, x31964, x31968, x31972, x31977, x31981, x31984, x31985;
  wire x31988, x31990, x31995, x31996, x31999, x32001, x32004, x32007;
  wire x32013, x32017, x32022, x32026, x32029, x32030, x32033, x32035;
  wire x32040, x32041, x32044, x32046, x32049, x32052, x32053, x32059;
  wire x32063, x32068, x32072, x32078, x32079, x32082, x32084, x32087;
  wire x32090, x32091, x32094, x32096, x32099, x32102, x32103, x32109;
  wire x32113, x32118, x32122, x32128, x32129, x32132, x32134, x32137;
  wire x32140, x32141, x32144, x32146, x32149, x32152, x32153, x32156;
  wire x32160, x32165, x32169, x32174, x32178, x32184, x32185, x32188;
  wire x32190, x32193, x32196, x32197, x32200, x32202, x32205, x32208;
  wire x32209, x32212, x32214, x32217, x32222, x32226, x32231, x32235;
  wire x32240, x32244, x32247, x32248, x32251, x32253, x32256, x32259;
  wire x32260, x32263, x32265, x32268, x32271, x32272, x32275, x32277;
  wire x32280, x32285, x32289, x32294, x32298, x32303, x32307, x32310;
  wire x32311, x32314, x32316, x32319, x32322, x32323, x32326, x32328;
  wire x32331, x32334, x32335, x32338, x32340, x32343, x32348, x32352;
  wire x32356, x32361, x32365, x32370, x32374, x32377, x32378, x32381;
  wire x32383, x32386, x32389, x32390, x32393, x32395, x32398, x32401;
  wire x32402, x32405, x32407, x32410, x32412, x32416, x32420, x32424;
  wire x32429, x32433, x32438, x32442, x32445, x32446, x32449, x32451;
  wire x32454, x32456, x32457, x32460, x32462, x32465, x32467, x32468;
  wire x32471, x32473, x32476, x32477, x32481, x32485, x32489, x32493;
  wire x32497, x32501, x32505, x32509, x32513, x32517, x32521, x32525;
  wire x32529, x32530, x32534, x32535, x32536, x32540, x32541, x32542;
  wire x32546, x32550, x32551, x32552, x32556, x32560, x32561, x32562;
  wire x32566, x32570, x32571, x32572, x32576, x32580, x32582, x32585;
  wire x32589, x32593, x32595, x32598, x32602, x32606, x32610, x32612;
  wire x32615, x32619, x32623, x32627, x32629, x32630, x32633, x32637;
  wire x32641, x32645, x32647, x32648, x32651, x32653, x32656, x32660;
  wire x32664, x32666, x32667, x32670, x32672, x32675, x32679, x32683;
  wire x32687, x32690, x32691, x32694, x32696, x32699, x32703, x32707;
  wire x32711, x32717, x32718, x32721, x32723, x32726, x32730, x32734;
  wire x32738, x32744, x32745, x32748, x32750, x32753, x32757, x32761;
  wire x32765, x32771, x32772, x32775, x32779, x32781, x32783, x32786;
  wire x32790, x32794, x32798, x32804, x32805, x32808, x32812, x32814;
  wire x32816, x32819, x32823, x32827, x32832, x32836, x32842, x32843;
  wire x32846, x32850, x32852, x32854, x32857, x32861, x32865, x32870;
  wire x32874, x32880, x32881, x32884, x32886, x32889, x32891, x32893;
  wire x32896, x32900, x32904, x32909, x32913, x32919, x32920, x32923;
  wire x32925, x32928, x32930, x32932, x32935, x32937, x32940, x32944;
  wire x32949, x32953, x32959, x32960, x32963, x32965, x32968, x32970;
  wire x32972, x32975, x32977, x32980, x32984, x32989, x32993, x32999;
  wire x33000, x33003, x33005, x33008, x33011, x33014, x33016, x33019;
  wire x33022, x33025, x33029, x33034, x33038, x33043, x33047, x33050;
  wire x33051, x33054, x33056, x33059, x33061, x33064, x33066, x33069;
  wire x33071, x33074, x33078, x33082, x33086, x33090, x33094, x33104;
  wire x33108, x33115, x33122, x33126, x33134, x33138, x33146, x33150;
  wire x33158, x33162, x33170, x33174, x33179, x33183, x33187, x33192;
  wire x33196, x33200, x33205, x33209, x33213, x33218, x33222, x33226;
  wire x33231, x33235, x33239, x33243, x33248, x33252, x33257, x33261;
  wire x33265, x33270, x33274, x33279, x33283, x33287, x33292, x33296;
  wire x33301, x33305, x33309, x33314, x33318, x33323, x33327, x33331;
  wire x33336, x33340, x33342, x33346, x33350, x33354, x33359, x33363;
  wire x33366, x33369, x33373, x33378, x33382, x33387, x33391, x33394;
  wire x33397, x33401, x33406, x33410, x33415, x33419, x33422, x33425;
  wire x33429, x33434, x33438, x33441, x33444, x33448, x33451, x33454;
  wire x33458, x33463, x33467, x33470, x33473, x33475, x33478, x33481;
  wire x33484, x33488, x33493, x33497, x33500, x33503, x33505, x33508;
  wire x33511, x33514, x33518, x33523, x33527, x33530, x33533, x33535;
  wire x33538, x33541, x33544, x33548, x33553, x33557, x33560, x33563;
  wire x33565, x33568, x33571, x33574, x33578, x33583, x33587, x33590;
  wire x33593, x33595, x33598, x33601, x33604, x33608, x33613, x33617;
  wire x33620, x33621, x33624, x33626, x33629, x33631, x33632, x33635;
  wire x33639, x33643, x33647, x33660, x33665, x33668, x33673, x33676;
  wire x33681, x33684, x33689, x33692, x33697, x33700, x33704, x33708;
  wire x33711, x33714, x33718, x33722, x33725, x33728, x33732, x33736;
  wire x33739, x33742, x33746, x33750, x33753, x33756, x33760, x33764;
  wire x33769, x33771, x33774, x33779, x33783, x33786, x33789, x33791;
  wire x33794, x33799, x33803, x33806, x33809, x33811, x33814, x33819;
  wire x33823, x33826, x33829, x33831, x33834, x33839, x33843, x33846;
  wire x33849, x33851, x33854, x33859, x33863, x33866, x33869, x33871;
  wire x33874, x33879, x33883, x33886, x33887, x33890, x33892, x33895;
  wire x33900, x33904, x33907, x33908, x33911, x33913, x33916, x33921;
  wire x33925, x33928, x33929, x33932, x33934, x33937, x33942, x33946;
  wire x33949, x33950, x33953, x33955, x33958, x33963, x33967, x33970;
  wire x33971, x33974, x33976, x33979, x33984, x33988, x33991, x33992;
  wire x33995, x33997, x34000, x34005, x34009, x34012, x34013, x34016;
  wire x34018, x34021, x34026, x34030, x34033, x34034, x34037, x34039;
  wire x34042, x34047, x34051, x34054, x34055, x34058, x34060, x34063;
  wire x34067, x34071, x34078, x34082, x34086, x34090, x34095, x34099;
  wire x34104, x34108, x34113, x34117, x34122, x34126, x34131, x34132;
  wire x34134, x34137, x34141, x34146, x34147, x34149, x34152, x34156;
  wire x34161, x34162, x34164, x34167, x34171, x34176, x34177, x34179;
  wire x34182, x34186, x34191, x34192, x34194, x34197, x34201, x34206;
  wire x34207, x34209, x34210, x34213, x34217, x34222, x34223, x34225;
  wire x34226, x34229, x34233, x34238, x34239, x34241, x34242, x34245;
  wire x34249, x34254, x34255, x34257, x34258, x34261, x34265, x34270;
  wire x34271, x34273, x34274, x34277, x34281, x34286, x34287, x34289;
  wire x34290, x34293, x34297, x34302, x34303, x34305, x34306, x34309;
  wire x34313, x34318, x34319, x34321, x34322, x34325, x34329, x34334;
  wire x34335, x34337, x34338, x34341, x34345, x34350, x34351, x34353;
  wire x34354, x34357, x34361, x34366, x34367, x34369, x34370, x34373;
  wire x34377, x34382, x34383, x34385, x34386, x34389, x34393, x34398;
  wire x34399, x34401, x34402, x34405, x34409, x34414, x34415, x34417;
  wire x34418, x34421, x34425, x34429, x34439, x34443, x34444, x34448;
  wire x34449, x34453, x34454, x34458, x34459, x34463, x34465, x34468;
  wire x34472, x34475, x34478, x34482, x34485, x34488, x34492, x34495;
  wire x34498, x34502, x34505, x34508, x34512, x34515, x34518, x34522;
  wire x34525, x34528, x34532, x34535, x34538, x34542, x34545, x34548;
  wire x34552, x34555, x34558, x34562, x34565, x34568, x34572, x34575;
  wire x34578, x34582, x34585, x34588, x34592, x34595, x34598, x34602;
  wire x34605, x34608, x34612, x34615, x34618, x34622, x34625, x34628;
  wire x34632, x34635, x34638, x34642, x34645, x34648, x34652, x34656;
  wire x34664, x34668, x34672, x34676, x34681, x34685, x34690, x34694;
  wire x34699, x34703, x34708, x34712, x34717, x34721, x34726, x34730;
  wire x34733, x34736, x34740, x34743, x34746, x34750, x34753, x34756;
  wire x34760, x34763, x34766, x34770, x34773, x34776, x34780, x34783;
  wire x34786, x34790, x34793, x34796, x34800, x34803, x34806, x34810;
  wire x34813, x34816, x34820, x34823, x34826, x34830, x34833, x34836;
  wire x34840, x34843, x34846, x34850, x34853, x34856, x34860, x34863;
  wire x34866, x34870, x34873, x34876, x34880, x34883, x34886, x34890;
  wire x34893, x34896, x34900, x34903, x34906, x34910, x34912, x34918;
  wire x34922, x34924, x34927, x34929, x34932, x34934, x34937, x34939;
  wire x34942, x34944, x34947, x34949, x34952, x34954, x34957, x34959;
  wire x34962, x34964, x34967, x34969, x34972, x34974, x34977, x34979;
  wire x34982, x34984, x34987, x34989, x34992, x34994, x34997, x34999;
  wire x35002, x35004, x35007, x35009, x35012, x35014, x35017, x35019;
  wire x35022, x35024, x35027, x35029, x35032, x35034, x35037, x35039;
  wire x35042, x35043, x35044, x35045, x35046, x35047, x35048, x35049;
  wire x35050, x35051, x35052, x35053, x35054, x35055, x35056, x35057;
  wire x35058, x35059, x35060, x35061, x35062, x35063, x35064, x35065;
  wire x35066, x35067, x35073, x35077, x35081, x35085, x35089, x35093;
  wire x35097, x35101, x35105, x35109, x35113, x35117, x35121, x35125;
  wire x35129, x35133, x35137, x35141, x35145, x35149, x35153, x35157;
  wire x35161, x35165, x35166, x35168, x35171, x35174, x35177, x35179;
  wire x35182, x35184, x35187, x35189, x35192, x35194, x35197, x35199;
  wire x35202, x35204, x35207, x35209, x35212, x35214, x35217, x35219;
  wire x35222, x35224, x35227, x35229, x35232, x35234, x35237, x35239;
  wire x35242, x35244, x35247, x35249, x35252, x35254, x35257, x35259;
  wire x35262, x35264, x35267, x35269, x35272, x35274, x35277, x35279;
  wire x35282, x35283, x35284, x35286, x35289, x35292, x35295, x35298;
  wire x35301, x35303, x35306, x35308, x35311, x35313, x35316, x35318;
  wire x35321, x35323, x35326, x35328, x35331, x35333, x35336, x35338;
  wire x35341, x35343, x35346, x35348, x35351, x35353, x35356, x35358;
  wire x35361, x35363, x35366, x35368, x35371, x35373, x35376, x35378;
  wire x35381, x35383, x35386, x35387, x35388, x35389, x35390, x35392;
  wire x35395, x35398, x35401, x35404, x35407, x35410, x35413, x35416;
  wire x35419, x35421, x35424, x35426, x35429, x35431, x35434, x35436;
  wire x35439, x35441, x35444, x35446, x35449, x35451, x35454, x35456;
  wire x35459, x35461, x35464, x35465, x35466, x35467, x35468, x35469;
  wire x35470, x35472, x35475, x35478, x35481, x35484, x35487, x35490;
  wire x35493, x35496, x35499, x35503, x35507, x35511, x35515, x35519;
  wire x35523, x35527, x35531, x35533, x35536, x35538, x35541, x35545;
  wire x35549, x35553, x35557, x35561, x35565, x35567, x35570, x35572;
  wire x35575, x35577, x35580, x35582, x35585, x35587, x35590, x35592;
  wire x35595, x35597, x35600, x35602, x35605, x35607, x35610, x35612;
  wire x35615, x35617, x35619, x35621, x35623, x35625, x35627, x35629;
  wire x35631, x35633, x35635, x35637, x35639, x35641, x35643, x35645;
  wire x35647, x35649, x35651, x35653, x35655, x35657, x35659, x35661;
  wire x35663, x35665, x35667, x35669, x35671, x35673, x35675, x35678;
  wire x35680, x35682, x35684, x35686, x35688, x35690, x35692, x35694;
  wire x35696, x35698, x35700, x35702, x35704, x35706, x35708, x35710;
  wire x35712, x35714, x35716, x35718, x35720, x35722, x35724, x35726;
  wire x35728, x35730, x35732, x35737, x35739, x35741, x35743, x35745;
  wire x35747, x35749, x35751, x35753, x35755, x35757, x35759, x35761;
  wire x35763, x35765, x35767, x35769, x35771, x35773, x35775, x35777;
  wire x35779, x35781, x35783, x35793, x35795, x35797, x35799, x35801;
  wire x35803, x35805, x35807, x35809, x35811, x35813, x35815, x35817;
  wire x35819, x35821, x35839, x35843, x35847, x35851, x35855, x35859;
  wire x35863, x35867, x35871, x35875, x35879, x35883, x35887, x35891;
  wire x35895, x35899, x35903, x35907, x35911, x35915, x35919, x35923;
  wire x35927, x35931, x35935, x35939, x35943, x35947, x35951, x35955;
  wire x35959, x35960, x35962, x35964, x35966, x35968, x35970, x35972;
  wire x35974, x35976, x35978, x35980, x35982, x35984, x35986, x35988;
  wire x35990, x35992, x36026, x36028, x36030, x36032, x36034, x36036;
  wire x36038, x36040, x36042, x36044, x36046, x36048, x36050, x36052;
  wire x36054, x36056, x36058, x36060, x36062, x36064, x36066, x36068;
  wire x36070, x36072, x36074, x36076, x36078, x36080, x36082, x36084;
  wire x36086, x36088, x38911, x38912, x38913, x38914, x38915, x38916;
  wire x38917, x38918, x38919, x38920, x38921, x38922, x38923, x38924;
  wire x38925, x38926, x38927, x38928, x38929, x38930, x38931, x38932;
  wire x38933, x38934, x38935, x38936, x38937, x38938, x38939, x38940;
  wire x38941, x38942, x39040, x39041, x39044, x39046, x39047, x39050;
  wire x39052, x39053, x39056, x39058, x39059, x39062, x39064, x39065;
  wire x39068, x39070, x39071, x39074, x39076, x39077, x39080, x39082;
  wire x39083, x39086, x39088, x39089, x39092, x39094, x39095, x39098;
  wire x39100, x39101, x39104, x39106, x39107, x39110, x39112, x39113;
  wire x39116, x39118, x39119, x39122, x39124, x39125, x39128, x39130;
  wire x39131, x39134, x39136, x39137, x39140, x39142, x39143, x39146;
  wire x39148, x39149, x39152, x39154, x39155, x39158, x39160, x39161;
  wire x39164, x39166, x39167, x39170, x39172, x39173, x39176, x39178;
  wire x39179, x39182, x39184, x39185, x39188, x39190, x39191, x39194;
  wire x39196, x39197, x39200, x39202, x39203, x39206, x39208, x39209;
  wire x39212, x39214, x39215, x39218, x39220, x39221, x39224, x39226;
  wire x39227, x39230, x39231, x39232, x39233, x39234, x39235, x39236;
  wire x39237, x39238, x39239, x39240, x39241, x39242, x39243, x39244;
  wire x39245, x39246, x39247, x39248, x39249, x39250, x39251, x39252;
  wire x39253, x39254, x39255, x39256, x39257, x39258, x39259, x39260;
  wire x39266, x39270, x39274, x39278, x39282, x39286, x39290, x39294;
  wire x39298, x39302, x39306, x39310, x39314, x39318, x39322, x39326;
  wire x39330, x39334, x39338, x39342, x39346, x39350, x39354, x39358;
  wire x39362, x39366, x39370, x39374, x39378, x39382, x39384, x39387;
  wire x39390, x39393, x39395, x39398, x39400, x39403, x39405, x39408;
  wire x39410, x39413, x39415, x39418, x39420, x39423, x39425, x39428;
  wire x39430, x39433, x39435, x39438, x39440, x39443, x39445, x39448;
  wire x39450, x39453, x39455, x39458, x39460, x39463, x39465, x39468;
  wire x39470, x39473, x39475, x39478, x39480, x39483, x39485, x39488;
  wire x39490, x39493, x39495, x39498, x39500, x39503, x39505, x39508;
  wire x39510, x39513, x39515, x39518, x39520, x39523, x39525, x39528;
  wire x39530, x39533, x39536, x39539, x39542, x39545, x39547, x39550;
  wire x39552, x39555, x39557, x39560, x39562, x39565, x39567, x39570;
  wire x39572, x39575, x39577, x39580, x39582, x39585, x39587, x39590;
  wire x39592, x39595, x39597, x39600, x39602, x39605, x39607, x39610;
  wire x39612, x39615, x39617, x39620, x39622, x39625, x39627, x39630;
  wire x39632, x39635, x39637, x39640, x39642, x39645, x39647, x39650;
  wire x39652, x39655, x39657, x39660, x39662, x39665, x39668, x39671;
  wire x39674, x39677, x39680, x39683, x39686, x39689, x39691, x39694;
  wire x39696, x39699, x39701, x39704, x39706, x39709, x39711, x39714;
  wire x39716, x39719, x39721, x39724, x39726, x39729, x39731, x39734;
  wire x39736, x39739, x39741, x39744, x39746, x39749, x39751, x39754;
  wire x39756, x39759, x39761, x39764, x39766, x39769, x39772, x39775;
  wire x39778, x39781, x39784, x39787, x39790, x39793, x39796, x39799;
  wire x39802, x39805, x39808, x39811, x39815, x39817, x39820, x39822;
  wire x39825, x39827, x39830, x39832, x39835, x39837, x39840, x39842;
  wire x39845, x39847, x39850, x39852, x39855, x39857, x39860, x39862;
  wire x39865, x39867, x39870, x39872, x39875, x39877, x39880, x39882;
  wire x39885, x39887, x39890, x39892, x39895, x39897, x39900, x39902;
  wire x39905, x39907, x39910, x39912, x39915, x39917, x39920, x39922;
  wire x39925, x39927, x39930, x39932, x39935, x39937, x39940, x39942;
  wire x39945, x39947, x39950, x39952, x39955, x39957, x39960, x39962;
  wire x39965, x39967, x39970, x39973, x39975, x39977, x39979, x39981;
  wire x39983, x39985, x39987, x39990, x39992, x39994, x39996, x39998;
  wire x40000, x40002, x40004, x40006, x40008, x40010, x40012, x40014;
  wire x40016, x40018, x40020, x40022, x40025, x40027, x40029, x40031;
  wire x40033, x40035, x40037, x40039, x40041, x40043, x40045, x40047;
  wire x40049, x40051, x40053, x40055, x40057, x40059, x40061, x40063;
  wire x40065, x40067, x40069, x40071, x40073, x40075, x40078, x40080;
  wire x40082, x40084, x40086, x40088, x40090, x40092, x40094, x40096;
  wire x40098, x40100, x40102, x40104, x40106, x40108, x40110, x40112;
  wire x40114, x40116, x40118, x40120, x40122, x40124, x40126, x40128;
  wire x40130, x40132, x40134, x40136, x40138, x40140, x40142, x40144;
  wire x40146, x40149, x40151, x40153, x40155, x40157, x40159, x40161;
  wire x40163, x40165, x40167, x40169, x40171, x40173, x40175, x40177;
  wire x40179, x40181, x40183, x40185, x40187, x40189, x40191, x40193;
  wire x40195, x40197, x40199, x40201, x40203, x40205, x40207, x40209;
  wire x40211, x40213, x40215, x40217, x40219, x40221, x40223, x40225;
  wire x40227, x40229, x40231, x40233, x40235, x40238, x40240, x40242;
  wire x40244, x40246, x40248, x40250, x40252, x40254, x40256, x40258;
  wire x40260, x40262, x40264, x40266, x40268, x40270, x40272, x40274;
  wire x40276, x40278, x40280, x40282, x40284, x40286, x40288, x40290;
  wire x40292, x40294, x40296, x40298, x40300, x40302, x40304, x40306;
  wire x40308, x40310, x40312, x40314, x40316, x40318, x40320, x40322;
  wire x40324, x40326, x40328, x40330, x40332, x40334, x40336, x40338;
  wire x40340, x40342, x40345, x40347, x40349, x40351, x40353, x40355;
  wire x40357, x40359, x40361, x40363, x40365, x40367, x40369, x40371;
  wire x40373, x40375, x40377, x40379, x40381, x40383, x40385, x40387;
  wire x40389, x40391, x40393, x40395, x40397, x40399, x40401, x40403;
  wire x40405, x40407, x40409, x40411, x40413, x40415, x40417, x40419;
  wire x40421, x40423, x40425, x40427, x40429, x40431, x40433, x40435;
  wire x40437, x40439, x40441, x40443, x40445, x40447, x40449, x40451;
  wire x40453, x40455, x40457, x40459, x40461, x40463, x40465, x40467;
  wire x40470, x40472, x40474, x40476, x40478, x40480, x40482, x40484;
  wire x40486, x40488, x40490, x40492, x40494, x40496, x40498, x40500;
  wire x40502, x40504, x40506, x40508, x40510, x40512, x40514, x40516;
  wire x40518, x40520, x40522, x40524, x40526, x40528, x40530, x40532;
  wire x40534, x40536, x40538, x40540, x40542, x40544, x40546, x40548;
  wire x40550, x40552, x40554, x40556, x40558, x40560, x40562, x40564;
  wire x40566, x40568, x40570, x40572, x40574, x40576, x40578, x40580;
  wire x40582, x40584, x40586, x40588, x40590, x40592, x40594, x40596;
  wire x40598, x40600, x40602, x40604, x40606, x40608, x40610, x40613;
  wire x40615, x40617, x40619, x40621, x40623, x40625, x40627, x40629;
  wire x40631, x40633, x40635, x40637, x40639, x40641, x40643, x40645;
  wire x40647, x40649, x40651, x40653, x40655, x40657, x40659, x40661;
  wire x40663, x40665, x40667, x40669, x40671, x40673, x40675, x40677;
  wire x40679, x40681, x40683, x40685, x40687, x40689, x40691, x40693;
  wire x40695, x40697, x40699, x40701, x40703, x40705, x40707, x40709;
  wire x40711, x40713, x40715, x40717, x40719, x40721, x40723, x40725;
  wire x40727, x40729, x40731, x40733, x40735, x40737, x40739, x40741;
  wire x40743, x40745, x40747, x40749, x40751, x40753, x40755, x40757;
  wire x40759, x40761, x40763, x40765, x40767, x40769, x40771, x40774;
  wire x40776, x40778, x40780, x40782, x40784, x40786, x40788, x40790;
  wire x40792, x40794, x40796, x40798, x40800, x40802, x40804, x40806;
  wire x40808, x40810, x40812, x40814, x40816, x40818, x40820, x40822;
  wire x40824, x40826, x40828, x40830, x40832, x40834, x40836, x40838;
  wire x40840, x40842, x40844, x40846, x40848, x40850, x40852, x40854;
  wire x40856, x40858, x40860, x40862, x40864, x40866, x40868, x40870;
  wire x40872, x40874, x40876, x40878, x40880, x40882, x40884, x40886;
  wire x40888, x40890, x40892, x40894, x40896, x40898, x40900, x40902;
  wire x40904, x40906, x40908, x40910, x40912, x40914, x40916, x40918;
  wire x40920, x40922, x40924, x40926, x40928, x40930, x40932, x40934;
  wire x40936, x40938, x40940, x40942, x40944, x40946, x40948, x40950;
  wire x40953, x40955, x40957, x40959, x40961, x40963, x40965, x40967;
  wire x40969, x40971, x40973, x40975, x40977, x40979, x40981, x40983;
  wire x40985, x40987, x40989, x40991, x40993, x40995, x40997, x40999;
  wire x41001, x41003, x41005, x41007, x41009, x41011, x41013, x41015;
  wire x41022, x41030, x41038, x41049, x41057, x41065, x41073, x41077;
  wire x41082, x41090, x41094, x41102, x41110, x41114, x41119, x41123;
  wire x41128, x41136, x41140, x41145, x41149, x41154, x41162, x41166;
  wire x41171, x41175, x41183, x41191, x41195, x41200, x41204, x41209;
  wire x41213, x41218, x41226, x41230, x41235, x41239, x41244, x41248;
  wire x41253, x41261, x41265, x41270, x41274, x41279, x41283, x41291;
  wire x41299, x41303, x41308, x41312, x41317, x41321, x41326, x41334;
  wire x41342, x41346, x41351, x41355, x41360, x41364, x41369, x41373;
  wire x41378, x41386, x41390, x41395, x41399, x41404, x41408, x41413;
  wire x41417, x41425, x41433, x41437, x41442, x41446, x41451, x41455;
  wire x41460, x41464, x41469, x41473, x41478, x41486, x41490, x41495;
  wire x41499, x41504, x41508, x41513, x41517, x41522, x41526, x41531;
  wire x41539, x41543, x41548, x41552, x41557, x41561, x41566, x41570;
  wire x41575, x41579, x41587, x41595, x41599, x41604, x41608, x41613;
  wire x41617, x41622, x41626, x41631, x41635, x41640, x41644, x41649;
  wire x41657, x41661, x41666, x41670, x41675, x41679, x41684, x41688;
  wire x41693, x41697, x41702, x41706, x41711, x41719, x41723, x41728;
  wire x41732, x41737, x41741, x41746, x41750, x41755, x41759, x41764;
  wire x41768, x41776, x41784, x41788, x41793, x41797, x41802, x41806;
  wire x41811, x41815, x41820, x41824, x41829, x41833, x41838, x41846;
  wire x41854, x41858, x41863, x41867, x41872, x41876, x41881, x41885;
  wire x41890, x41894, x41899, x41903, x41908, x41912, x41917, x41925;
  wire x41929, x41934, x41938, x41943, x41947, x41952, x41956, x41961;
  wire x41965, x41970, x41974, x41979, x41983, x41991, x41999, x42003;
  wire x42008, x42012, x42017, x42021, x42026, x42030, x42035, x42039;
  wire x42044, x42048, x42053, x42057, x42062, x42066, x42071, x42079;
  wire x42083, x42088, x42092, x42097, x42101, x42106, x42110, x42115;
  wire x42119, x42124, x42128, x42133, x42137, x42142, x42146, x42151;
  wire x42159, x42163, x42168, x42172, x42177, x42181, x42186, x42190;
  wire x42195, x42199, x42204, x42208, x42213, x42217, x42222, x42226;
  wire x42234, x42238, x42243, x42247, x42252, x42256, x42261, x42265;
  wire x42270, x42274, x42279, x42283, x42288, x42292, x42297, x42301;
  wire x42306, x42310, x42315, x42319, x42324, x42328, x42333, x42337;
  wire x42342, x42346, x42351, x42355, x42360, x42364, x42369, x42373;
  wire x42378, x42382, x42387, x42391, x42396, x42400, x42405, x42409;
  wire x42414, x42418, x42422, x42426, x42430, x42434, x42438, x42442;
  wire x42446, x42450, x42454, x42458, x42462, x42466, x42470, x42474;
  wire x42478, x42482, x42486, x42490, x42494, x42495, x42496, x42498;
  wire x42502, x42503, x42510, x42511, x42518, x42519, x42522, x42531;
  wire x42532, x42535, x42537, x42544, x42548, x42551, x42552, x42555;
  wire x42557, x42564, x42568, x42571, x42572, x42575, x42577, x42584;
  wire x42588, x42591, x42592, x42595, x42597, x42601, x42605, x42609;
  wire x42612, x42613, x42616, x42618, x42622, x42626, x42630, x42633;
  wire x42634, x42637, x42639, x42644, x42650, x42654, x42657, x42658;
  wire x42661, x42663, x42668, x42669, x42675, x42679, x42685, x42686;
  wire x42689, x42691, x42696, x42697, x42703, x42707, x42713, x42714;
  wire x42717, x42719, x42724, x42725, x42728, x42732, x42737, x42741;
  wire x42747, x42748, x42751, x42753, x42758, x42759, x42762, x42764;
  wire x42767, x42772, x42776, x42781, x42787, x42788, x42791, x42793;
  wire x42798, x42799, x42802, x42804, x42807, x42812, x42816, x42821;
  wire x42827, x42828, x42831, x42833, x42838, x42839, x42842, x42844;
  wire x42847, x42852, x42856, x42861, x42867, x42868, x42871, x42873;
  wire x42878, x42879, x42882, x42884, x42887, x42889, x42893, x42897;
  wire x42902, x42906, x42909, x42910, x42913, x42915, x42920, x42921;
  wire x42924, x42926, x42929, x42931, x42935, x42939, x42944, x42948;
  wire x42951, x42952, x42955, x42957, x42962, x42963, x42966, x42968;
  wire x42971, x42974, x42980, x42984, x42989, x42993, x42996, x42997;
  wire x43000, x43002, x43007, x43008, x43011, x43013, x43016, x43019;
  wire x43020, x43026, x43030, x43035, x43039, x43045, x43046, x43049;
  wire x43051, x43054, x43057, x43058, x43061, x43063, x43066, x43069;
  wire x43070, x43076, x43080, x43085, x43089, x43095, x43096, x43099;
  wire x43101, x43104, x43107, x43108, x43111, x43113, x43116, x43119;
  wire x43120, x43123, x43127, x43132, x43136, x43141, x43145, x43151;
  wire x43152, x43155, x43157, x43160, x43163, x43164, x43167, x43169;
  wire x43172, x43175, x43176, x43179, x43181, x43184, x43189, x43193;
  wire x43198, x43202, x43207, x43211, x43214, x43215, x43218, x43220;
  wire x43223, x43226, x43227, x43230, x43232, x43235, x43238, x43239;
  wire x43242, x43244, x43247, x43252, x43256, x43261, x43265, x43270;
  wire x43274, x43277, x43278, x43281, x43283, x43286, x43289, x43290;
  wire x43293, x43295, x43298, x43301, x43302, x43305, x43307, x43310;
  wire x43315, x43319, x43323, x43328, x43332, x43337, x43341, x43344;
  wire x43345, x43348, x43350, x43353, x43356, x43357, x43360, x43362;
  wire x43365, x43368, x43369, x43372, x43374, x43377, x43379, x43383;
  wire x43387, x43391, x43396, x43400, x43405, x43409, x43412, x43413;
  wire x43416, x43418, x43421, x43423, x43424, x43427, x43429, x43432;
  wire x43434, x43435, x43438, x43440, x43443, x43444, x43448, x43452;
  wire x43456, x43460, x43464, x43468, x43472, x43476, x43480, x43484;
  wire x43488, x43492, x43496, x43497, x43501, x43502, x43503, x43507;
  wire x43508, x43509, x43513, x43517, x43518, x43519, x43523, x43527;
  wire x43528, x43529, x43533, x43537, x43538, x43539, x43543, x43547;
  wire x43549, x43552, x43556, x43560, x43562, x43565, x43569, x43573;
  wire x43577, x43579, x43582, x43586, x43590, x43594, x43596, x43597;
  wire x43600, x43604, x43608, x43612, x43614, x43615, x43618, x43620;
  wire x43623, x43627, x43631, x43633, x43634, x43637, x43639, x43642;
  wire x43646, x43650, x43654, x43657, x43658, x43661, x43663, x43666;
  wire x43670, x43674, x43678, x43684, x43685, x43688, x43690, x43693;
  wire x43697, x43701, x43705, x43711, x43712, x43715, x43717, x43720;
  wire x43724, x43728, x43732, x43738, x43739, x43742, x43746, x43748;
  wire x43750, x43753, x43757, x43761, x43765, x43771, x43772, x43775;
  wire x43779, x43781, x43783, x43786, x43790, x43794, x43799, x43803;
  wire x43809, x43810, x43813, x43817, x43819, x43821, x43824, x43828;
  wire x43832, x43837, x43841, x43847, x43848, x43851, x43853, x43856;
  wire x43858, x43860, x43863, x43867, x43871, x43876, x43880, x43886;
  wire x43887, x43890, x43892, x43895, x43897, x43899, x43902, x43904;
  wire x43907, x43911, x43916, x43920, x43926, x43927, x43930, x43932;
  wire x43935, x43937, x43939, x43942, x43944, x43947, x43951, x43956;
  wire x43960, x43966, x43967, x43970, x43972, x43975, x43978, x43981;
  wire x43983, x43986, x43989, x43992, x43996, x44001, x44005, x44010;
  wire x44014, x44017, x44018, x44021, x44023, x44026, x44028, x44031;
  wire x44033, x44036, x44038, x44041, x44045, x44049, x44053, x44057;
  wire x44061, x44071, x44075, x44082, x44089, x44093, x44101, x44105;
  wire x44113, x44117, x44125, x44129, x44137, x44141, x44146, x44150;
  wire x44154, x44159, x44163, x44167, x44172, x44176, x44180, x44185;
  wire x44189, x44193, x44198, x44202, x44206, x44210, x44215, x44219;
  wire x44224, x44228, x44232, x44237, x44241, x44246, x44250, x44254;
  wire x44259, x44263, x44268, x44272, x44276, x44281, x44285, x44290;
  wire x44294, x44298, x44303, x44307, x44309, x44313, x44317, x44321;
  wire x44326, x44330, x44333, x44336, x44340, x44345, x44349, x44354;
  wire x44358, x44361, x44364, x44368, x44373, x44377, x44382, x44386;
  wire x44389, x44392, x44396, x44401, x44405, x44408, x44411, x44415;
  wire x44418, x44421, x44425, x44430, x44434, x44437, x44440, x44442;
  wire x44445, x44448, x44451, x44455, x44460, x44464, x44467, x44470;
  wire x44472, x44475, x44478, x44481, x44485, x44490, x44494, x44497;
  wire x44500, x44502, x44505, x44508, x44511, x44515, x44520, x44524;
  wire x44527, x44530, x44532, x44535, x44538, x44541, x44545, x44550;
  wire x44554, x44557, x44560, x44562, x44565, x44568, x44571, x44575;
  wire x44580, x44584, x44587, x44588, x44591, x44593, x44596, x44598;
  wire x44599, x44602, x44606, x44610, x44614, x44627, x44632, x44635;
  wire x44640, x44643, x44648, x44651, x44656, x44659, x44664, x44667;
  wire x44671, x44675, x44678, x44681, x44685, x44689, x44692, x44695;
  wire x44699, x44703, x44706, x44709, x44713, x44717, x44720, x44723;
  wire x44727, x44731, x44736, x44738, x44741, x44746, x44750, x44753;
  wire x44756, x44758, x44761, x44766, x44770, x44773, x44776, x44778;
  wire x44781, x44786, x44790, x44793, x44796, x44798, x44801, x44806;
  wire x44810, x44813, x44816, x44818, x44821, x44826, x44830, x44833;
  wire x44836, x44838, x44841, x44846, x44850, x44853, x44854, x44857;
  wire x44859, x44862, x44867, x44871, x44874, x44875, x44878, x44880;
  wire x44883, x44888, x44892, x44895, x44896, x44899, x44901, x44904;
  wire x44909, x44913, x44916, x44917, x44920, x44922, x44925, x44930;
  wire x44934, x44937, x44938, x44941, x44943, x44946, x44951, x44955;
  wire x44958, x44959, x44962, x44964, x44967, x44972, x44976, x44979;
  wire x44980, x44983, x44985, x44988, x44993, x44997, x45000, x45001;
  wire x45004, x45006, x45009, x45014, x45018, x45021, x45022, x45025;
  wire x45027, x45030, x45034, x45038, x45045, x45049, x45053, x45057;
  wire x45062, x45066, x45071, x45075, x45080, x45084, x45089, x45093;
  wire x45098, x45099, x45101, x45104, x45108, x45113, x45114, x45116;
  wire x45119, x45123, x45128, x45129, x45131, x45134, x45138, x45143;
  wire x45144, x45146, x45149, x45153, x45158, x45159, x45161, x45164;
  wire x45168, x45173, x45174, x45176, x45177, x45180, x45184, x45189;
  wire x45190, x45192, x45193, x45196, x45200, x45205, x45206, x45208;
  wire x45209, x45212, x45216, x45221, x45222, x45224, x45225, x45228;
  wire x45232, x45237, x45238, x45240, x45241, x45244, x45248, x45253;
  wire x45254, x45256, x45257, x45260, x45264, x45269, x45270, x45272;
  wire x45273, x45276, x45280, x45285, x45286, x45288, x45289, x45292;
  wire x45296, x45301, x45302, x45304, x45305, x45308, x45312, x45317;
  wire x45318, x45320, x45321, x45324, x45328, x45333, x45334, x45336;
  wire x45337, x45340, x45344, x45349, x45350, x45352, x45353, x45356;
  wire x45360, x45365, x45366, x45368, x45369, x45372, x45376, x45381;
  wire x45382, x45384, x45385, x45388, x45392, x45396, x45406, x45410;
  wire x45411, x45415, x45416, x45420, x45421, x45425, x45426, x45430;
  wire x45432, x45435, x45439, x45442, x45445, x45449, x45452, x45455;
  wire x45459, x45462, x45465, x45469, x45472, x45475, x45479, x45482;
  wire x45485, x45489, x45492, x45495, x45499, x45502, x45505, x45509;
  wire x45512, x45515, x45519, x45522, x45525, x45529, x45532, x45535;
  wire x45539, x45542, x45545, x45549, x45552, x45555, x45559, x45562;
  wire x45565, x45569, x45572, x45575, x45579, x45582, x45585, x45589;
  wire x45592, x45595, x45599, x45602, x45605, x45609, x45612, x45615;
  wire x45619, x45623, x45631, x45635, x45639, x45643, x45648, x45652;
  wire x45657, x45661, x45666, x45670, x45675, x45679, x45684, x45688;
  wire x45693, x45697, x45700, x45703, x45707, x45710, x45713, x45717;
  wire x45720, x45723, x45727, x45730, x45733, x45737, x45740, x45743;
  wire x45747, x45750, x45753, x45757, x45760, x45763, x45767, x45770;
  wire x45773, x45777, x45780, x45783, x45787, x45790, x45793, x45797;
  wire x45800, x45803, x45807, x45810, x45813, x45817, x45820, x45823;
  wire x45827, x45830, x45833, x45837, x45840, x45843, x45847, x45850;
  wire x45853, x45857, x45860, x45863, x45867, x45870, x45873, x45877;
  wire x45879, x45885, x45889, x45891, x45894, x45896, x45899, x45901;
  wire x45904, x45906, x45909, x45911, x45914, x45916, x45919, x45921;
  wire x45924, x45926, x45929, x45931, x45934, x45936, x45939, x45941;
  wire x45944, x45946, x45949, x45951, x45954, x45956, x45959, x45961;
  wire x45964, x45966, x45969, x45971, x45974, x45976, x45979, x45981;
  wire x45984, x45986, x45989, x45991, x45994, x45996, x45999, x46001;
  wire x46004, x46006, x46009, x46010, x46011, x46012, x46013, x46014;
  wire x46015, x46016, x46017, x46018, x46019, x46020, x46021, x46022;
  wire x46023, x46024, x46025, x46026, x46027, x46028, x46029, x46030;
  wire x46031, x46032, x46033, x46034, x46040, x46044, x46048, x46052;
  wire x46056, x46060, x46064, x46068, x46072, x46076, x46080, x46084;
  wire x46088, x46092, x46096, x46100, x46104, x46108, x46112, x46116;
  wire x46120, x46124, x46128, x46132, x46133, x46135, x46138, x46141;
  wire x46144, x46146, x46149, x46151, x46154, x46156, x46159, x46161;
  wire x46164, x46166, x46169, x46171, x46174, x46176, x46179, x46181;
  wire x46184, x46186, x46189, x46191, x46194, x46196, x46199, x46201;
  wire x46204, x46206, x46209, x46211, x46214, x46216, x46219, x46221;
  wire x46224, x46226, x46229, x46231, x46234, x46236, x46239, x46241;
  wire x46244, x46246, x46249, x46250, x46251, x46253, x46256, x46259;
  wire x46262, x46265, x46268, x46270, x46273, x46275, x46278, x46280;
  wire x46283, x46285, x46288, x46290, x46293, x46295, x46298, x46300;
  wire x46303, x46305, x46308, x46310, x46313, x46315, x46318, x46320;
  wire x46323, x46325, x46328, x46330, x46333, x46335, x46338, x46340;
  wire x46343, x46345, x46348, x46350, x46353, x46354, x46355, x46356;
  wire x46357, x46359, x46362, x46365, x46368, x46371, x46374, x46377;
  wire x46380, x46383, x46386, x46388, x46391, x46393, x46396, x46398;
  wire x46401, x46403, x46406, x46408, x46411, x46413, x46416, x46418;
  wire x46421, x46423, x46426, x46428, x46431, x46432, x46433, x46434;
  wire x46435, x46436, x46437, x46439, x46442, x46445, x46448, x46451;
  wire x46454, x46457, x46460, x46463, x46466, x46470, x46474, x46478;
  wire x46482, x46486, x46490, x46494, x46498, x46500, x46503, x46505;
  wire x46508, x46512, x46516, x46520, x46524, x46528, x46532, x46534;
  wire x46537, x46539, x46542, x46544, x46547, x46549, x46552, x46554;
  wire x46557, x46559, x46562, x46564, x46567, x46569, x46572, x46574;
  wire x46577, x46579, x46582, x46584, x46586, x46588, x46590, x46592;
  wire x46594, x46596, x46598, x46600, x46602, x46604, x46606, x46608;
  wire x46610, x46612, x46614, x46616, x46618, x46620, x46622, x46624;
  wire x46626, x46628, x46630, x46632, x46634, x46636, x46638, x46640;
  wire x46642, x46645, x46647, x46649, x46651, x46653, x46655, x46657;
  wire x46659, x46661, x46663, x46665, x46667, x46669, x46671, x46673;
  wire x46675, x46677, x46679, x46681, x46683, x46685, x46687, x46689;
  wire x46691, x46693, x46695, x46697, x46699, x46704, x46706, x46708;
  wire x46710, x46712, x46714, x46716, x46718, x46720, x46722, x46724;
  wire x46726, x46728, x46730, x46732, x46734, x46736, x46738, x46740;
  wire x46742, x46744, x46746, x46748, x46750, x46760, x46762, x46764;
  wire x46766, x46768, x46770, x46772, x46774, x46776, x46778, x46780;
  wire x46782, x46784, x46786, x46788, x46806, x46810, x46814, x46818;
  wire x46822, x46826, x46830, x46834, x46838, x46842, x46846, x46850;
  wire x46854, x46858, x46862, x46866, x46870, x46874, x46878, x46882;
  wire x46886, x46890, x46894, x46898, x46902, x46906, x46910, x46914;
  wire x46918, x46922, x46926, x46927, x46929, x46931, x46933, x46935;
  wire x46937, x46939, x46941, x46943, x46945, x46947, x46949, x46951;
  wire x46953, x46955, x46957, x46959, x46993, x46995, x46997, x46999;
  wire x47001, x47003, x47005, x47007, x47009, x47011, x47013, x47015;
  wire x47017, x47019, x47021, x47023, x47025, x47027, x47029, x47031;
  wire x47033, x47035, x47037, x47039, x47041, x47043, x47045, x47047;
  wire x47049, x47051, x47053, x47055, x49878, x49879, x49880, x49881;
  wire x49882, x49883, x49884, x49885, x49886, x49887, x49888, x49889;
  wire x49890, x49891, x49892, x49893, x49894, x49895, x49896, x49897;
  wire x49898, x49899, x49900, x49901, x49902, x49903, x49904, x49905;
  wire x49906, x49907, x49908, x49909, x50007, x50008, x50011, x50013;
  wire x50014, x50017, x50019, x50020, x50023, x50025, x50026, x50029;
  wire x50031, x50032, x50035, x50037, x50038, x50041, x50043, x50044;
  wire x50047, x50049, x50050, x50053, x50055, x50056, x50059, x50061;
  wire x50062, x50065, x50067, x50068, x50071, x50073, x50074, x50077;
  wire x50079, x50080, x50083, x50085, x50086, x50089, x50091, x50092;
  wire x50095, x50097, x50098, x50101, x50103, x50104, x50107, x50109;
  wire x50110, x50113, x50115, x50116, x50119, x50121, x50122, x50125;
  wire x50127, x50128, x50131, x50133, x50134, x50137, x50139, x50140;
  wire x50143, x50145, x50146, x50149, x50151, x50152, x50155, x50157;
  wire x50158, x50161, x50163, x50164, x50167, x50169, x50170, x50173;
  wire x50175, x50176, x50179, x50181, x50182, x50185, x50187, x50188;
  wire x50191, x50193, x50194, x50197, x50198, x50199, x50200, x50201;
  wire x50202, x50203, x50204, x50205, x50206, x50207, x50208, x50209;
  wire x50210, x50211, x50212, x50213, x50214, x50215, x50216, x50217;
  wire x50218, x50219, x50220, x50221, x50222, x50223, x50224, x50225;
  wire x50226, x50227, x50233, x50237, x50241, x50245, x50249, x50253;
  wire x50257, x50261, x50265, x50269, x50273, x50277, x50281, x50285;
  wire x50289, x50293, x50297, x50301, x50305, x50309, x50313, x50317;
  wire x50321, x50325, x50329, x50333, x50337, x50341, x50345, x50349;
  wire x50351, x50354, x50357, x50360, x50362, x50365, x50367, x50370;
  wire x50372, x50375, x50377, x50380, x50382, x50385, x50387, x50390;
  wire x50392, x50395, x50397, x50400, x50402, x50405, x50407, x50410;
  wire x50412, x50415, x50417, x50420, x50422, x50425, x50427, x50430;
  wire x50432, x50435, x50437, x50440, x50442, x50445, x50447, x50450;
  wire x50452, x50455, x50457, x50460, x50462, x50465, x50467, x50470;
  wire x50472, x50475, x50477, x50480, x50482, x50485, x50487, x50490;
  wire x50492, x50495, x50497, x50500, x50503, x50506, x50509, x50512;
  wire x50514, x50517, x50519, x50522, x50524, x50527, x50529, x50532;
  wire x50534, x50537, x50539, x50542, x50544, x50547, x50549, x50552;
  wire x50554, x50557, x50559, x50562, x50564, x50567, x50569, x50572;
  wire x50574, x50577, x50579, x50582, x50584, x50587, x50589, x50592;
  wire x50594, x50597, x50599, x50602, x50604, x50607, x50609, x50612;
  wire x50614, x50617, x50619, x50622, x50624, x50627, x50629, x50632;
  wire x50635, x50638, x50641, x50644, x50647, x50650, x50653, x50656;
  wire x50658, x50661, x50663, x50666, x50668, x50671, x50673, x50676;
  wire x50678, x50681, x50683, x50686, x50688, x50691, x50693, x50696;
  wire x50698, x50701, x50703, x50706, x50708, x50711, x50713, x50716;
  wire x50718, x50721, x50723, x50726, x50728, x50731, x50733, x50736;
  wire x50739, x50742, x50745, x50748, x50751, x50754, x50757, x50760;
  wire x50763, x50766, x50769, x50772, x50775, x50778, x50782, x50784;
  wire x50787, x50789, x50792, x50794, x50797, x50799, x50802, x50804;
  wire x50807, x50809, x50812, x50814, x50817, x50819, x50822, x50824;
  wire x50827, x50829, x50832, x50834, x50837, x50839, x50842, x50844;
  wire x50847, x50849, x50852, x50854, x50857, x50859, x50862, x50864;
  wire x50867, x50869, x50872, x50874, x50877, x50879, x50882, x50884;
  wire x50887, x50889, x50892, x50894, x50897, x50899, x50902, x50904;
  wire x50907, x50909, x50912, x50914, x50917, x50919, x50922, x50924;
  wire x50927, x50929, x50932, x50934, x50937, x50940, x50942, x50944;
  wire x50946, x50948, x50950, x50952, x50954, x50957, x50959, x50961;
  wire x50963, x50965, x50967, x50969, x50971, x50973, x50975, x50977;
  wire x50979, x50981, x50983, x50985, x50987, x50989, x50992, x50994;
  wire x50996, x50998, x51000, x51002, x51004, x51006, x51008, x51010;
  wire x51012, x51014, x51016, x51018, x51020, x51022, x51024, x51026;
  wire x51028, x51030, x51032, x51034, x51036, x51038, x51040, x51042;
  wire x51045, x51047, x51049, x51051, x51053, x51055, x51057, x51059;
  wire x51061, x51063, x51065, x51067, x51069, x51071, x51073, x51075;
  wire x51077, x51079, x51081, x51083, x51085, x51087, x51089, x51091;
  wire x51093, x51095, x51097, x51099, x51101, x51103, x51105, x51107;
  wire x51109, x51111, x51113, x51116, x51118, x51120, x51122, x51124;
  wire x51126, x51128, x51130, x51132, x51134, x51136, x51138, x51140;
  wire x51142, x51144, x51146, x51148, x51150, x51152, x51154, x51156;
  wire x51158, x51160, x51162, x51164, x51166, x51168, x51170, x51172;
  wire x51174, x51176, x51178, x51180, x51182, x51184, x51186, x51188;
  wire x51190, x51192, x51194, x51196, x51198, x51200, x51202, x51205;
  wire x51207, x51209, x51211, x51213, x51215, x51217, x51219, x51221;
  wire x51223, x51225, x51227, x51229, x51231, x51233, x51235, x51237;
  wire x51239, x51241, x51243, x51245, x51247, x51249, x51251, x51253;
  wire x51255, x51257, x51259, x51261, x51263, x51265, x51267, x51269;
  wire x51271, x51273, x51275, x51277, x51279, x51281, x51283, x51285;
  wire x51287, x51289, x51291, x51293, x51295, x51297, x51299, x51301;
  wire x51303, x51305, x51307, x51309, x51312, x51314, x51316, x51318;
  wire x51320, x51322, x51324, x51326, x51328, x51330, x51332, x51334;
  wire x51336, x51338, x51340, x51342, x51344, x51346, x51348, x51350;
  wire x51352, x51354, x51356, x51358, x51360, x51362, x51364, x51366;
  wire x51368, x51370, x51372, x51374, x51376, x51378, x51380, x51382;
  wire x51384, x51386, x51388, x51390, x51392, x51394, x51396, x51398;
  wire x51400, x51402, x51404, x51406, x51408, x51410, x51412, x51414;
  wire x51416, x51418, x51420, x51422, x51424, x51426, x51428, x51430;
  wire x51432, x51434, x51437, x51439, x51441, x51443, x51445, x51447;
  wire x51449, x51451, x51453, x51455, x51457, x51459, x51461, x51463;
  wire x51465, x51467, x51469, x51471, x51473, x51475, x51477, x51479;
  wire x51481, x51483, x51485, x51487, x51489, x51491, x51493, x51495;
  wire x51497, x51499, x51501, x51503, x51505, x51507, x51509, x51511;
  wire x51513, x51515, x51517, x51519, x51521, x51523, x51525, x51527;
  wire x51529, x51531, x51533, x51535, x51537, x51539, x51541, x51543;
  wire x51545, x51547, x51549, x51551, x51553, x51555, x51557, x51559;
  wire x51561, x51563, x51565, x51567, x51569, x51571, x51573, x51575;
  wire x51577, x51580, x51582, x51584, x51586, x51588, x51590, x51592;
  wire x51594, x51596, x51598, x51600, x51602, x51604, x51606, x51608;
  wire x51610, x51612, x51614, x51616, x51618, x51620, x51622, x51624;
  wire x51626, x51628, x51630, x51632, x51634, x51636, x51638, x51640;
  wire x51642, x51644, x51646, x51648, x51650, x51652, x51654, x51656;
  wire x51658, x51660, x51662, x51664, x51666, x51668, x51670, x51672;
  wire x51674, x51676, x51678, x51680, x51682, x51684, x51686, x51688;
  wire x51690, x51692, x51694, x51696, x51698, x51700, x51702, x51704;
  wire x51706, x51708, x51710, x51712, x51714, x51716, x51718, x51720;
  wire x51722, x51724, x51726, x51728, x51730, x51732, x51734, x51736;
  wire x51738, x51741, x51743, x51745, x51747, x51749, x51751, x51753;
  wire x51755, x51757, x51759, x51761, x51763, x51765, x51767, x51769;
  wire x51771, x51773, x51775, x51777, x51779, x51781, x51783, x51785;
  wire x51787, x51789, x51791, x51793, x51795, x51797, x51799, x51801;
  wire x51803, x51805, x51807, x51809, x51811, x51813, x51815, x51817;
  wire x51819, x51821, x51823, x51825, x51827, x51829, x51831, x51833;
  wire x51835, x51837, x51839, x51841, x51843, x51845, x51847, x51849;
  wire x51851, x51853, x51855, x51857, x51859, x51861, x51863, x51865;
  wire x51867, x51869, x51871, x51873, x51875, x51877, x51879, x51881;
  wire x51883, x51885, x51887, x51889, x51891, x51893, x51895, x51897;
  wire x51899, x51901, x51903, x51905, x51907, x51909, x51911, x51913;
  wire x51915, x51917, x51920, x51922, x51924, x51926, x51928, x51930;
  wire x51932, x51934, x51936, x51938, x51940, x51942, x51944, x51946;
  wire x51948, x51950, x51952, x51954, x51956, x51958, x51960, x51962;
  wire x51964, x51966, x51968, x51970, x51972, x51974, x51976, x51978;
  wire x51980, x51982, x51989, x51997, x52005, x52016, x52024, x52032;
  wire x52040, x52044, x52049, x52057, x52061, x52069, x52077, x52081;
  wire x52086, x52090, x52095, x52103, x52107, x52112, x52116, x52121;
  wire x52129, x52133, x52138, x52142, x52150, x52158, x52162, x52167;
  wire x52171, x52176, x52180, x52185, x52193, x52197, x52202, x52206;
  wire x52211, x52215, x52220, x52228, x52232, x52237, x52241, x52246;
  wire x52250, x52258, x52266, x52270, x52275, x52279, x52284, x52288;
  wire x52293, x52301, x52309, x52313, x52318, x52322, x52327, x52331;
  wire x52336, x52340, x52345, x52353, x52357, x52362, x52366, x52371;
  wire x52375, x52380, x52384, x52392, x52400, x52404, x52409, x52413;
  wire x52418, x52422, x52427, x52431, x52436, x52440, x52445, x52453;
  wire x52457, x52462, x52466, x52471, x52475, x52480, x52484, x52489;
  wire x52493, x52498, x52506, x52510, x52515, x52519, x52524, x52528;
  wire x52533, x52537, x52542, x52546, x52554, x52562, x52566, x52571;
  wire x52575, x52580, x52584, x52589, x52593, x52598, x52602, x52607;
  wire x52611, x52616, x52624, x52628, x52633, x52637, x52642, x52646;
  wire x52651, x52655, x52660, x52664, x52669, x52673, x52678, x52686;
  wire x52690, x52695, x52699, x52704, x52708, x52713, x52717, x52722;
  wire x52726, x52731, x52735, x52743, x52751, x52755, x52760, x52764;
  wire x52769, x52773, x52778, x52782, x52787, x52791, x52796, x52800;
  wire x52805, x52813, x52821, x52825, x52830, x52834, x52839, x52843;
  wire x52848, x52852, x52857, x52861, x52866, x52870, x52875, x52879;
  wire x52884, x52892, x52896, x52901, x52905, x52910, x52914, x52919;
  wire x52923, x52928, x52932, x52937, x52941, x52946, x52950, x52958;
  wire x52966, x52970, x52975, x52979, x52984, x52988, x52993, x52997;
  wire x53002, x53006, x53011, x53015, x53020, x53024, x53029, x53033;
  wire x53038, x53046, x53050, x53055, x53059, x53064, x53068, x53073;
  wire x53077, x53082, x53086, x53091, x53095, x53100, x53104, x53109;
  wire x53113, x53118, x53126, x53130, x53135, x53139, x53144, x53148;
  wire x53153, x53157, x53162, x53166, x53171, x53175, x53180, x53184;
  wire x53189, x53193, x53201, x53205, x53210, x53214, x53219, x53223;
  wire x53228, x53232, x53237, x53241, x53246, x53250, x53255, x53259;
  wire x53264, x53268, x53273, x53277, x53282, x53286, x53291, x53295;
  wire x53300, x53304, x53309, x53313, x53318, x53322, x53327, x53331;
  wire x53336, x53340, x53345, x53349, x53354, x53358, x53363, x53367;
  wire x53372, x53376, x53381, x53385, x53389, x53393, x53397, x53401;
  wire x53405, x53409, x53413, x53417, x53421, x53425, x53429, x53433;
  wire x53437, x53441, x53445, x53449, x53453, x53457, x53461, x53462;
  wire x53463, x53465, x53469, x53470, x53477, x53478, x53485, x53486;
  wire x53489, x53498, x53499, x53502, x53504, x53511, x53515, x53518;
  wire x53519, x53522, x53524, x53531, x53535, x53538, x53539, x53542;
  wire x53544, x53551, x53555, x53558, x53559, x53562, x53564, x53568;
  wire x53572, x53576, x53579, x53580, x53583, x53585, x53589, x53593;
  wire x53597, x53600, x53601, x53604, x53606, x53611, x53617, x53621;
  wire x53624, x53625, x53628, x53630, x53635, x53636, x53642, x53646;
  wire x53652, x53653, x53656, x53658, x53663, x53664, x53670, x53674;
  wire x53680, x53681, x53684, x53686, x53691, x53692, x53695, x53699;
  wire x53704, x53708, x53714, x53715, x53718, x53720, x53725, x53726;
  wire x53729, x53731, x53734, x53739, x53743, x53748, x53754, x53755;
  wire x53758, x53760, x53765, x53766, x53769, x53771, x53774, x53779;
  wire x53783, x53788, x53794, x53795, x53798, x53800, x53805, x53806;
  wire x53809, x53811, x53814, x53819, x53823, x53828, x53834, x53835;
  wire x53838, x53840, x53845, x53846, x53849, x53851, x53854, x53856;
  wire x53860, x53864, x53869, x53873, x53876, x53877, x53880, x53882;
  wire x53887, x53888, x53891, x53893, x53896, x53898, x53902, x53906;
  wire x53911, x53915, x53918, x53919, x53922, x53924, x53929, x53930;
  wire x53933, x53935, x53938, x53941, x53947, x53951, x53956, x53960;
  wire x53963, x53964, x53967, x53969, x53974, x53975, x53978, x53980;
  wire x53983, x53986, x53987, x53993, x53997, x54002, x54006, x54012;
  wire x54013, x54016, x54018, x54021, x54024, x54025, x54028, x54030;
  wire x54033, x54036, x54037, x54043, x54047, x54052, x54056, x54062;
  wire x54063, x54066, x54068, x54071, x54074, x54075, x54078, x54080;
  wire x54083, x54086, x54087, x54090, x54094, x54099, x54103, x54108;
  wire x54112, x54118, x54119, x54122, x54124, x54127, x54130, x54131;
  wire x54134, x54136, x54139, x54142, x54143, x54146, x54148, x54151;
  wire x54156, x54160, x54165, x54169, x54174, x54178, x54181, x54182;
  wire x54185, x54187, x54190, x54193, x54194, x54197, x54199, x54202;
  wire x54205, x54206, x54209, x54211, x54214, x54219, x54223, x54228;
  wire x54232, x54237, x54241, x54244, x54245, x54248, x54250, x54253;
  wire x54256, x54257, x54260, x54262, x54265, x54268, x54269, x54272;
  wire x54274, x54277, x54282, x54286, x54290, x54295, x54299, x54304;
  wire x54308, x54311, x54312, x54315, x54317, x54320, x54323, x54324;
  wire x54327, x54329, x54332, x54335, x54336, x54339, x54341, x54344;
  wire x54346, x54350, x54354, x54358, x54363, x54367, x54372, x54376;
  wire x54379, x54380, x54383, x54385, x54388, x54390, x54391, x54394;
  wire x54396, x54399, x54401, x54402, x54405, x54407, x54410, x54411;
  wire x54415, x54419, x54423, x54427, x54431, x54435, x54439, x54443;
  wire x54447, x54451, x54455, x54459, x54463, x54464, x54468, x54469;
  wire x54470, x54474, x54475, x54476, x54480, x54484, x54485, x54486;
  wire x54490, x54494, x54495, x54496, x54500, x54504, x54505, x54506;
  wire x54510, x54514, x54516, x54519, x54523, x54527, x54529, x54532;
  wire x54536, x54540, x54544, x54546, x54549, x54553, x54557, x54561;
  wire x54563, x54564, x54567, x54571, x54575, x54579, x54581, x54582;
  wire x54585, x54587, x54590, x54594, x54598, x54600, x54601, x54604;
  wire x54606, x54609, x54613, x54617, x54621, x54624, x54625, x54628;
  wire x54630, x54633, x54637, x54641, x54645, x54651, x54652, x54655;
  wire x54657, x54660, x54664, x54668, x54672, x54678, x54679, x54682;
  wire x54684, x54687, x54691, x54695, x54699, x54705, x54706, x54709;
  wire x54713, x54715, x54717, x54720, x54724, x54728, x54732, x54738;
  wire x54739, x54742, x54746, x54748, x54750, x54753, x54757, x54761;
  wire x54766, x54770, x54776, x54777, x54780, x54784, x54786, x54788;
  wire x54791, x54795, x54799, x54804, x54808, x54814, x54815, x54818;
  wire x54820, x54823, x54825, x54827, x54830, x54834, x54838, x54843;
  wire x54847, x54853, x54854, x54857, x54859, x54862, x54864, x54866;
  wire x54869, x54871, x54874, x54878, x54883, x54887, x54893, x54894;
  wire x54897, x54899, x54902, x54904, x54906, x54909, x54911, x54914;
  wire x54918, x54923, x54927, x54933, x54934, x54937, x54939, x54942;
  wire x54945, x54948, x54950, x54953, x54956, x54959, x54963, x54968;
  wire x54972, x54977, x54981, x54984, x54985, x54988, x54990, x54993;
  wire x54995, x54998, x55000, x55003, x55005, x55008, x55012, x55016;
  wire x55020, x55024, x55028, x55038, x55042, x55049, x55056, x55060;
  wire x55068, x55072, x55080, x55084, x55092, x55096, x55104, x55108;
  wire x55113, x55117, x55121, x55126, x55130, x55134, x55139, x55143;
  wire x55147, x55152, x55156, x55160, x55165, x55169, x55173, x55177;
  wire x55182, x55186, x55191, x55195, x55199, x55204, x55208, x55213;
  wire x55217, x55221, x55226, x55230, x55235, x55239, x55243, x55248;
  wire x55252, x55257, x55261, x55265, x55270, x55274, x55276, x55280;
  wire x55284, x55288, x55293, x55297, x55300, x55303, x55307, x55312;
  wire x55316, x55321, x55325, x55328, x55331, x55335, x55340, x55344;
  wire x55349, x55353, x55356, x55359, x55363, x55368, x55372, x55375;
  wire x55378, x55382, x55385, x55388, x55392, x55397, x55401, x55404;
  wire x55407, x55409, x55412, x55415, x55418, x55422, x55427, x55431;
  wire x55434, x55437, x55439, x55442, x55445, x55448, x55452, x55457;
  wire x55461, x55464, x55467, x55469, x55472, x55475, x55478, x55482;
  wire x55487, x55491, x55494, x55497, x55499, x55502, x55505, x55508;
  wire x55512, x55517, x55521, x55524, x55527, x55529, x55532, x55535;
  wire x55538, x55542, x55547, x55551, x55554, x55555, x55558, x55560;
  wire x55563, x55565, x55566, x55569, x55573, x55577, x55581, x55594;
  wire x55599, x55602, x55607, x55610, x55615, x55618, x55623, x55626;
  wire x55631, x55634, x55638, x55642, x55645, x55648, x55652, x55656;
  wire x55659, x55662, x55666, x55670, x55673, x55676, x55680, x55684;
  wire x55687, x55690, x55694, x55698, x55703, x55705, x55708, x55713;
  wire x55717, x55720, x55723, x55725, x55728, x55733, x55737, x55740;
  wire x55743, x55745, x55748, x55753, x55757, x55760, x55763, x55765;
  wire x55768, x55773, x55777, x55780, x55783, x55785, x55788, x55793;
  wire x55797, x55800, x55803, x55805, x55808, x55813, x55817, x55820;
  wire x55821, x55824, x55826, x55829, x55834, x55838, x55841, x55842;
  wire x55845, x55847, x55850, x55855, x55859, x55862, x55863, x55866;
  wire x55868, x55871, x55876, x55880, x55883, x55884, x55887, x55889;
  wire x55892, x55897, x55901, x55904, x55905, x55908, x55910, x55913;
  wire x55918, x55922, x55925, x55926, x55929, x55931, x55934, x55939;
  wire x55943, x55946, x55947, x55950, x55952, x55955, x55960, x55964;
  wire x55967, x55968, x55971, x55973, x55976, x55981, x55985, x55988;
  wire x55989, x55992, x55994, x55997, x56001, x56005, x56012, x56016;
  wire x56020, x56024, x56029, x56033, x56038, x56042, x56047, x56051;
  wire x56056, x56060, x56065, x56066, x56068, x56071, x56075, x56080;
  wire x56081, x56083, x56086, x56090, x56095, x56096, x56098, x56101;
  wire x56105, x56110, x56111, x56113, x56116, x56120, x56125, x56126;
  wire x56128, x56131, x56135, x56140, x56141, x56143, x56144, x56147;
  wire x56151, x56156, x56157, x56159, x56160, x56163, x56167, x56172;
  wire x56173, x56175, x56176, x56179, x56183, x56188, x56189, x56191;
  wire x56192, x56195, x56199, x56204, x56205, x56207, x56208, x56211;
  wire x56215, x56220, x56221, x56223, x56224, x56227, x56231, x56236;
  wire x56237, x56239, x56240, x56243, x56247, x56252, x56253, x56255;
  wire x56256, x56259, x56263, x56268, x56269, x56271, x56272, x56275;
  wire x56279, x56284, x56285, x56287, x56288, x56291, x56295, x56300;
  wire x56301, x56303, x56304, x56307, x56311, x56316, x56317, x56319;
  wire x56320, x56323, x56327, x56332, x56333, x56335, x56336, x56339;
  wire x56343, x56348, x56349, x56351, x56352, x56355, x56359, x56363;
  wire x56373, x56377, x56378, x56382, x56383, x56387, x56388, x56392;
  wire x56393, x56397, x56399, x56402, x56406, x56409, x56412, x56416;
  wire x56419, x56422, x56426, x56429, x56432, x56436, x56439, x56442;
  wire x56446, x56449, x56452, x56456, x56459, x56462, x56466, x56469;
  wire x56472, x56476, x56479, x56482, x56486, x56489, x56492, x56496;
  wire x56499, x56502, x56506, x56509, x56512, x56516, x56519, x56522;
  wire x56526, x56529, x56532, x56536, x56539, x56542, x56546, x56549;
  wire x56552, x56556, x56559, x56562, x56566, x56569, x56572, x56576;
  wire x56579, x56582, x56586, x56590, x56598, x56602, x56606, x56610;
  wire x56615, x56619, x56624, x56628, x56633, x56637, x56642, x56646;
  wire x56651, x56655, x56660, x56664, x56667, x56670, x56674, x56677;
  wire x56680, x56684, x56687, x56690, x56694, x56697, x56700, x56704;
  wire x56707, x56710, x56714, x56717, x56720, x56724, x56727, x56730;
  wire x56734, x56737, x56740, x56744, x56747, x56750, x56754, x56757;
  wire x56760, x56764, x56767, x56770, x56774, x56777, x56780, x56784;
  wire x56787, x56790, x56794, x56797, x56800, x56804, x56807, x56810;
  wire x56814, x56817, x56820, x56824, x56827, x56830, x56834, x56837;
  wire x56840, x56844, x56846, x56852, x56856, x56858, x56861, x56863;
  wire x56866, x56868, x56871, x56873, x56876, x56878, x56881, x56883;
  wire x56886, x56888, x56891, x56893, x56896, x56898, x56901, x56903;
  wire x56906, x56908, x56911, x56913, x56916, x56918, x56921, x56923;
  wire x56926, x56928, x56931, x56933, x56936, x56938, x56941, x56943;
  wire x56946, x56948, x56951, x56953, x56956, x56958, x56961, x56963;
  wire x56966, x56968, x56971, x56973, x56976, x56977, x56978, x56979;
  wire x56980, x56981, x56982, x56983, x56984, x56985, x56986, x56987;
  wire x56988, x56989, x56990, x56991, x56992, x56993, x56994, x56995;
  wire x56996, x56997, x56998, x56999, x57000, x57001, x57007, x57011;
  wire x57015, x57019, x57023, x57027, x57031, x57035, x57039, x57043;
  wire x57047, x57051, x57055, x57059, x57063, x57067, x57071, x57075;
  wire x57079, x57083, x57087, x57091, x57095, x57099, x57100, x57102;
  wire x57105, x57108, x57111, x57113, x57116, x57118, x57121, x57123;
  wire x57126, x57128, x57131, x57133, x57136, x57138, x57141, x57143;
  wire x57146, x57148, x57151, x57153, x57156, x57158, x57161, x57163;
  wire x57166, x57168, x57171, x57173, x57176, x57178, x57181, x57183;
  wire x57186, x57188, x57191, x57193, x57196, x57198, x57201, x57203;
  wire x57206, x57208, x57211, x57213, x57216, x57217, x57218, x57220;
  wire x57223, x57226, x57229, x57232, x57235, x57237, x57240, x57242;
  wire x57245, x57247, x57250, x57252, x57255, x57257, x57260, x57262;
  wire x57265, x57267, x57270, x57272, x57275, x57277, x57280, x57282;
  wire x57285, x57287, x57290, x57292, x57295, x57297, x57300, x57302;
  wire x57305, x57307, x57310, x57312, x57315, x57317, x57320, x57321;
  wire x57322, x57323, x57324, x57326, x57329, x57332, x57335, x57338;
  wire x57341, x57344, x57347, x57350, x57353, x57355, x57358, x57360;
  wire x57363, x57365, x57368, x57370, x57373, x57375, x57378, x57380;
  wire x57383, x57385, x57388, x57390, x57393, x57395, x57398, x57399;
  wire x57400, x57401, x57402, x57403, x57404, x57406, x57409, x57412;
  wire x57415, x57418, x57421, x57424, x57427, x57430, x57433, x57437;
  wire x57441, x57445, x57449, x57453, x57457, x57461, x57465, x57467;
  wire x57470, x57472, x57475, x57479, x57483, x57487, x57491, x57495;
  wire x57499, x57501, x57504, x57506, x57509, x57511, x57514, x57516;
  wire x57519, x57521, x57524, x57526, x57529, x57531, x57534, x57536;
  wire x57539, x57541, x57544, x57546, x57549, x57551, x57553, x57555;
  wire x57557, x57559, x57561, x57563, x57565, x57567, x57569, x57571;
  wire x57573, x57575, x57577, x57579, x57581, x57583, x57585, x57587;
  wire x57589, x57591, x57593, x57595, x57597, x57599, x57601, x57603;
  wire x57605, x57607, x57609, x57612, x57614, x57616, x57618, x57620;
  wire x57622, x57624, x57626, x57628, x57630, x57632, x57634, x57636;
  wire x57638, x57640, x57642, x57644, x57646, x57648, x57650, x57652;
  wire x57654, x57656, x57658, x57660, x57662, x57664, x57666, x57671;
  wire x57673, x57675, x57677, x57679, x57681, x57683, x57685, x57687;
  wire x57689, x57691, x57693, x57695, x57697, x57699, x57701, x57703;
  wire x57705, x57707, x57709, x57711, x57713, x57715, x57717, x57727;
  wire x57729, x57731, x57733, x57735, x57737, x57739, x57741, x57743;
  wire x57745, x57747, x57749, x57751, x57753, x57755, x57773, x57777;
  wire x57781, x57785, x57789, x57793, x57797, x57801, x57805, x57809;
  wire x57813, x57817, x57821, x57825, x57829, x57833, x57837, x57841;
  wire x57845, x57849, x57853, x57857, x57861, x57865, x57869, x57873;
  wire x57877, x57881, x57885, x57889, x57893, x57894, x57896, x57898;
  wire x57900, x57902, x57904, x57906, x57908, x57910, x57912, x57914;
  wire x57916, x57918, x57920, x57922, x57924, x57926, x57960, x57962;
  wire x57964, x57966, x57968, x57970, x57972, x57974, x57976, x57978;
  wire x57980, x57982, x57984, x57986, x57988, x57990, x57992, x57994;
  wire x57996, x57998, x58000, x58002, x58004, x58006, x58008, x58010;
  wire x58012, x58014, x58016, x58018, x58020, x58022, x60842, x60843;
  wire x60844, x60846, x60847, x60849, x60850, x60852, x60853, x60855;
  wire x60856, x60858, x60859, x60861, x60862, x60864, x60865, x60867;
  wire x60868, x60870, x60871, x60873, x60874, x60876, x60877, x60879;
  wire x60880, x60882, x60883, x60885, x60886, x60888, x60889, x60891;
  wire x60892, x60894, x60895, x60897, x60898, x60900, x60901, x60903;
  wire x60904, x60906, x60907, x60909, x60910, x60912, x60913, x60915;
  wire x60916, x60918, x60919, x60921, x60922, x60924, x60925, x60927;
  wire x60928, x60930, x60931, x60933, x60934, x60937, x60938, x60939;
  wire x60942, x60943, x60944, x60955, x60962, x60967, x60970, x60977;
  wire x60978, x60980, x60981, x60983, x60984, x60986, x60987, x60989;
  wire x60990, x60992, x60993, x60995, x60996, x60998, x60999, x61001;
  wire x61002, x61004, x61005, x61007, x61008, x61010, x61011, x61013;
  wire x61014, x61016, x61017, x61019, x61020, x61022, x61023, x61025;
  wire x61026, x61028, x61029, x61031, x61032, x61034, x61035, x61037;
  wire x61038, x61040, x61041, x61043, x61044, x61046, x61047, x61049;
  wire x61050, x61052, x61053, x61055, x61056, x61058, x61059, x61061;
  wire x61062, x61064, x61065, x61067, x61068, x61071, x61072, x61073;
  wire x61076, x61077, x61106, x61107, x61109, x61110, x61112, x61113;
  wire x61115, x61116, x61118, x61119, x61121, x61122, x61124, x61125;
  wire x61127, x61128, x61130, x61131, x61133, x61134, x61136, x61137;
  wire x61139, x61140, x61142, x61143, x61145, x61146, x61148, x61149;
  wire x61151, x61152, x61154, x61155, x61157, x61158, x61160, x61161;
  wire x61163, x61164, x61166, x61167, x61169, x61170, x61172, x61173;
  wire x61175, x61176, x61178, x61179, x61181, x61182, x61184, x61185;
  wire x61187, x61188, x61190, x61191, x61193, x61194, x61196, x61197;
  wire x61200, x61201, x61202, x61205, x61206, x61235, x61236, x61238;
  wire x61239, x61241, x61242, x61244, x61245, x61247, x61248, x61250;
  wire x61251, x61253, x61254, x61256, x61257, x61259, x61260, x61262;
  wire x61263, x61265, x61266, x61268, x61269, x61271, x61272, x61274;
  wire x61275, x61277, x61278, x61280, x61281, x61283, x61284, x61286;
  wire x61287, x61289, x61290, x61292, x61293, x61295, x61296, x61298;
  wire x61299, x61301, x61302, x61304, x61305, x61307, x61308, x61310;
  wire x61311, x61313, x61314, x61316, x61317, x61319, x61320, x61322;
  wire x61323, x61325, x61326, x61329, x61330, x61331, x61334, x61335;
  wire x61425, x61427, x61686, x61975, x62931, x62933, x63027, x63028;
  wire x63032, x63033, x63036, x63038, x63039, x63042, x63044, x63045;
  wire x63048, x63050, x63051, x63054, x63056, x63057, x63060, x63062;
  wire x63063, x63066, x63068, x63069, x63072, x63074, x63075, x63078;
  wire x63080, x63081, x63084, x63086, x63087, x63090, x63092, x63093;
  wire x63096, x63098, x63099, x63102, x63104, x63105, x63108, x63110;
  wire x63111, x63114, x63116, x63117, x63120, x63122, x63123, x63126;
  wire x63128, x63129, x63132, x63134, x63135, x63138, x63140, x63141;
  wire x63144, x63146, x63147, x63150, x63152, x63153, x63156, x63158;
  wire x63159, x63162, x63164, x63165, x63168, x63170, x63171, x63174;
  wire x63176, x63177, x63180, x63182, x63183, x63186, x63188, x63189;
  wire x63192, x63194, x63195, x63198, x63200, x63201, x63204, x63206;
  wire x63207, x63210, x63211, x63212, x63213, x63214, x63215, x63216;
  wire x63217, x63218, x63219, x63220, x63221, x63222, x63223, x63224;
  wire x63225, x63226, x63227, x63228, x63229, x63230, x63231, x63232;
  wire x63233, x63234, x63235, x63236, x63237, x63238, x63239, x63245;
  wire x63249, x63253, x63257, x63261, x63265, x63269, x63273, x63277;
  wire x63281, x63285, x63289, x63293, x63297, x63301, x63305, x63309;
  wire x63313, x63317, x63321, x63325, x63329, x63333, x63337, x63341;
  wire x63345, x63349, x63353, x63354, x63356, x63359, x63362, x63365;
  wire x63367, x63370, x63372, x63375, x63377, x63380, x63382, x63385;
  wire x63387, x63390, x63392, x63395, x63397, x63400, x63402, x63405;
  wire x63407, x63410, x63412, x63415, x63417, x63420, x63422, x63425;
  wire x63427, x63430, x63432, x63435, x63437, x63440, x63442, x63445;
  wire x63447, x63450, x63452, x63455, x63457, x63460, x63462, x63465;
  wire x63467, x63470, x63472, x63475, x63477, x63480, x63482, x63485;
  wire x63487, x63490, x63491, x63493, x63496, x63499, x63502, x63505;
  wire x63508, x63510, x63513, x63515, x63518, x63520, x63523, x63525;
  wire x63528, x63530, x63533, x63535, x63538, x63540, x63543, x63545;
  wire x63548, x63550, x63553, x63555, x63558, x63560, x63563, x63565;
  wire x63568, x63570, x63573, x63575, x63578, x63580, x63583, x63585;
  wire x63588, x63590, x63593, x63595, x63598, x63600, x63603, x63605;
  wire x63608, x63610, x63613, x63614, x63616, x63619, x63622, x63625;
  wire x63628, x63631, x63634, x63637, x63640, x63643, x63645, x63648;
  wire x63650, x63653, x63655, x63658, x63660, x63663, x63665, x63668;
  wire x63670, x63673, x63675, x63678, x63680, x63683, x63685, x63688;
  wire x63690, x63693, x63695, x63698, x63700, x63703, x63705, x63708;
  wire x63709, x63711, x63714, x63717, x63720, x63723, x63726, x63729;
  wire x63732, x63735, x63738, x63741, x63744, x63747, x63750, x63757;
  wire x63759, x63762, x63766, x63768, x63771, x63773, x63776, x63778;
  wire x63781, x63785, x63787, x63790, x63792, x63796, x63800, x63804;
  wire x63808, x63812, x63819, x63823, x63827, x63831, x63835, x63839;
  wire x63843, x63847, x63851, x63855, x63859, x63863, x63867, x63871;
  wire x63875, x63914, x64009, x64102, x64191, x64272, x64337, x64339;
  wire x64341, x64343, x64345, x64347, x64349, x64351, x64353, x64355;
  wire x64357, x64359, x64361, x64363, x64365, x64367, x64369, x64371;
  wire x64373, x64375, x64377, x64379, x64381, x64383, x64385, x64387;
  wire x64389, x64391, x64393, x64395, x64397, x64429, x64433, x64436;
  wire x64438, x64441, x64443, x64446, x64448, x64451, x64453, x64456;
  wire x64458, x64461, x64463, x64466, x64468, x64471, x64473, x64476;
  wire x64477, x64478, x64479, x64480, x64481, x64482, x64483, x64484;
  wire x64490, x64494, x64498, x64502, x64506, x64510, x64514, x64515;
  wire x64517, x64520, x64523, x64526, x64528, x64531, x64533, x64536;
  wire x64538, x64541, x64543, x64546, x64547, x64549, x64552, x64555;
  wire x64558, x64561, x64564, x64565, x64567, x64574, x64576, x64579;
  wire x64583, x64585, x64588, x64590, x64593, x64595, x64598, x64602;
  wire x64604, x64607, x64646, x64741, x64834, x64923, x65004, x65099;
  wire x65103, x65106, x65108, x65111, x65113, x65116, x65118, x65121;
  wire x65123, x65126, x65128, x65131, x65133, x65136, x65138, x65141;
  wire x65143, x65146, x65147, x65148, x65149, x65150, x65151, x65152;
  wire x65153, x65154, x65160, x65164, x65168, x65172, x65176, x65180;
  wire x65184, x65185, x65187, x65190, x65193, x65196, x65198, x65201;
  wire x65203, x65206, x65208, x65211, x65213, x65216, x65217, x65219;
  wire x65222, x65225, x65228, x65231, x65234, x65235, x65237, x65244;
  wire x65246, x65249, x65253, x65255, x65258, x65260, x65263, x65265;
  wire x65268, x65272, x65274, x65277, x65316, x65411, x65504, x65593;
  wire x65674, x65769, x65773, x65776, x65778, x65781, x65783, x65786;
  wire x65788, x65791, x65793, x65796, x65798, x65801, x65803, x65806;
  wire x65808, x65811, x65813, x65816, x65817, x65818, x65819, x65820;
  wire x65821, x65822, x65823, x65824, x65830, x65834, x65838, x65842;
  wire x65846, x65850, x65854, x65855, x65857, x65860, x65863, x65866;
  wire x65868, x65871, x65873, x65876, x65878, x65881, x65883, x65886;
  wire x65887, x65889, x65892, x65895, x65898, x65901, x65904, x65905;
  wire x65907, x65914, x65916, x65919, x65923, x65925, x65928, x65930;
  wire x65933, x65935, x65938, x65942, x65944, x65947, x65986, x66081;
  wire x66174, x66263, x66344, x66409, x66470, x66472, x66603, x67463;
  wire x67465, x67596, x68458, x68459, x68461, x68464, x68467, x68469;
  wire x68470, x68471, x68473, x68475, x68478, x68480, x68483, x68485;
  wire x68488, x68491, x68494, x68498, x68501, x68502, x68505, x68509;
  wire x68511, x68514, x68516, x68519, x68521, x68524, x68526, x68529;
  wire x68530, x68533, x68535, x68537, x68541, x68545, x68549, x68553;
  wire x68557, x68561, x68563, x68570, x68624, x68625, x68626, x68627;
  wire x68628, x68629, x68639, x68640, x68641, x68643, x68654, x68655;
  wire x68656, x68658, x68660, x68661, x68662, x68663, x68671, x68677;
  wire x68679, x68681, x68682, x68683, x68684, x68692, x68698, x68700;
  wire x68702, x68703, x68720, x68721, x68745, x68810, x71027, x71028;
  wire x71032, x71033, x71037, x71038, x71042, x71043, x71047, x71048;
  wire x71052, x71053, x71057, x71059, x71061, x71063, x71065, x71067;
  wire x71069, x71071, x71073, x71075, x71077, x71078, x71082, x71083;
  wire x71087, x71088, x71092, x71093, x71097, x71098, x71102, x71103;
  wire x71107, x71109, x71111, x71113, x71115, x71117, x71119, x71121;
  wire x71123, x71125, x71126, x71127, x71132, x71133, x71135, x71136;
  wire x71138, x71139, x83383, x83384, x83385, x83386, x83387, x83388;
  wire x83389, x83390, x83391, x83392, x83393, x83394, x83395, x83396;
  wire x83397, x83398, x83399, x83400, x83401, x83402, x83403, x83404;
  wire x83405, x83406, x83407, x83408, x83409, x83410, x83411, x83412;
  wire x83413, x83414, x83415, x83416, x83417, x83418, x83419, x83420;
  wire x83421, x83422, x83423, x83424, x83425, x83426, x83427, x83428;
  wire x83429, x83430, x83431, x83432, x83433, x83434, x83435, x83436;
  wire x83437, x83438, x83439, x83440, x83441, x83442, x83443, x83444;
  wire x83445, x83446, x83447, x83448, x83449, x83450, x83451, x83452;
  wire x83453, x83454, x83455, x83456, x83457, x83458, x83459, x83460;
  wire x83461, x83462, x83463, x83464, x83465, x83466, x83467, x83468;
  wire x83469, x83470, x83471, x83472, x83473, x83474, x83475, x83476;
  wire x83477, x83478, x83479, x83480, x83481, x83482, x83483, x83484;
  wire x83485, x83486, x83487, x83488, x83489, x83490, x83491, x83492;
  wire x83493, x83494, x83495, x83496, x83497, x83498, x83499, x83500;
  wire x83501, x83502, x83503, x83504, x83505, x83506, x83507, x83508;
  wire x83509, x83510, x83511, x83512, x83513, x83514, x83515, x83516;
  wire x83517, x83518, x83519, x83520, x83521, x83522, x83523, x83524;
  wire x83525, x83526, x83527, x83528, x83529, x83530, x83531, x83532;
  wire x83533, x83534, x83535, x83536, x83537, x83538, x83539, x83540;
  wire x83541, x83542, x83543, x83544, x83545, x83546, x83547, x83548;
  wire x83549, x83550, x83551, x83552, x83553, x83554, x83555, x83556;
  wire x83557, x83558, x83559, x83560, x83561, x83562, x83563, x83564;
  wire x83565, x83566, x83567, x83568, x83569, x83570, x83571, x83572;
  wire x83573, x83574, x83575, x83576, x83577, x83578, x83579, x83580;
  wire x83581, x83582, x83583, x83584, x83585, x83586, x83587, x83588;
  wire x83589, x83590, x83591, x83592, x83593, x83594, x83595, x83596;
  wire x83597, x83598, x83599, x83600, x83601, x83602, x83603, x83604;
  wire x83605, x83606, x83607, x83608, x83609, x83610, x83611, x83612;
  wire x83613, x83614, x83615, x83616, x83617, x83618, x83619, x83620;
  wire x83621, x83622, x83623, x83624, x83625, x83626, x83627, x83628;
  wire x83629, x83630, x83631, x83632, x83633, x83634, x83635, x83636;
  wire x83637, x83638, x83639, x83640, x83641, x83642, x83643, x83644;
  wire x83645, x83646, x83647, x83648, x83649, x83650, x83651, x83652;
  wire x83653, x83654, x83655, x83656, x83657, x83658, x83659, x83660;
  wire x83661, x83662, x83663, x83664, x83665, x83666, x83667, x83668;
  wire x83669, x83670, x83671, x83672, x83673, x83674, x83675, x83676;
  wire x83677, x83678, x83679, x83680, x83681, x83682, x83683, x83684;
  wire x83685, x83686, x83687, x83688, x83689, x83690, x83691, x83692;
  wire x83693, x83694, x83695, x83696, x83697, x83698, x83699, x83700;
  wire x83701, x83702, x83703, x83704, x83705, x83706, x83707, x83708;
  wire x83709, x83710, x83711, x83712, x83713, x83714, x83715, x83716;
  wire x83717, x83718, x83719, x83720, x83721, x83722, x83723, x83724;
  wire x83725, x83726, x83727, x83728, x83729, x83730, x83731, x83732;
  wire x83733, x83734, x83735, x83736, x83737, x83738, x83739, x83740;
  wire x83741, x83742, x83743, x83744, x83745, x83746, x83747, x83748;
  wire x83749, x83750, x83751, x83752, x83753, x83754, x83755, x83756;
  wire x83757, x83758, x83759, x83760, x83761, x83762, x83763, x83764;
  wire x83765, x83766, x83767, x83768, x83769, x83770, x83771, x83772;
  wire x83773, x83774, x83775, x83776, x83777, x83778, x83779, x83780;
  wire x83781, x83782, x83783, x83784, x83785, x83786, x83787, x83788;
  wire x83789, x83790, x83791, x83792, x83793, x83794, x83795, x83796;
  wire x83797, x83798, x83799, x83800, x83801, x83802, x83803, x83804;
  wire x83805, x83806, x83807, x83808, x83809, x83810, x83811, x83812;
  wire x83813, x83814, x83815, x83816, x83817, x83818, x83819, x83820;
  wire x83821, x83822, x83823, x83824, x83825, x83826, x83827, x83828;
  wire x83829, x83830, x83831, x83832, x83833, x83834, x83835, x83836;
  wire x83837, x83838, x83839, x83840, x83841, x83842, x83843, x83844;
  wire x83845, x83846, x83847, x83848, x83849, x83850, x83851, x83852;
  wire x83853, x83854, x83855, x83856, x83857, x83858, x83859, x83860;
  wire x83861, x83862, x83863, x83864, x83865, x83866, x83867, x83868;
  wire x83869, x83870, x83871, x83872, x83873, x83874, x83875, x83876;
  wire x83877, x83878, x83879, x83880, x83881, x83882, x83883, x83884;
  wire x83885, x83886, x83887, x83888, x83889, x83890, x83891, x83892;
  wire x83893, x83894, x83895, x83896, x83897, x83898, x83899, x83900;
  wire x83901, x83902, x83903, x83904, x83905, x83906, x83907, x83908;
  wire x83909, x83910, x83911, x83912, x83913, x83914, x83915, x83916;
  wire x83917, x83918, x83919, x83920, x83921, x83922, x83923, x83924;
  wire x83925, x83926, x83927, x83928, x83929, x83930, x83931, x83932;
  wire x83933, x83934, x83935, x83936, x83937, x83938, x83939, x83940;
  wire x83941, x83942, x83943, x83944, x83945, x83946, x83947, x83948;
  wire x83949, x83950, x83951, x83952, x83953, x83954, x83955, x83956;
  wire x83957, x83958, x83959, x83960, x83961, x83962, x83963, x83964;
  wire x83965, x83966, x83967, x83968, x83969, x83970, x83971, x83972;
  wire x83973, x83974, x83975, x83976, x83977, x83978, x83979, x83980;
  wire x83981, x83982, x83983, x83984, x83985, x83986, x83987, x83988;
  wire x83989, x83990, x83991, x83992, x83993, x83994, x83995, x83996;
  wire x83997, x83998, x83999, x84000, x84001, x84002, x84003, x84004;
  wire x84005, x84006, x84007, x84008, x84009, x84010, x84011, x84012;
  wire x84013, x84014, x84015, x84016, x84017, x84018, x84019, x84020;
  wire x84021, x84022, x84023, x84024, x84025, x84026, x84027, x84028;
  wire x84029, x84030, x84031, x84032, x84033, x84034, x84035, x84036;
  wire x84037, x84038, x84039, x84040, x84041, x84042, x84043, x84044;
  wire x84045, x84046, x84047, x84048, x84049, x84050, x84051, x84052;
  wire x84053, x84054, x84055, x84056, x84057, x84058, x84059, x84060;
  wire x84061, x84062, x84063, x84064, x84065, x84066, x84067, x84068;
  wire x84069, x84070, x84071, x84072, x84073, x84074, x84075, x84076;
  wire x84077, x84078, x84079, x84080, x84081, x84082, x84083, x84084;
  wire x84085, x84086, x84087, x84088, x84089, x84090, x84091, x84092;
  wire x84093, x84094, x84095, x84096, x84097, x84098, x84099, x84100;
  wire x84101, x84102, x84103, x84104, x84105, x84106, x84107, x84108;
  wire x84109, x84110, x84111, x84112, x84113, x84114, x84115, x84116;
  wire x84117, x84118, x84119, x84120, x84121, x84122, x84123, x84124;
  wire x84125, x84126, x84127, x84128, x84129, x84130, x84131, x84132;
  wire x84133, x84134, x84135, x84136, x84137, x84138, x84139, x84140;
  wire x84141, x84142, x84143, x84144, x84145, x84146, x84147, x84148;
  wire x84149, x84150, x84151, x84152, x84153, x84154, x84155, x84156;
  wire x84157, x84158, x84159, x84160, x84161, x84162, x84163, x84164;
  wire x84165, x84166, x84167, x84168, x84169, x84170, x84171, x84172;
  wire x84173, x84174, x84175, x84176, x84177, x84178, x84179, x84180;
  wire x84181, x84182, x84183, x84184, x84185, x84186, x84187, x84188;
  wire x84189, x84190, x84191, x84192, x84193, x84194, x84195, x84196;
  wire x84197, x84198, x84199, x84200, x84201, x84202, x84203, x84204;
  wire x84205, x84206, x84207, x84208, x84209, x84210, x84211, x84212;
  wire x84213, x84214, x84215, x84216, x84217, x84218, x84219, x84220;
  wire x84221, x84222, x84223, x84224, x84225, x84226, x84227, x84228;
  wire x84229, x84230, x84231, x84232, x84233, x84234, x84235, x84236;
  wire x84237, x84238, x84239, x84240, x84241, x84242, x84243, x84244;
  wire x84245, x84246, x84247, x84248, x84249, x84250, x84251, x84252;
  wire x84253, x84254, x84255, x84256, x84257, x84258, x84259, x84260;
  wire x84261, x84262, x84263, x84264, x84265, x84266, x84267, x84268;
  wire x84269, x84270, x84271, x84272, x84273, x84274, x84275, x84276;
  wire x84277, x84278, x84279, x84280, x84281, x84282, x84283, x84284;
  wire x84285, x84286, x84287, x84288, x84289, x84290, x84291, x84292;
  wire x84293, x84294, x84295, x84296, x84297, x84298, x84299, x84300;
  wire x84301, x84302, x84303, x84304, x84305, x84306, x84307, x84308;
  wire x84309, x84310, x84311, x84312, x84313, x84314, x84315, x84316;
  wire x84317, x84318, x84319, x84320, x84321, x84322, x84323, x84324;
  wire x84325, x84326, x84327, x84328, x84329, x84330, x84331, x84332;
  wire x84333, x84334, x84335, x84336, x84337, x84338, x84339, x84340;
  wire x84341, x84342, x84343, x84344, x84345, x84346, x84347, x84348;
  wire x84349, x84350, x84351, x84352, x84353, x84354, x84355, x84356;
  wire x84357, x84358, x84359, x84360, x84361, x84362, x84363, x84364;
  wire x84365, x84366, x84367, x84368, x84369, x84370, x84371, x84372;
  wire x84373, x84374, x84375, x84376, x84377, x84378, x84379, x84380;
  wire x84381, x84382, x84383, x84384, x84385, x84386, x84387, x84388;
  wire x84389, x84390, x84391, x84392, x84393, x84394, x84395, x84396;
  wire x84397, x84398, x84399, x84400, x84401, x84402, x84403, x84404;
  wire x84405, x84406, x84407, x84408, x84409, x84410, x84411, x84412;
  wire x84413, x84414, x84415, x84416, x84417, x84418, x84419, x84420;
  wire x84421, x84422, x84423, x84424, x84425, x84426, x84427, x84428;
  wire x84429, x84430, x84431, x84432, x84433, x84434, x84435, x84436;
  wire x84437, x84438, x84439, x84440, x84441, x84442, x84443, x84444;
  wire x84445, x84446, x84447, x84448, x84449, x84450, x84451, x84452;
  wire x84453, x84454, x84455, x84456, x84457, x84458, x84459, x84460;
  wire x84461, x84462, x84463, x84464, x84465, x84466, x84467, x84468;
  wire x84469, x84470, x84471, x84472, x84473, x84474, x84475, x84476;
  wire x84477, x84478, x84479, x84480, x84481, x84482, x84483, x84484;
  wire x84485, x84486, x84487, x84488, x84489, x84490, x84491, x84492;
  wire x84493, x84494, x84495, x84496, x84497, x84498, x84499, x84500;
  wire x84501, x84502, x84503, x84504, x84505, x84506, x84507, x84508;
  wire x84509, x84510, x84511, x84512, x84513, x84514, x84515, x84516;
  wire x84517, x84518, x84519, x84520, x84521, x84522, x84523, x84524;
  wire x84525, x84526, x84527, x84528, x84529, x84530, x84531, x84532;
  wire x84533, x84534, x84535, x84536, x84537, x84538, x84539, x84540;
  wire x84541, x84542, x84543, x84544, x84545, x84546, x84547, x84548;
  wire x84549, x84550, x84551, x84552, x84553, x84554, x84555, x84556;
  wire x84557, x84558, x84559, x84560, x84561, x84562, x84563, x84564;
  wire x84565, x84566, x84567, x84568, x84569, x84570, x84571, x84572;
  wire x84573, x84574, x84575, x84576, x84577, x84578, x84579, x84580;
  wire x84581, x84582, x84583, x84584, x84585, x84586, x84587, x84588;
  wire x84589, x84590, x84591, x84592, x84593, x84594, x84595, x84596;
  wire x84597, x84598, x84599, x84600, x84601, x84602, x84603, x84604;
  wire x84605, x84606, x84607, x84608, x84609, x84610, x84611, x84612;
  wire x84613, x84614, x84615, x84616, x84617, x84618, x84619, x84620;
  wire x84621, x84622, x84623, x84624, x84625, x84626, x84627, x84628;
  wire x84629, x84630, x84631, x84632, x84633, x84634, x84635, x84636;
  wire x84637, x84638, x84639, x84640, x84641, x84642, x84643, x84644;
  wire x84645, x84646, x84647, x84648, x84649, x84650, x84651, x84652;
  wire x84653, x84654, x84655, x84656, x84657, x84658, x84659, x84660;
  wire x84661, x84662, x84663, x84664, x84665, x84666, x84667, x84668;
  wire x84669, x84670, x84671, x84672, x84673, x84674, x84675, x84676;
  wire x84677, x84678, x84679, x84680, x84681, x84682, x84683, x84684;
  wire x84685, x84686, x84687, x84688, x84689, x84690, x84691, x84692;
  wire x84693, x84694, x84695, x84696, x84697, x84698, x84699, x84700;
  wire x84701, x84702, x84703, x84704, x84705, x84706, x84707, x84708;
  wire x84709, x84710, x84711, x84712, x84713, x84714, x84715, x84716;
  wire x84717, x84718, x84719, x84720, x84721, x84722, x84723, x84724;
  wire x84725, x84726, x84727, x84728, x84729, x84730, x84731, x84732;
  wire x84733, x84734, x84735, x84736, x84737, x84738, x84739, x84740;
  wire x84741, x84742, x84743, x84744, x84745, x84746, x84747, x84748;
  wire x84749, x84750, x84751, x84752, x84753, x84754, x84755, x84756;
  wire x84757, x84758, x84759, x84760, x84761, x84762, x84763, x84764;
  wire x84765, x84766, x84767, x84768, x84769, x84770, x84771, x84772;
  wire x84773, x84774, x84775, x84776, x84777, x84778, x84779, x84780;
  wire x84781, x84782, x84783, x84784, x84785, x84786, x84787, x84788;
  wire x84789, x84790, x84791, x84792, x84793, x84794, x84795, x84796;
  wire x84797, x84798, x84799, x84800, x84801, x84802, x84803, x84804;
  wire x84805, x84806, x84807, x84808, x84809, x84810, x84811, x84812;
  wire x84813, x84814, x84815, x84816, x84817, x84818, x84819, x84820;
  wire x84821, x84822, x84823, x84824, x84825, x84826, x84827, x84828;
  wire x84829, x84830, x84831, x84832, x84833, x84834, x84835, x84836;
  wire x84837, x84838, x84839, x84840, x84841, x84842, x84843, x84844;
  wire x84845, x84846, x84847, x84848, x84849, x84850, x84851, x84852;
  wire x84853, x84854, x84855, x84856, x84857, x84858, x84859, x84860;
  wire x84861, x84862, x84863, x84864, x84865, x84866, x84867, x84868;
  wire x84869, x84870, x84871, x84872, x84873, x84874, x84875, x84876;
  wire x84877, x84878, x84879, x84880, x84881, x84882, x84883, x84884;
  wire x84885, x84886, x84887, x84888, x84889, x84890, x84891, x84892;
  wire x84893, x84894, x84895, x84896, x84897, x84898, x84899, x84900;
  wire x84901, x84902, x84903, x84904, x84905, x84906, x84907, x84908;
  wire x84909, x84910, x84911, x84912, x84913, x84914, x84915, x84916;
  wire x84917, x84918, x84919, x84920, x84921, x84922, x84923, x84924;
  wire x84925, x84926, x84927, x84928, x84929, x84930, x84931, x84932;
  wire x84933, x84934, x84935, x84936, x84937, x84938, x84939, x84940;
  wire x84941, x84942, x84943, x84944, x84945, x84946, x84947, x84948;
  wire x84949, x84950, x84951, x84952, x84953, x84954, x84955, x84956;
  wire x84957, x84958, x84959, x84960, x84961, x84962, x84963, x84964;
  wire x84965, x84966, x84967, x84968, x84969, x84970, x84971, x84972;
  wire x84973, x84974, x84975, x84976, x84977, x84978, x84979, x84980;
  wire x84981, x84982, x84983, x84984, x84985, x84986, x84987, x84988;
  wire x84989, x84990, x84991, x84992, x84993, x84994, x84995, x84996;
  wire x84997, x84998, x84999, x85000, x85001, x85002, x85003, x85004;
  wire x85005, x85006, x85007, x85008, x85009, x85010, x85011, x85012;
  wire x85013, x85014, x85015, x85016, x85017, x85018, x85019, x85020;
  wire x85021, x85022, x85023, x85024, x85025, x85026, x85027, x85028;
  wire x85029, x85030, x85031, x85032, x85033, x85034, x85035, x85036;
  wire x85037, x85038, x85039, x85040, x85041, x85042, x85043, x85044;
  wire x85045, x85046, x85047, x85048, x85049, x85050, x85051, x85052;
  wire x85053, x85054, x85055, x85056, x85057, x85058, x85059, x85060;
  wire x85061, x85062, x85063, x85064, x85065, x85066, x85067, x85068;
  wire x85069, x85070, x85071, x85072, x85073, x85074, x85075, x85076;
  wire x85077, x85078, x85079, x85080, x85081, x85082, x85083, x85084;
  wire x85085, x85086, x85087, x85088, x85089, x85090, x85091, x85092;
  wire x85093, x85094, x85095, x85096, x85097, x85098, x85099, x85100;
  wire x85101, x85102, x85103, x85104, x85105, x85106, x85107, x85108;
  wire x85109, x85110, x85111, x85112, x85113, x85114, x85115, x85116;
  wire x85117, x85118, x85119, x85120, x85121, x85122, x85123, x85124;
  wire x85125, x85126, x85127, x85128, x85129, x85130, x85131, x85132;
  wire x85133, x85134, x85135, x85136, x85137, x85138, x85139, x85140;
  wire x85141, x85142, x85143, x85144, x85145, x85146, x85147, x85148;
  wire x85149, x85150, x85151, x85152, x85153, x85154, x85155, x85156;
  wire x85157, x85158, x85159, x85160, x85161, x85162, x85163, x85164;
  wire x85165, x85166, x85167, x85168, x85169, x85170, x85171, x85172;
  wire x85173, x85174, x85175, x85176, x85177, x85178, x85179, x85180;
  wire x85181, x85182, x85183, x85184, x85185, x85186, x85187, x85188;
  wire x85189, x85190, x85191, x85192, x85193, x85194, x85195, x85196;
  wire x85197, x85198, x85199, x85200, x85201, x85202, x85203, x85204;
  wire x85205, x85206, x85207, x85208, x85209, x85210, x85211, x85212;
  wire x85213, x85214, x85215, x85216, x85217, x85218, x85219, x85220;
  wire x85221, x85222, x85223, x85224, x85225, x85226, x85227, x85228;
  wire x85229, x85230, x85231, x85232, x85233, x85234, x85235, x85236;
  wire x85237, x85238, x85239, x85240, x85241, x85242, x85243, x85244;
  wire x85245, x85246, x85247, x85248, x85249, x85250, x85251, x85252;
  wire x85253, x85254, x85255, x85256, x85257, x85258, x85259, x85260;
  wire x85261, x85262, x85263, x85264, x85265, x85266, x85267, x85268;
  wire x85269, x85270, x85271, x85272, x85273, x85274, x85275, x85276;
  wire x85277, x85278, x85279, x85280, x85281, x85282, x85283, x85284;
  wire x85285, x85286, x85287, x85288, x85289, x85290, x85291, x85292;
  wire x85293, x85294, x85295, x85296, x85297, x85298, x85299, x85300;
  wire x85301, x85302, x85303, x85304, x85305, x85306, x85307, x85308;
  wire x85309, x85310, x85311, x85312, x85313, x85314, x85315, x85316;
  wire x85317, x85318, x85319, x85320, x85321, x85322, x85323, x85324;
  wire x85325, x85326, x85327, x85328, x85329, x85330, x85331, x85332;
  wire x85333, x85334, x85335, x85336, x85337, x85338, x85339, x85340;
  wire x85341, x85342, x85343, x85344, x85345, x85346, x85347, x85348;
  wire x85349, x85350, x85351, x85352, x85353, x85354, x85355, x85356;
  wire x85357, x85358, x85359, x85360, x85361, x85362, x85363, x85364;
  wire x85365, x85366, x85367, x85368, x85369, x85370, x85371, x85372;
  wire x85373, x85374, x85375, x85376, x85377, x85378, x85379, x85380;
  wire x85381, x85382, x85383, x85384, x85385, x85386, x85387, x85388;
  wire x85389, x85390, x85391, x85392, x85393, x85394, x85395, x85396;
  wire x85397, x85398, x85399, x85400, x85401, x85402, x85403, x85404;
  wire x85405, x85406, x85407, x85408, x85409, x85410, x85411, x85412;
  wire x85413, x85414, x85415, x85416, x85417, x85418, x85419, x85420;
  wire x85421, x85422, x85423, x85424, x85425, x85426, x85427, x85428;
  wire x85429, x85430, x85431, x85432, x85433, x85434, x85435, x85436;
  wire x85437, x85438, x85439, x85440, x85441, x85442, x85443, x85444;
  wire x85445, x85446, x85447, x85448, x85449, x85450, x85451, x85452;
  wire x85453, x85454, x85455, x85456, x85457, x85458, x85459, x85460;
  wire x85461, x85462, x85463, x85464, x85465, x85466, x85467, x85468;
  wire x85469, x85470, x85471, x85472, x85473, x85474, x85475, x85476;
  wire x85477, x85478, x85479, x85480, x85481, x85482, x85483, x85484;
  wire x85485, x85486, x85487, x85488, x85489, x85490, x85491, x85492;
  wire x85493, x85494, x85495, x85496, x85497, x85498, x85499, x85500;
  wire x85501, x85502, x85503, x85504, x85505, x85506, x85507, x85508;
  wire x85509, x85510, x85511, x85512, x85513, x85514, x85515, x85516;
  wire x85517, x85518, x85519, x85520, x85521, x85522, x85523, x85524;
  wire x85525, x85526, x85527, x85528, x85529, x85530, x85531, x85532;
  wire x85533, x85534, x85535, x85536, x85537, x85538, x85539, x85540;
  wire x85541, x85542, x85543, x85544, x85545, x85546, x85547, x85548;
  wire x85549, x85550, x85551, x85552, x85553, x85554, x85555, x85556;
  wire x85557, x85558, x85559, x85560, x85561, x85562, x85563, x85564;
  wire x85565, x85566, x85567, x85568, x85569, x85570, x85571, x85572;
  wire x85573, x85574, x85575, x85576, x85577, x85578, x85579, x85580;
  wire x85581, x85582, x85583, x85584, x85585, x85586, x85587, x85588;
  wire x85589, x85590, x85591, x85592, x85593, x85594, x85595, x85596;
  wire x85597, x85598, x85599, x85600, x85601, x85602, x85603, x85604;
  wire x85605, x85606, x85607, x85608, x85609, x85610, x85611, x85612;
  wire x85613, x85614, x85615, x85616, x85617, x85618, x85619, x85620;
  wire x85621, x85622, x85623, x85624, x85625, x85626, x85627, x85628;
  wire x85629, x85630, x85631, x85632, x85633, x85634, x85635, x85636;
  wire x85637, x85638, x85639, x85640, x85641, x85642, x85643, x85644;
  wire x85645, x85646, x85647, x85648, x85649, x85650, x85651, x85652;
  wire x85653, x85654, x85655, x85656, x85657, x85658, x85659, x85660;
  wire x85661, x85662, x85663, x85664, x85665, x85666, x85667, x85668;
  wire x85669, x85670, x85671, x85672, x85673, x85674, x85675, x85676;
  wire x85677, x85678, x85679, x85680, x85681, x85682, x85683, x85684;
  wire x85685, x85686, x85687, x85688, x85689, x85690, x85691, x85692;
  wire x85693, x85694, x85695, x85696, x85697, x85698, x85699, x85700;
  wire x85701, x85702, x85703, x85704, x85705, x85706, x85707, x85708;
  wire x85709, x85710, x85711, x85712, x85713, x85714, x85715, x85716;
  wire x85717, x85718, x85719, x85720, x85721, x85722, x85723, x85724;
  wire x85725, x85726, x85727, x85728, x85729, x85730, x85731, x85732;
  wire x85733, x85734, x85735, x85736, x85737, x85738, x85739, x85740;
  wire x85741, x85742, x85743, x85744, x85745, x85746, x85747, x85748;
  wire x85749, x85750, x85751, x85752, x85753, x85754, x85755, x85756;
  wire x85757, x85758, x85759, x85760, x85761, x85762, x85763, x85764;
  wire x85765, x85766, x85767, x85768, x85769, x85770, x85771, x85772;
  wire x85773, x85774, x85775, x85776, x85777, x85778, x85779, x85780;
  wire x85781, x85782, x85783, x85784, x85785, x85786, x85787, x85788;
  wire x85789, x85790, x85791, x85792, x85793, x85794, x85795, x85796;
  wire x85797, x85798, x85799, x85800, x85801, x85802, x85803, x85804;
  wire x85805, x85806, x85807, x85808, x85809, x85810, x85811, x85812;
  wire x85813, x85814, x85815, x85816, x85817, x85818, x85819, x85820;
  wire x85821, x85822, x85823, x85824, x85825, x85826, x85827, x85828;
  wire x85829, x85830, x85831, x85832, x85833, x85834, x85835, x85836;
  wire x85837, x85838, x85839, x85840, x85841, x85842, x85843, x85844;
  wire x85845, x85846, x85847, x85848, x85849, x85850, x85851, x85852;
  wire x85853, x85854, x85855, x85856, x85857, x85858, x85859, x85860;
  wire x85861, x85862, x85863, x85864, x85865, x85866, x85867, x85868;
  wire x85869, x85870, x85871, x85872, x85873, x85874, x85875, x85876;
  wire x85877, x85878, x85879, x85880, x85881, x85882, x85883, x85884;
  wire x85885, x85886, x85887, x85888, x85889, x85890, x85891, x85892;
  wire x85893, x85894, x85895, x85896, x85897, x85898, x85899, x85900;
  wire x85901, x85902, x85903, x85904, x85905, x85906, x85907, x85908;
  wire x85909, x85910, x85911, x85912, x85913, x85914, x85915, x85916;
  wire x85917, x85918, x85919, x85920, x85921, x85922, x85923, x85924;
  wire x85925, x85926, x85927, x85928, x85929, x85930, x85931, x85932;
  wire x85933, x85934, x85935, x85936, x85937, x85938, x85939, x85940;
  wire x85941, x85942, x85943, x85944, x85945, x85946, x85947, x85948;
  wire x85949, x85950, x85951, x85952, x85953, x85954, x85955, x85956;
  wire x85957, x85958, x85959, x85960, x85961, x85962, x85963, x85964;
  wire x85965, x85966, x85967, x85968, x85969, x85970, x85971, x85972;
  wire x85973, x85974, x85975, x85976, x85977, x85978, x85979, x85980;
  wire x85981, x85982, x85983, x85984, x85985, x85986, x85987, x85988;
  wire x85989, x85990, x85991, x85992, x85993, x85994, x85995, x85996;
  wire x85997, x85998, x85999, x86000, x86001, x86002, x86003, x86004;
  wire x86005, x86006, x86007, x86008, x86009, x86010, x86011, x86012;
  wire x86013, x86014, x86015, x86016, x86017, x86018, x86019, x86020;
  wire x86021, x86022, x86023, x86024, x86025, x86026, x86027, x86028;
  wire x86029, x86030, x86031, x86032, x86033, x86034, x86035, x86036;
  wire x86037, x86038, x86039, x86040, x86041, x86042, x86043, x86044;
  wire x86045, x86046, x86047, x86048, x86049, x86050, x86051, x86052;
  wire x86053, x86054, x86055, x86056, x86057, x86058, x86059, x86060;
  wire x86061, x86062, x86063, x86064, x86065, x86066, x86067, x86068;
  wire x86069, x86070, x86071, x86072, x86073, x86074, x86075, x86076;
  wire x86077, x86078, x86079, x86080, x86081, x86082, x86083, x86084;
  wire x86085, x86086, x86087, x86088, x86089, x86090, x86091, x86092;
  wire x86093, x86094, x86095, x86096, x86097, x86098, x86099, x86100;
  wire x86101, x86102, x86103, x86104, x86105, x86106, x86107, x86108;
  wire x86109, x86110, x86111, x86112, x86113, x86114, x86115, x86116;
  wire x86117, x86118, x86119, x86120, x86121, x86122, x86123, x86124;
  wire x86125, x86126, x86127, x86128, x86129, x86130, x86131, x86132;
  wire x86133, x86134, x86135, x86136, x86137, x86138, x86139, x86140;
  wire x86141, x86142, x86143, x86144, x86145, x86146, x86147, x86148;
  wire x86149, x86150, x86151, x86152, x86153, x86154, x86155, x86156;
  wire x86157, x86158, x86159, x86160, x86161, x86162, x86163, x86164;
  wire x86165, x86166, x86167, x86168, x86169, x86170, x86171, x86172;
  wire x86173, x86174, x86175, x86176, x86177, x86178, x86179, x86180;
  wire x86181, x86182, x86183, x86184, x86185, x86186, x86187, x86188;
  wire x86189, x86190, x86191, x86192, x86193, x86194, x86195, x86196;
  wire x86197, x86198, x86199, x86200, x86201, x86202, x86203, x86204;
  wire x86205, x86206, x86207, x86208, x86209, x86210, x86211, x86212;
  wire x86213, x86214, x86215, x86216, x86217, x86218, x86219, x86220;
  wire x86221, x86222, x86223, x86224, x86225, x86226, x86227, x86228;
  wire x86229, x86230, x86231, x86232, x86233, x86234, x86235, x86236;
  wire x86237, x86238, x86239, x86240, x86241, x86242, x86243, x86244;
  wire x86245, x86246, x86247, x86248, x86249, x86250, x86251, x86252;
  wire x86253, x86254, x86255, x86256, x86257, x86258, x86259, x86260;
  wire x86261, x86262, x86263, x86264, x86265, x86266, x86267, x86268;
  wire x86269, x86270, x86271, x86272, x86273, x86274, x86275, x86276;
  wire x86277, x86278, x86279, x86280, x86281, x86282, x86283, x86284;
  wire x86285, x86286, x86287, x86288, x86289, x86290, x86291, x86292;
  wire x86293, x86294, x86295, x86296, x86297, x86298, x86299, x86300;
  wire x86301, x86302, x86303, x86304, x86305, x86306, x86307, x86308;
  wire x86309, x86310, x86311, x86312, x86313, x86314, x86315, x86316;
  wire x86317, x86318, x86319, x86320, x86321, x86322, x86323, x86324;
  wire x86325, x86326, x86327, x86328, x86329, x86330, x86331, x86332;
  wire x86333, x86334, x86335, x86336, x86337, x86338, x86339, x86340;
  wire x86341, x86342, x86343, x86344, x86345, x86346, x86347, x86348;
  wire x86349, x86350, x86351, x86352, x86353, x86354, x86355, x86356;
  wire x86357, x86358, x86359, x86360, x86361, x86362, x86363, x86364;
  wire x86365, x86366, x86367, x86368, x86369, x86370, x86371, x86372;
  wire x86373, x86374, x86375, x86376, x86377, x86378, x86379, x86380;
  wire x86381, x86382, x86383, x86384, x86385, x86386, x86387, x86388;
  wire x86389, x86390, x86391, x86392, x86393, x86394, x86395, x86396;
  wire x86397, x86398, x86399, x86400, x86401, x86402, x86403, x86404;
  wire x86405, x86406, x86407, x86408, x86409, x86410, x86411, x86412;
  wire x86413, x86414, x86415, x86416, x86417, x86418, x86419, x86420;
  wire x86421, x86422, x86423, x86424, x86425, x86426, x86427, x86428;
  wire x86429, x86430, x86431, x86432, x86433, x86434, x86435, x86436;
  wire x86437, x86438, x86439, x86440, x86441, x86442, x86443, x86444;
  wire x86445, x86446, x86447, x86448, x86449, x86450, x86451, x86452;
  wire x86453, x86454, x86455, x86456, x86457, x86458, x86459, x86460;
  wire x86461, x86462, x86463, x86464, x86465, x86466, x86467, x86468;
  wire x86469, x86470, x86471, x86472, x86473, x86474, x86475, x86476;
  wire x86477, x86478, x86479, x86480, x86481, x86482, x86483, x86484;
  wire x86485, x86486, x86487, x86488, x86489, x86490, x86491, x86492;
  wire x86493, x86494, x86495, x86496, x86497, x86498, x86499, x86500;
  wire x86501, x86502, x86503, x86504, x86505, x86506, x86507, x86508;
  wire x86509, x86510, x86511, x86512, x86513, x86514, x86515, x86516;
  wire x86517, x86518, x86519, x86520, x86521, x86522, x86523, x86524;
  wire x86525, x86526, x86527, x86528, x86529, x86530, x86531, x86532;
  wire x86533, x86534, x86535, x86536, x86537, x86538, x86539, x86540;
  wire x86541, x86542, x86543, x86544, x86545, x86546, x86547, x86548;
  wire x86549, x86550, x86551, x86552, x86553, x86554, x86555, x86556;
  wire x86557, x86558, x86559, x86560, x86561, x86562, x86563, x86564;
  wire x86565, x86566, x86567, x86568, x86569, x86570, x86571, x86572;
  wire x86573, x86574, x86575, x86576, x86577, x86578, x86579, x86580;
  wire x86581, x86582, x86583, x86584, x86585, x86586, x86587, x86588;
  wire x86589, x86590, x86591, x86592, x86593, x86594, x86595, x86596;
  wire x86597, x86598, x86599, x86600, x86601, x86602, x86603, x86604;
  wire x86605, x86606, x86607, x86608, x86609, x86610, x86611, x86612;
  wire x86613, x86614, x86615, x86616, x86617, x86618, x86619, x86620;
  wire x86621, x86622, x86623, x86624, x86625, x86626, x86627, x86628;
  wire x86629, x86630, x86631, x86632, x86633, x86634, x86635, x86636;
  wire x86637, x86638, x86639, x86640, x86641, x86642, x86643, x86644;
  wire x86645, x86646, x86647, x86648, x86649, x86650, x86651, x86652;
  wire x86653, x86654, x86655, x86656, x86657, x86658, x86659, x86660;
  wire x86661, x86662, x86663, x86664, x86665, x86666, x86667, x86668;
  wire x86669, x86670, x86671, x86672, x86673, x86674, x86675, x86676;
  wire x86677, x86678, x86679, x86680, x86681, x86682, x86683, x86684;
  wire x86685, x86686, x86687, x86688, x86689, x86690, x86691, x86692;
  wire x86693, x86694, x86695, x86696, x86697, x86698, x86699, x86700;
  wire x86701, x86702, x86703, x86704, x86705, x86706, x86707, x86708;
  wire x86709, x86710, x86711, x86712, x86713, x86714, x86715, x86716;
  wire x86717, x86718, x86719, x86720, x86721, x86722, x86723, x86724;
  wire x86725, x86726, x86727, x86728, x86729, x86730, x86731, x86732;
  wire x86733, x86734, x86735, x86736, x86737, x86738, x86739, x86740;
  wire x86741, x86742, x86743, x86744, x86745, x86746, x86747, x86748;
  wire x86749, x86750, x86751, x86752, x86753, x86754, x86755, x86756;
  wire x86757, x86758, x86759, x86760, x86761, x86762, x86763, x86764;
  wire x86765, x86766, x86767, x86768, x86769, x86770, x86771, x86772;
  wire x86773, x86774, x86775, x86776, x86777, x86778, x86779, x86780;
  wire x86781, x86782, x86783, x86784, x86785, x86786, x86787, x86788;
  wire x86789, x86790, x86791, x86792, x86793, x86794, x86795, x86796;
  wire x86797, x86798, x86799, x86800, x86801, x86802, x86803, x86804;
  wire x86805, x86806, x86807, x86808, x86809, x86810, x86811, x86812;
  wire x86813, x86814, x86815, x86816, x86817, x86818, x86819, x86820;
  wire x86821, x86822, x86823, x86824, x86825, x86826, x86827, x86828;
  wire x86829, x86830, x86831, x86832, x86833, x86834, x86835, x86836;
  wire x86837, x86838, x86839, x86840, x86841, x86842, x86843, x86844;
  wire x86845, x86846, x86847, x86848, x86849, x86850, x86851, x86852;
  wire x86853, x86854, x86855, x86856, x86857, x86858, x86859, x86860;
  wire x86861, x86862, x86863, x86864, x86865, x86866, x86867, x86868;
  wire x86869, x86870, x86871, x86872, x86873, x86874, x86875, x86876;
  wire x86877, x86878, x86879, x86880, x86881, x86882, x86883, x86884;
  wire x86885, x86886, x86887, x86888, x86889, x86890, x86891, x86892;
  wire x86893, x86894, x86895, x86896, x86897, x86898, x86899, x86900;
  wire x86901, x86902, x86903, x86904, x86905, x86906, x86907, x86908;
  wire x86909, x86910, x86911, x86912, x86913, x86914, x86915, x86916;
  wire x86917, x86918, x86919, x86920, x86921, x86922, x86923, x86924;
  wire x86925, x86926, x86927, x86928, x86929, x86930, x86931, x86932;
  wire x86933, x86934, x86935, x86936, x86937, x86938, x86939, x86940;
  wire x86941, x86942, x86943, x86944, x86945, x86946, x86947, x86948;
  wire x86949, x86950, x86951, x86952, x86953, x86954, x86955, x86956;
  wire x86957, x86958, x86959, x86960, x86961, x86962, x86963, x86964;
  wire x86965, x86966, x86967, x86968, x86969, x86970, x86971, x86972;
  wire x86973, x86974, x86975, x86976, x86977, x86978, x86979, x86980;
  wire x86981, x86982, x86983, x86984, x86985, x86986, x86987, x86988;
  wire x86989, x86990, x86991, x86992, x86993, x86994, x86995, x86996;
  wire x86997, x86998, x86999, x87000, x87001, x87002, x87003, x87004;
  wire x87005, x87006, x87007, x87008, x87009, x87010, x87011, x87012;
  wire x87013, x87014, x87015, x87016, x87017, x87018, x87019, x87020;
  wire x87021, x87022, x87023, x87024, x87025, x87026, x87027, x87028;
  wire x87029, x87030, x87031, x87032, x87033, x87034, x87035, x87036;
  wire x87037, x87038, x87039, x87040, x87041, x87042, x87043, x87044;
  wire x87045, x87046, x87047, x87048, x87049, x87050, x87051, x87052;
  wire x87053, x87054, x87055, x87056, x87057, x87058, x87059, x87060;
  wire x87061, x87062, x87063, x87064, x87065, x87066, x87067, x87068;
  wire x87069, x87070, x87071, x87072, x87073, x87074, x87075, x87076;
  wire x87077, x87078, x87079, x87080, x87081, x87082, x87083, x87084;
  wire x87085, x87086, x87087, x87088, x87089, x87090, x87091, x87092;
  wire x87093, x87094, x87095, x87096, x87097, x87098, x87099, x87100;
  wire x87101, x87102, x87103, x87104, x87105, x87106, x87107, x87108;
  wire x87109, x87110, x87111, x87112, x87113, x87114, x87115, x87116;
  wire x87117, x87118, x87119, x87120, x87121, x87122, x87123, x87124;
  wire x87125, x87126, x87127, x87128, x87129, x87130, x87131, x87132;
  wire x87133, x87134, x87135, x87136, x87137, x87138, x87139, x87140;
  wire x87141, x87142, x87143, x87144, x87145, x87146, x87147, x87148;
  wire x87149, x87150, x87151, x87152, x87153, x87154, x87155, x87156;
  wire x87157, x87158, x87159, x87160, x87161, x87162, x87163, x87164;
  wire x87165, x87166, x87167, x87168, x87169, x87170, x87171, x87172;
  wire x87173, x87174, x87175, x87176, x87177, x87178, x87179, x87180;
  wire x87181, x87182, x87183, x87184, x87185, x87186, x87187, x87188;
  wire x87189, x87190, x87191, x87192, x87193, x87194, x87195, x87196;
  wire x87197, x87198, x87199, x87200, x87201, x87202, x87203, x87204;
  wire x87205, x87206, x87207, x87208, x87209, x87210, x87211, x87212;
  wire x87213, x87214, x87215, x87216, x87217, x87218, x87219, x87220;
  wire x87221, x87222, x87223, x87224, x87225, x87226, x87227, x87228;
  wire x87229, x87230, x87231, x87232, x87233, x87234, x87235, x87236;
  wire x87237, x87238, x87239, x87240, x87241, x87242, x87243, x87244;
  wire x87245, x87246, x87247, x87248, x87249, x87250, x87251, x87252;
  wire x87253, x87254, x87255, x87256, x87257, x87258, x87259, x87260;
  wire x87261, x87262, x87263, x87264;

  nand n2(x2, x1, x0);
  nand n9(x9, x59, x58);
  nand n10(x10, x60, x59);
  nand n12(x12, x61, x60);
  nand n14(x14, x62, x61);
  nand n16(x16, x11, x58);
  nand n17(x17, x13, x83383);
  nand n18(x18, x15, x11);
  nand n20(x20, x19, x58);
  nand n21(x21, x3, x8);
  nand n22(x22, x21, x9);
  nand n24(x24, x60, x83383);
  nand n25(x25, x4, x9);
  nand n26(x26, x25, x24);
  nand n28(x28, x61, x83384);
  nand n29(x29, x5, x16);
  nand n30(x30, x29, x28);
  nand n32(x32, x62, x83385);
  nand n33(x33, x6, x17);
  nand n34(x34, x33, x32);
  nand n36(x36, x63, x83386);
  nand n37(x37, x7, x20);
  nand n38(x38, x37, x36);
  nand n40(x40, x71140, x58);
  nand n41(x41, x1, x8);
  nand n42(x42, x41, x40);
  nand n43(x43, x71140, x59);
  nand n44(x44, x1, x23);
  nand n45(x45, x44, x43);
  nand n46(x46, x71140, x60);
  nand n47(x47, x1, x27);
  nand n48(x48, x47, x46);
  nand n49(x49, x71140, x61);
  nand n50(x50, x1, x31);
  nand n51(x51, x50, x49);
  nand n52(x52, x71140, x62);
  nand n53(x53, x1, x35);
  nand n54(x54, x53, x52);
  nand n55(x55, x71140, x63);
  nand n56(x56, x1, x39);
  nand n57(x57, x56, x55);
  nand n94(x94, x605, x604);
  nand n95(x95, x606, x605);
  nand n97(x97, x607, x606);
  nand n99(x99, x608, x607);
  nand n101(x101, x609, x608);
  nand n103(x103, x610, x609);
  nand n105(x105, x611, x610);
  nand n107(x107, x612, x611);
  nand n109(x109, x613, x612);
  nand n111(x111, x614, x613);
  nand n113(x113, x615, x614);
  nand n115(x115, x616, x615);
  nand n117(x117, x617, x616);
  nand n119(x119, x618, x617);
  nand n121(x121, x619, x618);
  nand n123(x123, x620, x619);
  nand n125(x125, x621, x620);
  nand n127(x127, x622, x621);
  nand n129(x129, x623, x622);
  nand n131(x131, x624, x623);
  nand n133(x133, x625, x624);
  nand n135(x135, x626, x625);
  nand n137(x137, x627, x626);
  nand n139(x139, x628, x627);
  nand n141(x141, x629, x628);
  nand n143(x143, x630, x629);
  nand n145(x145, x631, x630);
  nand n147(x147, x632, x631);
  nand n149(x149, x96, x604);
  nand n150(x150, x98, x83387);
  nand n151(x151, x100, x96);
  nand n153(x153, x102, x98);
  nand n155(x155, x104, x100);
  nand n157(x157, x106, x102);
  nand n159(x159, x108, x104);
  nand n161(x161, x110, x106);
  nand n163(x163, x112, x108);
  nand n165(x165, x114, x110);
  nand n167(x167, x116, x112);
  nand n169(x169, x118, x114);
  nand n171(x171, x120, x116);
  nand n173(x173, x122, x118);
  nand n175(x175, x124, x120);
  nand n177(x177, x126, x122);
  nand n179(x179, x128, x124);
  nand n181(x181, x130, x126);
  nand n183(x183, x132, x128);
  nand n185(x185, x134, x130);
  nand n187(x187, x136, x132);
  nand n189(x189, x138, x134);
  nand n191(x191, x140, x136);
  nand n193(x193, x142, x138);
  nand n195(x195, x144, x140);
  nand n197(x197, x146, x142);
  nand n199(x199, x148, x144);
  nand n201(x201, x152, x604);
  nand n202(x202, x154, x83387);
  nand n203(x203, x156, x83388);
  nand n204(x204, x158, x83389);
  nand n205(x205, x160, x152);
  nand n207(x207, x162, x154);
  nand n209(x209, x164, x156);
  nand n211(x211, x166, x158);
  nand n213(x213, x168, x160);
  nand n215(x215, x170, x162);
  nand n217(x217, x172, x164);
  nand n219(x219, x174, x166);
  nand n221(x221, x176, x168);
  nand n223(x223, x178, x170);
  nand n225(x225, x180, x172);
  nand n227(x227, x182, x174);
  nand n229(x229, x184, x176);
  nand n231(x231, x186, x178);
  nand n233(x233, x188, x180);
  nand n235(x235, x190, x182);
  nand n237(x237, x192, x184);
  nand n239(x239, x194, x186);
  nand n241(x241, x196, x188);
  nand n243(x243, x198, x190);
  nand n245(x245, x200, x192);
  nand n247(x247, x206, x604);
  nand n248(x248, x208, x83387);
  nand n249(x249, x210, x83388);
  nand n250(x250, x212, x83389);
  nand n251(x251, x214, x83390);
  nand n252(x252, x216, x83391);
  nand n253(x253, x218, x83392);
  nand n254(x254, x220, x83393);
  nand n255(x255, x222, x206);
  nand n257(x257, x224, x208);
  nand n259(x259, x226, x210);
  nand n261(x261, x228, x212);
  nand n263(x263, x230, x214);
  nand n265(x265, x232, x216);
  nand n267(x267, x234, x218);
  nand n269(x269, x236, x220);
  nand n271(x271, x238, x222);
  nand n273(x273, x240, x224);
  nand n275(x275, x242, x226);
  nand n277(x277, x244, x228);
  nand n279(x279, x246, x230);
  nand n281(x281, x256, x604);
  nand n282(x282, x258, x83387);
  nand n283(x283, x260, x83388);
  nand n284(x284, x262, x83389);
  nand n285(x285, x264, x83390);
  nand n286(x286, x266, x83391);
  nand n287(x287, x268, x83392);
  nand n288(x288, x270, x83393);
  nand n289(x289, x272, x83394);
  nand n290(x290, x274, x83395);
  nand n291(x291, x276, x83396);
  nand n292(x292, x278, x83397);
  nand n293(x293, x280, x83398);
  nand n294(x294, x64, x93);
  nand n295(x295, x294, x94);
  nand n297(x297, x606, x83387);
  nand n298(x298, x65, x94);
  nand n299(x299, x298, x297);
  nand n301(x301, x607, x83388);
  nand n302(x302, x66, x149);
  nand n303(x303, x302, x301);
  nand n305(x305, x608, x83389);
  nand n306(x306, x67, x150);
  nand n307(x307, x306, x305);
  nand n309(x309, x609, x83390);
  nand n310(x310, x68, x201);
  nand n311(x311, x310, x309);
  nand n313(x313, x610, x83391);
  nand n314(x314, x69, x202);
  nand n315(x315, x314, x313);
  nand n317(x317, x611, x83392);
  nand n318(x318, x70, x203);
  nand n319(x319, x318, x317);
  nand n321(x321, x612, x83393);
  nand n322(x322, x71, x204);
  nand n323(x323, x322, x321);
  nand n325(x325, x613, x83394);
  nand n326(x326, x72, x247);
  nand n327(x327, x326, x325);
  nand n329(x329, x614, x83395);
  nand n330(x330, x73, x248);
  nand n331(x331, x330, x329);
  nand n333(x333, x615, x83396);
  nand n334(x334, x74, x249);
  nand n335(x335, x334, x333);
  nand n337(x337, x616, x83397);
  nand n338(x338, x75, x250);
  nand n339(x339, x338, x337);
  nand n341(x341, x617, x83398);
  nand n342(x342, x76, x251);
  nand n343(x343, x342, x341);
  nand n345(x345, x618, x83399);
  nand n346(x346, x77, x252);
  nand n347(x347, x346, x345);
  nand n349(x349, x619, x83400);
  nand n350(x350, x78, x253);
  nand n351(x351, x350, x349);
  nand n353(x353, x620, x83401);
  nand n354(x354, x79, x254);
  nand n355(x355, x354, x353);
  nand n357(x357, x621, x83402);
  nand n358(x358, x80, x281);
  nand n359(x359, x358, x357);
  nand n361(x361, x622, x83403);
  nand n362(x362, x81, x282);
  nand n363(x363, x362, x361);
  nand n365(x365, x623, x83404);
  nand n366(x366, x82, x283);
  nand n367(x367, x366, x365);
  nand n369(x369, x624, x83405);
  nand n370(x370, x83, x284);
  nand n371(x371, x370, x369);
  nand n373(x373, x625, x83406);
  nand n374(x374, x84, x285);
  nand n375(x375, x374, x373);
  nand n377(x377, x626, x83407);
  nand n378(x378, x85, x286);
  nand n379(x379, x378, x377);
  nand n381(x381, x627, x83408);
  nand n382(x382, x86, x287);
  nand n383(x383, x382, x381);
  nand n385(x385, x628, x83409);
  nand n386(x386, x87, x288);
  nand n387(x387, x386, x385);
  nand n389(x389, x629, x83410);
  nand n390(x390, x88, x289);
  nand n391(x391, x390, x389);
  nand n393(x393, x630, x83411);
  nand n394(x394, x89, x290);
  nand n395(x395, x394, x393);
  nand n397(x397, x631, x83412);
  nand n398(x398, x90, x291);
  nand n399(x399, x398, x397);
  nand n401(x401, x632, x83413);
  nand n402(x402, x91, x292);
  nand n403(x403, x402, x401);
  nand n405(x405, x633, x83414);
  nand n406(x406, x92, x293);
  nand n407(x407, x406, x405);
  nand n409(x409, x2, x602);
  nand n411(x411, x410, x602);
  nand n412(x412, x411, x409);
  nand n413(x413, x2, x603);
  nand n414(x414, x410, x603);
  nand n415(x415, x414, x413);
  nand n416(x416, x2, x604);
  nand n417(x417, x410, x93);
  nand n418(x418, x417, x416);
  nand n419(x419, x2, x605);
  nand n420(x420, x410, x296);
  nand n421(x421, x420, x419);
  nand n422(x422, x2, x606);
  nand n423(x423, x410, x300);
  nand n424(x424, x423, x422);
  nand n425(x425, x2, x607);
  nand n426(x426, x410, x304);
  nand n427(x427, x426, x425);
  nand n428(x428, x2, x608);
  nand n429(x429, x410, x308);
  nand n430(x430, x429, x428);
  nand n431(x431, x2, x609);
  nand n432(x432, x410, x312);
  nand n433(x433, x432, x431);
  nand n434(x434, x2, x610);
  nand n435(x435, x410, x316);
  nand n436(x436, x435, x434);
  nand n437(x437, x2, x611);
  nand n438(x438, x410, x320);
  nand n439(x439, x438, x437);
  nand n440(x440, x2, x612);
  nand n441(x441, x410, x324);
  nand n442(x442, x441, x440);
  nand n443(x443, x2, x613);
  nand n444(x444, x410, x328);
  nand n445(x445, x444, x443);
  nand n446(x446, x2, x614);
  nand n447(x447, x410, x332);
  nand n448(x448, x447, x446);
  nand n449(x449, x2, x615);
  nand n450(x450, x410, x336);
  nand n451(x451, x450, x449);
  nand n452(x452, x2, x616);
  nand n453(x453, x410, x340);
  nand n454(x454, x453, x452);
  nand n455(x455, x2, x617);
  nand n456(x456, x410, x344);
  nand n457(x457, x456, x455);
  nand n458(x458, x2, x618);
  nand n459(x459, x410, x348);
  nand n460(x460, x459, x458);
  nand n461(x461, x2, x619);
  nand n462(x462, x410, x352);
  nand n463(x463, x462, x461);
  nand n464(x464, x2, x620);
  nand n465(x465, x410, x356);
  nand n466(x466, x465, x464);
  nand n467(x467, x2, x621);
  nand n468(x468, x410, x360);
  nand n469(x469, x468, x467);
  nand n470(x470, x2, x622);
  nand n471(x471, x410, x364);
  nand n472(x472, x471, x470);
  nand n473(x473, x2, x623);
  nand n474(x474, x410, x368);
  nand n475(x475, x474, x473);
  nand n476(x476, x2, x624);
  nand n477(x477, x410, x372);
  nand n478(x478, x477, x476);
  nand n479(x479, x2, x625);
  nand n480(x480, x410, x376);
  nand n481(x481, x480, x479);
  nand n482(x482, x2, x626);
  nand n483(x483, x410, x380);
  nand n484(x484, x483, x482);
  nand n485(x485, x2, x627);
  nand n486(x486, x410, x384);
  nand n487(x487, x486, x485);
  nand n488(x488, x2, x628);
  nand n489(x489, x410, x388);
  nand n490(x490, x489, x488);
  nand n491(x491, x2, x629);
  nand n492(x492, x410, x392);
  nand n493(x493, x492, x491);
  nand n494(x494, x2, x630);
  nand n495(x495, x410, x396);
  nand n496(x496, x495, x494);
  nand n497(x497, x2, x631);
  nand n498(x498, x410, x400);
  nand n499(x499, x498, x497);
  nand n500(x500, x2, x632);
  nand n501(x501, x410, x404);
  nand n502(x502, x501, x500);
  nand n503(x503, x2, x633);
  nand n504(x504, x410, x408);
  nand n505(x505, x504, x503);
  nand n506(x506, x15229, x16412);
  nand n507(x507, x15228, x412);
  nand n508(x508, x507, x506);
  nand n509(x509, x15229, x16415);
  nand n510(x510, x15228, x415);
  nand n511(x511, x510, x509);
  nand n512(x512, x15229, x16418);
  nand n513(x513, x15228, x418);
  nand n514(x514, x513, x512);
  nand n515(x515, x15229, x16421);
  nand n516(x516, x15228, x421);
  nand n517(x517, x516, x515);
  nand n518(x518, x15229, x16424);
  nand n519(x519, x15228, x424);
  nand n520(x520, x519, x518);
  nand n521(x521, x15229, x16427);
  nand n522(x522, x15228, x427);
  nand n523(x523, x522, x521);
  nand n524(x524, x15229, x16430);
  nand n525(x525, x15228, x430);
  nand n526(x526, x525, x524);
  nand n527(x527, x15229, x16433);
  nand n528(x528, x15228, x433);
  nand n529(x529, x528, x527);
  nand n530(x530, x15229, x16436);
  nand n531(x531, x15228, x436);
  nand n532(x532, x531, x530);
  nand n533(x533, x15229, x16439);
  nand n534(x534, x15228, x439);
  nand n535(x535, x534, x533);
  nand n536(x536, x15229, x16442);
  nand n537(x537, x15228, x442);
  nand n538(x538, x537, x536);
  nand n539(x539, x15229, x16445);
  nand n540(x540, x15228, x445);
  nand n541(x541, x540, x539);
  nand n542(x542, x15229, x16448);
  nand n543(x543, x15228, x448);
  nand n544(x544, x543, x542);
  nand n545(x545, x15229, x16451);
  nand n546(x546, x15228, x451);
  nand n547(x547, x546, x545);
  nand n548(x548, x15229, x16454);
  nand n549(x549, x15228, x454);
  nand n550(x550, x549, x548);
  nand n551(x551, x15229, x16457);
  nand n552(x552, x15228, x457);
  nand n553(x553, x552, x551);
  nand n554(x554, x15229, x16460);
  nand n555(x555, x15228, x460);
  nand n556(x556, x555, x554);
  nand n557(x557, x15229, x16463);
  nand n558(x558, x15228, x463);
  nand n559(x559, x558, x557);
  nand n560(x560, x15229, x16466);
  nand n561(x561, x15228, x466);
  nand n562(x562, x561, x560);
  nand n563(x563, x15229, x16469);
  nand n564(x564, x15228, x469);
  nand n565(x565, x564, x563);
  nand n566(x566, x15229, x16472);
  nand n567(x567, x15228, x472);
  nand n568(x568, x567, x566);
  nand n569(x569, x15229, x16475);
  nand n570(x570, x15228, x475);
  nand n571(x571, x570, x569);
  nand n572(x572, x15229, x16478);
  nand n573(x573, x15228, x478);
  nand n574(x574, x573, x572);
  nand n575(x575, x15229, x16481);
  nand n576(x576, x15228, x481);
  nand n577(x577, x576, x575);
  nand n578(x578, x15229, x16484);
  nand n579(x579, x15228, x484);
  nand n580(x580, x579, x578);
  nand n581(x581, x15229, x16487);
  nand n582(x582, x15228, x487);
  nand n583(x583, x582, x581);
  nand n584(x584, x15229, x16490);
  nand n585(x585, x15228, x490);
  nand n586(x586, x585, x584);
  nand n587(x587, x15229, x16493);
  nand n588(x588, x15228, x493);
  nand n589(x589, x588, x587);
  nand n590(x590, x15229, x16496);
  nand n591(x591, x15228, x496);
  nand n592(x592, x591, x590);
  nand n593(x593, x15229, x16499);
  nand n594(x594, x15228, x499);
  nand n595(x595, x594, x593);
  nand n596(x596, x15229, x16502);
  nand n597(x597, x15228, x502);
  nand n598(x598, x597, x596);
  nand n599(x599, x15229, x16505);
  nand n600(x600, x15228, x505);
  nand n601(x601, x600, x599);
  nand n638(x638, x675, x674);
  nand n639(x639, x676, x675);
  nand n641(x641, x640, x674);
  nand n642(x642, x634, x637);
  nand n643(x643, x642, x638);
  nand n645(x645, x676, x83415);
  nand n646(x646, x635, x638);
  nand n647(x647, x646, x645);
  nand n649(x649, x677, x83416);
  nand n650(x650, x636, x641);
  nand n651(x651, x650, x649);
  nand n653(x653, x635, x677);
  nand n655(x655, x674, x634);
  nand n657(x657, x656, x654);
  nand n658(x658, x657, x637);
  nand n659(x659, x657, x644);
  nand n660(x660, x657, x648);
  nand n661(x661, x657, x652);
  nand n662(x662, x71140, x674);
  nand n663(x663, x1, x83417);
  nand n664(x664, x663, x662);
  nand n665(x665, x71140, x675);
  nand n666(x666, x1, x83418);
  nand n667(x667, x666, x665);
  nand n668(x668, x71140, x676);
  nand n669(x669, x1, x83419);
  nand n670(x670, x669, x668);
  nand n671(x671, x71140, x677);
  nand n672(x672, x1, x83420);
  nand n673(x673, x672, x671);
  nand n679(x679, x604, x93);
  nand n680(x680, x605, x679);
  nand n681(x681, x64, x604);
  nand n682(x682, x606, x83421);
  nand n683(x683, x606, x83422);
  nand n684(x684, x65, x83421);
  nand n685(x685, x684, x683);
  nand n686(x686, x65, x83423);
  nand n687(x687, x607, x83424);
  nand n688(x688, x66, x685);
  nand n689(x689, x688, x687);
  nand n690(x690, x66, x83425);
  nand n691(x691, x608, x689);
  nand n692(x692, x67, x83426);
  nand n693(x693, x692, x691);
  nand n694(x694, x68, x693);
  nand n695(x695, x69, x83427);
  nand n696(x696, x70, x83428);
  nand n697(x697, x606, x83423);
  nand n698(x698, x65, x83387);
  nand n699(x699, x698, x697);
  nand n700(x700, x66, x83430);
  nand n701(x701, x66, x699);
  nand n702(x702, x608, x83431);
  nand n703(x703, x67, x83432);
  nand n704(x704, x703, x702);
  nand n705(x705, x68, x704);
  nand n706(x706, x69, x83433);
  nand n707(x707, x70, x83434);
  nand n708(x708, x605, x93);
  nand n709(x709, x64, x679);
  nand n710(x710, x65, x83436);
  nand n711(x711, x710, x683);
  nand n712(x712, x606, x83436);
  nand n713(x713, x65, x83437);
  nand n714(x714, x713, x712);
  nand n715(x715, x607, x83430);
  nand n716(x716, x66, x711);
  nand n717(x717, x716, x715);
  nand n718(x718, x607, x714);
  nand n719(x719, x66, x83438);
  nand n720(x720, x719, x718);
  nand n721(x721, x608, x717);
  nand n722(x722, x67, x720);
  nand n723(x723, x722, x721);
  nand n724(x724, x68, x723);
  nand n725(x725, x69, x83439);
  nand n726(x726, x70, x83440);
  nand n727(x727, x681, x708);
  nand n728(x728, x65, x727);
  nand n729(x729, x606, x727);
  nand n730(x730, x66, x83442);
  nand n731(x731, x730, x715);
  nand n732(x732, x607, x83443);
  nand n733(x733, x66, x83444);
  nand n734(x734, x733, x732);
  nand n735(x735, x608, x731);
  nand n736(x736, x67, x734);
  nand n737(x737, x736, x735);
  nand n738(x738, x68, x737);
  nand n739(x739, x69, x83445);
  nand n740(x740, x70, x83446);
  nand n741(x741, x66, x83448);
  nand n742(x742, x741, x715);
  nand n743(x743, x608, x742);
  nand n744(x744, x67, x83449);
  nand n745(x745, x744, x743);
  nand n746(x746, x68, x745);
  nand n747(x747, x69, x83450);
  nand n748(x748, x70, x83451);
  nand n749(x749, x686, x297);
  nand n750(x750, x607, x749);
  nand n751(x751, x67, x83453);
  nand n752(x752, x751, x735);
  nand n753(x753, x68, x752);
  nand n754(x754, x69, x83454);
  nand n755(x755, x70, x83455);
  nand n756(x756, x607, x83425);
  nand n757(x757, x719, x756);
  nand n758(x758, x67, x757);
  nand n759(x759, x758, x735);
  nand n760(x760, x68, x759);
  nand n761(x761, x69, x83457);
  nand n762(x762, x70, x83458);
  nand n763(x763, x681, x680);
  nand n764(x764, x65, x763);
  nand n765(x765, x66, x83460);
  nand n766(x766, x765, x715);
  nand n767(x767, x608, x766);
  nand n768(x768, x67, x83461);
  nand n769(x769, x768, x767);
  nand n770(x770, x68, x769);
  nand n771(x771, x69, x83462);
  nand n772(x772, x70, x83463);
  nand n773(x773, x294, x708);
  nand n774(x774, x606, x83437);
  nand n775(x775, x65, x773);
  nand n776(x776, x775, x774);
  nand n777(x777, x686, x697);
  nand n778(x778, x607, x776);
  nand n779(x779, x765, x778);
  nand n780(x780, x607, x777);
  nand n781(x781, x608, x779);
  nand n782(x782, x67, x83465);
  nand n783(x783, x782, x781);
  nand n784(x784, x68, x783);
  nand n785(x785, x69, x83466);
  nand n786(x786, x70, x83467);
  nand n787(x787, x775, x697);
  nand n788(x788, x607, x787);
  nand n789(x789, x765, x788);
  nand n790(x790, x608, x789);
  nand n791(x791, x768, x790);
  nand n792(x792, x68, x791);
  nand n793(x793, x69, x83469);
  nand n794(x794, x70, x83470);
  nand n795(x795, x709, x94);
  nand n796(x796, x709, x680);
  nand n797(x797, x606, x795);
  nand n798(x798, x764, x797);
  nand n799(x799, x606, x773);
  nand n800(x800, x65, x796);
  nand n801(x801, x800, x799);
  nand n802(x802, x607, x798);
  nand n803(x803, x66, x801);
  nand n804(x804, x803, x802);
  nand n805(x805, x66, x83472);
  nand n806(x806, x805, x780);
  nand n807(x807, x608, x804);
  nand n808(x808, x67, x806);
  nand n809(x809, x808, x807);
  nand n810(x810, x68, x809);
  nand n811(x811, x69, x83473);
  nand n812(x812, x70, x83474);
  nand n813(x813, x65, x295);
  nand n814(x814, x813, x774);
  nand n815(x815, x606, x295);
  nand n816(x816, x65, x795);
  nand n817(x817, x816, x815);
  nand n818(x818, x607, x814);
  nand n819(x819, x66, x817);
  nand n820(x820, x819, x818);
  nand n821(x821, x66, x83476);
  nand n822(x822, x821, x756);
  nand n823(x823, x608, x820);
  nand n824(x824, x67, x822);
  nand n825(x825, x824, x823);
  nand n826(x826, x68, x825);
  nand n827(x827, x69, x83477);
  nand n828(x828, x70, x83478);
  nand n829(x829, x709, x708);
  nand n830(x830, x681, x94);
  nand n831(x831, x65, x829);
  nand n832(x832, x831, x774);
  nand n833(x833, x65, x830);
  nand n834(x834, x833, x729);
  nand n835(x835, x607, x832);
  nand n836(x836, x66, x834);
  nand n837(x837, x836, x835);
  nand n838(x838, x608, x837);
  nand n839(x839, x768, x838);
  nand n840(x840, x68, x839);
  nand n841(x841, x69, x83480);
  nand n842(x842, x70, x83481);
  nand n843(x843, x294, x680);
  nand n844(x844, x65, x843);
  nand n845(x845, x844, x797);
  nand n846(x846, x606, x830);
  nand n847(x847, x833, x846);
  nand n848(x848, x833, x797);
  nand n849(x849, x606, x843);
  nand n850(x850, x764, x849);
  nand n851(x851, x66, x83483);
  nand n852(x852, x607, x845);
  nand n853(x853, x66, x847);
  nand n854(x854, x853, x852);
  nand n855(x855, x607, x848);
  nand n856(x856, x66, x850);
  nand n857(x857, x856, x855);
  nand n858(x858, x67, x83484);
  nand n859(x859, x608, x854);
  nand n860(x860, x67, x857);
  nand n861(x861, x860, x859);
  nand n862(x862, x609, x83485);
  nand n863(x863, x68, x861);
  nand n864(x864, x863, x862);
  nand n865(x865, x69, x864);
  nand n866(x866, x70, x83486);
  nand n867(x867, x684, x774);
  nand n868(x868, x764, x682);
  nand n869(x869, x686, x815);
  nand n870(x870, x684, x729);
  nand n871(x871, x607, x867);
  nand n872(x872, x66, x868);
  nand n873(x873, x872, x871);
  nand n874(x874, x607, x869);
  nand n875(x875, x66, x870);
  nand n876(x876, x875, x874);
  nand n877(x877, x608, x873);
  nand n878(x878, x67, x876);
  nand n879(x879, x878, x877);
  nand n880(x880, x68, x879);
  nand n881(x881, x880, x862);
  nand n882(x882, x69, x881);
  nand n883(x883, x70, x83488);
  nand n884(x884, x831, x697);
  nand n885(x885, x606, x796);
  nand n886(x886, x686, x885);
  nand n887(x887, x607, x884);
  nand n888(x888, x66, x886);
  nand n889(x889, x888, x887);
  nand n890(x890, x608, x889);
  nand n891(x891, x768, x890);
  nand n892(x892, x68, x891);
  nand n893(x893, x69, x83490);
  nand n894(x894, x70, x83491);
  nand n895(x895, x844, x697);
  nand n896(x896, x833, x849);
  nand n897(x897, x800, x815);
  nand n898(x898, x800, x729);
  nand n899(x899, x607, x895);
  nand n900(x900, x66, x896);
  nand n901(x901, x900, x899);
  nand n902(x902, x607, x897);
  nand n903(x903, x66, x898);
  nand n904(x904, x903, x902);
  nand n905(x905, x608, x901);
  nand n906(x906, x67, x904);
  nand n907(x907, x906, x905);
  nand n908(x908, x68, x907);
  nand n909(x909, x69, x83493);
  nand n910(x910, x70, x83494);
  nand n911(x911, x775, x849);
  nand n912(x912, x710, x712);
  nand n913(x913, x607, x83448);
  nand n914(x914, x66, x911);
  nand n915(x915, x914, x913);
  nand n916(x916, x607, x83472);
  nand n917(x917, x66, x912);
  nand n918(x918, x917, x916);
  nand n919(x919, x608, x915);
  nand n920(x920, x67, x918);
  nand n921(x921, x920, x919);
  nand n922(x922, x68, x921);
  nand n923(x923, x922, x862);
  nand n924(x924, x69, x923);
  nand n925(x925, x70, x83496);
  nand n926(x926, x606, x763);
  nand n927(x927, x831, x926);
  nand n928(x928, x800, x683);
  nand n929(x929, x800, x682);
  nand n930(x930, x713, x797);
  nand n931(x931, x607, x927);
  nand n932(x932, x66, x928);
  nand n933(x933, x932, x931);
  nand n934(x934, x607, x929);
  nand n935(x935, x66, x930);
  nand n936(x936, x935, x934);
  nand n937(x937, x608, x933);
  nand n938(x938, x67, x936);
  nand n939(x939, x938, x937);
  nand n940(x940, x68, x939);
  nand n941(x941, x940, x862);
  nand n942(x942, x69, x941);
  nand n943(x943, x70, x83498);
  nand n944(x944, x713, x697);
  nand n945(x945, x698, x682);
  nand n946(x946, x66, x777);
  nand n947(x947, x946, x916);
  nand n948(x948, x607, x944);
  nand n949(x949, x66, x945);
  nand n950(x950, x949, x948);
  nand n951(x951, x608, x947);
  nand n952(x952, x67, x950);
  nand n953(x953, x952, x951);
  nand n954(x954, x68, x953);
  nand n955(x955, x954, x862);
  nand n956(x956, x69, x955);
  nand n957(x957, x70, x83500);
  nand n958(x958, x800, x885);
  nand n959(x959, x728, x885);
  nand n960(x960, x713, x682);
  nand n961(x961, x698, x729);
  nand n962(x962, x607, x958);
  nand n963(x963, x66, x959);
  nand n964(x964, x963, x962);
  nand n965(x965, x607, x960);
  nand n966(x966, x66, x961);
  nand n967(x967, x966, x965);
  nand n968(x968, x608, x964);
  nand n969(x969, x67, x967);
  nand n970(x970, x969, x968);
  nand n971(x971, x68, x970);
  nand n972(x972, x971, x862);
  nand n973(x973, x69, x972);
  nand n974(x974, x70, x83502);
  nand n975(x975, x813, x682);
  nand n976(x976, x831, x815);
  nand n977(x977, x607, x928);
  nand n978(x978, x66, x975);
  nand n979(x979, x978, x977);
  nand n980(x980, x607, x685);
  nand n981(x981, x66, x976);
  nand n982(x982, x981, x980);
  nand n983(x983, x608, x979);
  nand n984(x984, x67, x982);
  nand n985(x985, x984, x983);
  nand n986(x986, x68, x985);
  nand n987(x987, x69, x83504);
  nand n988(x988, x70, x83505);
  nand n989(x989, x65, x83422);
  nand n990(x990, x607, x83507);
  nand n991(x991, x67, x83508);
  nand n992(x992, x68, x83509);
  nand n993(x993, x69, x83510);
  nand n994(x994, x70, x83511);
  nand n995(x995, x608, x83426);
  nand n996(x996, x991, x995);
  nand n997(x997, x68, x996);
  nand n998(x998, x69, x83513);
  nand n999(x999, x70, x83514);
  nand n1002(x1002, x71265, x1001);
  nand n1004(x1004, x71255, x71260);
  nand n1006(x1006, x1000, x71250);
  nand n1008(x1008, x1005, x1003);
  nand n1010(x1010, x1009, x1007);
  nand n1013(x1013, x71265, x71270);
  nand n1015(x1015, x1012, x71260);
  nand n1017(x1017, x71245, x1011);
  nand n1019(x1019, x1016, x1014);
  nand n1021(x1021, x1020, x1018);
  nand n1023(x1023, x71255, x1022);
  nand n1025(x1025, x1000, x1011);
  nand n1027(x1027, x1024, x1014);
  nand n1029(x1029, x1028, x1026);
  nand n1030(x1030, x1012, x1022);
  nand n1032(x1032, x71245, x71250);
  nand n1034(x1034, x1031, x1014);
  nand n1036(x1036, x1035, x1033);
  nand n1037(x1037, x1009, x1026);
  nand n1039(x1039, x1038, x1001);
  nand n1041(x1041, x1024, x1040);
  nand n1043(x1043, x1042, x1007);
  nand n1044(x1044, x1042, x1018);
  nand n1045(x1045, x1044, x1043);
  nand n1047(x1047, x1046, x1037);
  nand n1049(x1049, x1048, x1036);
  nand n1051(x1051, x1050, x1029);
  nand n1053(x1053, x1052, x1021);
  nand n1054(x1054, x1020, x1026);
  nand n1055(x1055, x1028, x1033);
  nand n1056(x1056, x1028, x1007);
  nand n1057(x1057, x1028, x1018);
  nand n1058(x1058, x1031, x1003);
  nand n1060(x1060, x1059, x1026);
  nand n1061(x1061, x1005, x1040);
  nand n1063(x1063, x1062, x1033);
  nand n1064(x1064, x1062, x1007);
  nand n1065(x1065, x1062, x1018);
  nand n1066(x1066, x1062, x1026);
  nand n1067(x1067, x1016, x1040);
  nand n1069(x1069, x1068, x1033);
  nand n1070(x1070, x1068, x1007);
  nand n1071(x1071, x1068, x1018);
  nand n1072(x1072, x1068, x1026);
  nand n1073(x1073, x1042, x1033);
  nand n1074(x1074, x1073, x1072);
  nand n1076(x1076, x1075, x1071);
  nand n1078(x1078, x1077, x1070);
  nand n1080(x1080, x1079, x1069);
  nand n1082(x1082, x1081, x1066);
  nand n1084(x1084, x1083, x1065);
  nand n1086(x1086, x1085, x1064);
  nand n1088(x1088, x1087, x1063);
  nand n1090(x1090, x1089, x1060);
  nand n1092(x1092, x1091, x1057);
  nand n1094(x1094, x1093, x1056);
  nand n1096(x1096, x1095, x1055);
  nand n1098(x1098, x1097, x1054);
  nand n1099(x1099, x1009, x1018);
  nand n1100(x1100, x1038, x71270);
  nand n1102(x1102, x1024, x1101);
  nand n1104(x1104, x1103, x1018);
  nand n1105(x1105, x1016, x1003);
  nand n1107(x1107, x1106, x1033);
  nand n1108(x1108, x1107, x1104);
  nand n1109(x1109, x1031, x1101);
  nand n1111(x1111, x1110, x1033);
  nand n1112(x1112, x1106, x1007);
  nand n1113(x1113, x1106, x1018);
  nand n1114(x1114, x1106, x1026);
  nand n1115(x1115, x1024, x1003);
  nand n1117(x1117, x1116, x1033);
  nand n1118(x1118, x1116, x1007);
  nand n1119(x1119, x1116, x1018);
  nand n1120(x1120, x1116, x1026);
  nand n1121(x1121, x1059, x1033);
  nand n1122(x1122, x1059, x1007);
  nand n1123(x1123, x1059, x1018);
  nand n1124(x1124, x1123, x1122);
  nand n1126(x1126, x1125, x1121);
  nand n1128(x1128, x1127, x1120);
  nand n1130(x1130, x1129, x1119);
  nand n1132(x1132, x1131, x1118);
  nand n1134(x1134, x1133, x1117);
  nand n1136(x1136, x1135, x1114);
  nand n1138(x1138, x1137, x1113);
  nand n1140(x1140, x1139, x1112);
  nand n1142(x1142, x1141, x1111);
  nand n1143(x1143, x1103, x1026);
  nand n1144(x1144, x1005, x1101);
  nand n1146(x1146, x1145, x1026);
  nand n1147(x1147, x1016, x1101);
  nand n1149(x1149, x1148, x1033);
  nand n1150(x1150, x1103, x1007);
  nand n1151(x1151, x1150, x1149);
  nand n1153(x1153, x1152, x1146);
  nand n1154(x1154, x1148, x1007);
  nand n1155(x1155, x1148, x1018);
  nand n1156(x1156, x1148, x1026);
  nand n1157(x1157, x1103, x1033);
  nand n1158(x1158, x1157, x1156);
  nand n1160(x1160, x1159, x1155);
  nand n1165(x1165, x1162, x1161);
  nand n1166(x1166, x1099, x1163);
  nand n1167(x1167, x1010, x1164);
  nand n1171(x1171, x1170, x1169);
  nand n1173(x1173, x1172, x1168);
  nand n1174(x1174, x1154, x1161);
  nand n1176(x1176, x1175, x1163);
  nand n1178(x1178, x1177, x1164);
  nand n1182(x1182, x1181, x1180);
  nand n1184(x1184, x1183, x1179);
  nand n1185(x1185, x1099, x1180);
  nand n1187(x1187, x1143, x1162);
  nand n1189(x1189, x1188, x1179);
  nand n1191(x1191, x71122, x71124);
  nand n1192(x1192, x71118, x71120);
  nand n1195(x1195, x1194, x1193);
  nand n1197(x1197, x1196, x1195);
  nand n1199(x1199, x70929, x1195);
  nand n1202(x1202, x1201, x1198);
  nand n1204(x1204, x70913, x1198);
  nand n1206(x1206, x1201, x1200);
  nand n1208(x1208, x70913, x1200);
  nand n1211(x1211, x1210, x1203);
  nand n1213(x1213, x70897, x1203);
  nand n1215(x1215, x1210, x1205);
  nand n1217(x1217, x70897, x1205);
  nand n1219(x1219, x1210, x1207);
  nand n1221(x1221, x70897, x1207);
  nand n1223(x1223, x1210, x1209);
  nand n1225(x1225, x70897, x1209);
  nand n1227(x1227, x1212, x71119);
  nand n1229(x1229, x1228, x70833);
  nand n1230(x1230, x1227, x1232);
  nand n1231(x1231, x1230, x1229);
  nand n1233(x1233, x1214, x71119);
  nand n1235(x1235, x1234, x70833);
  nand n1236(x1236, x1233, x1238);
  nand n1237(x1237, x1236, x1235);
  nand n1239(x1239, x1216, x71119);
  nand n1241(x1241, x1240, x70833);
  nand n1242(x1242, x1239, x1244);
  nand n1243(x1243, x1242, x1241);
  nand n1245(x1245, x1218, x71119);
  nand n1247(x1247, x1246, x70833);
  nand n1248(x1248, x1245, x1250);
  nand n1249(x1249, x1248, x1247);
  nand n1251(x1251, x1220, x71119);
  nand n1253(x1253, x1252, x70833);
  nand n1254(x1254, x1251, x1256);
  nand n1255(x1255, x1254, x1253);
  nand n1257(x1257, x1222, x71119);
  nand n1259(x1259, x1258, x70833);
  nand n1260(x1260, x1257, x1262);
  nand n1261(x1261, x1260, x1259);
  nand n1263(x1263, x1224, x71119);
  nand n1265(x1265, x1264, x70833);
  nand n1266(x1266, x1263, x1268);
  nand n1267(x1267, x1266, x1265);
  nand n1269(x1269, x1226, x71119);
  nand n1271(x1271, x1270, x70833);
  nand n1272(x1272, x1269, x1274);
  nand n1273(x1273, x1272, x1271);
  nand n1275(x1275, x1212, x71121);
  nand n1277(x1277, x1276, x70849);
  nand n1278(x1278, x1275, x1282);
  nand n1279(x1279, x1278, x1277);
  nand n1283(x1283, x1214, x71121);
  nand n1285(x1285, x1284, x70849);
  nand n1286(x1286, x1283, x1288);
  nand n1287(x1287, x1286, x1285);
  nand n1289(x1289, x1216, x71121);
  nand n1291(x1291, x1290, x70849);
  nand n1292(x1292, x1289, x1294);
  nand n1293(x1293, x1292, x1291);
  nand n1295(x1295, x1218, x71121);
  nand n1297(x1297, x1296, x70849);
  nand n1298(x1298, x1295, x1300);
  nand n1299(x1299, x1298, x1297);
  nand n1301(x1301, x1220, x71121);
  nand n1303(x1303, x1302, x70849);
  nand n1304(x1304, x1301, x1306);
  nand n1305(x1305, x1304, x1303);
  nand n1307(x1307, x1222, x71121);
  nand n1309(x1309, x1308, x70849);
  nand n1310(x1310, x1307, x1312);
  nand n1311(x1311, x1310, x1309);
  nand n1313(x1313, x1224, x71121);
  nand n1315(x1315, x1314, x70849);
  nand n1316(x1316, x1313, x1318);
  nand n1317(x1317, x1316, x1315);
  nand n1319(x1319, x1226, x71121);
  nand n1321(x1321, x1320, x70849);
  nand n1322(x1322, x1319, x1324);
  nand n1323(x1323, x1322, x1321);
  nand n1325(x1325, x1212, x71123);
  nand n1327(x1327, x1326, x70865);
  nand n1328(x1328, x1325, x1330);
  nand n1329(x1329, x1328, x1327);
  nand n1331(x1331, x1214, x71123);
  nand n1333(x1333, x1332, x70865);
  nand n1334(x1334, x1331, x1336);
  nand n1335(x1335, x1334, x1333);
  nand n1337(x1337, x1216, x71123);
  nand n1339(x1339, x1338, x70865);
  nand n1340(x1340, x1337, x1342);
  nand n1341(x1341, x1340, x1339);
  nand n1343(x1343, x1218, x71123);
  nand n1345(x1345, x1344, x70865);
  nand n1346(x1346, x1343, x1348);
  nand n1347(x1347, x1346, x1345);
  nand n1349(x1349, x1220, x71123);
  nand n1351(x1351, x1350, x70865);
  nand n1352(x1352, x1349, x1354);
  nand n1353(x1353, x1352, x1351);
  nand n1355(x1355, x1222, x71123);
  nand n1357(x1357, x1356, x70865);
  nand n1358(x1358, x1355, x1360);
  nand n1359(x1359, x1358, x1357);
  nand n1361(x1361, x1224, x71123);
  nand n1363(x1363, x1362, x70865);
  nand n1364(x1364, x1361, x1366);
  nand n1365(x1365, x1364, x1363);
  nand n1367(x1367, x1226, x71123);
  nand n1369(x1369, x1368, x70865);
  nand n1370(x1370, x1367, x1372);
  nand n1371(x1371, x1370, x1369);
  nand n1373(x1373, x1212, x71125);
  nand n1375(x1375, x1374, x70881);
  nand n1376(x1376, x1373, x1380);
  nand n1377(x1377, x1376, x1375);
  nand n1381(x1381, x1214, x71125);
  nand n1383(x1383, x1382, x70881);
  nand n1384(x1384, x1381, x1386);
  nand n1385(x1385, x1384, x1383);
  nand n1387(x1387, x1216, x71125);
  nand n1389(x1389, x1388, x70881);
  nand n1390(x1390, x1387, x1392);
  nand n1391(x1391, x1390, x1389);
  nand n1393(x1393, x1218, x71125);
  nand n1395(x1395, x1394, x70881);
  nand n1396(x1396, x1393, x1398);
  nand n1397(x1397, x1396, x1395);
  nand n1399(x1399, x1220, x71125);
  nand n1401(x1401, x1400, x70881);
  nand n1402(x1402, x1399, x1404);
  nand n1403(x1403, x1402, x1401);
  nand n1405(x1405, x1222, x71125);
  nand n1407(x1407, x1406, x70881);
  nand n1408(x1408, x1405, x1410);
  nand n1409(x1409, x1408, x1407);
  nand n1411(x1411, x1224, x71125);
  nand n1413(x1413, x1412, x70881);
  nand n1414(x1414, x1411, x1416);
  nand n1415(x1415, x1414, x1413);
  nand n1417(x1417, x1226, x71125);
  nand n1419(x1419, x1418, x70881);
  nand n1420(x1420, x1417, x1422);
  nand n1421(x1421, x1420, x1419);
  nand n1423(x1423, x71215, x1274);
  nand n1425(x1425, x1424, x1268);
  nand n1426(x1426, x1425, x1423);
  nand n1427(x1427, x71215, x1262);
  nand n1428(x1428, x1424, x1256);
  nand n1429(x1429, x1428, x1427);
  nand n1430(x1430, x71215, x1250);
  nand n1431(x1431, x1424, x1244);
  nand n1432(x1432, x1431, x1430);
  nand n1433(x1433, x71215, x1238);
  nand n1434(x1434, x1424, x1232);
  nand n1435(x1435, x1434, x1433);
  nand n1436(x1436, x71220, x1426);
  nand n1438(x1438, x1437, x1429);
  nand n1439(x1439, x1438, x1436);
  nand n1440(x1440, x71220, x1432);
  nand n1441(x1441, x1437, x1435);
  nand n1442(x1442, x1441, x1440);
  nand n1443(x1443, x71225, x1439);
  nand n1445(x1445, x1444, x1442);
  nand n1446(x1446, x1445, x1443);
  nand n1447(x1447, x71202, x1274);
  nand n1449(x1449, x1448, x1268);
  nand n1450(x1450, x1449, x1447);
  nand n1451(x1451, x71202, x1262);
  nand n1452(x1452, x1448, x1256);
  nand n1453(x1453, x1452, x1451);
  nand n1454(x1454, x71202, x1250);
  nand n1455(x1455, x1448, x1244);
  nand n1456(x1456, x1455, x1454);
  nand n1457(x1457, x71202, x1238);
  nand n1458(x1458, x1448, x1232);
  nand n1459(x1459, x1458, x1457);
  nand n1460(x1460, x71205, x1450);
  nand n1462(x1462, x1461, x1453);
  nand n1463(x1463, x1462, x1460);
  nand n1464(x1464, x71205, x1456);
  nand n1465(x1465, x1461, x1459);
  nand n1466(x1466, x1465, x1464);
  nand n1467(x1467, x71210, x1463);
  nand n1469(x1469, x1468, x1466);
  nand n1470(x1470, x1469, x1467);
  nand n1471(x1471, x71275, x1274);
  nand n1473(x1473, x1472, x1268);
  nand n1474(x1474, x1473, x1471);
  nand n1475(x1475, x71275, x1262);
  nand n1476(x1476, x1472, x1256);
  nand n1477(x1477, x1476, x1475);
  nand n1478(x1478, x71275, x1250);
  nand n1479(x1479, x1472, x1244);
  nand n1480(x1480, x1479, x1478);
  nand n1481(x1481, x71275, x1238);
  nand n1482(x1482, x1472, x1232);
  nand n1483(x1483, x1482, x1481);
  nand n1484(x1484, x71277, x1474);
  nand n1486(x1486, x1485, x1477);
  nand n1487(x1487, x1486, x1484);
  nand n1488(x1488, x71277, x1480);
  nand n1489(x1489, x1485, x1483);
  nand n1490(x1490, x1489, x1488);
  nand n1491(x1491, x71279, x1487);
  nand n1493(x1493, x1492, x1490);
  nand n1494(x1494, x1493, x1491);
  nand n1495(x1495, x71215, x1324);
  nand n1496(x1496, x1424, x1318);
  nand n1497(x1497, x1496, x1495);
  nand n1498(x1498, x71215, x1312);
  nand n1499(x1499, x1424, x1306);
  nand n1500(x1500, x1499, x1498);
  nand n1501(x1501, x71215, x1300);
  nand n1502(x1502, x1424, x1294);
  nand n1503(x1503, x1502, x1501);
  nand n1504(x1504, x71215, x1288);
  nand n1505(x1505, x1424, x1282);
  nand n1506(x1506, x1505, x1504);
  nand n1507(x1507, x71220, x1497);
  nand n1508(x1508, x1437, x1500);
  nand n1509(x1509, x1508, x1507);
  nand n1510(x1510, x71220, x1503);
  nand n1511(x1511, x1437, x1506);
  nand n1512(x1512, x1511, x1510);
  nand n1513(x1513, x71225, x1509);
  nand n1514(x1514, x1444, x1512);
  nand n1515(x1515, x1514, x1513);
  nand n1516(x1516, x71202, x1324);
  nand n1517(x1517, x1448, x1318);
  nand n1518(x1518, x1517, x1516);
  nand n1519(x1519, x71202, x1312);
  nand n1520(x1520, x1448, x1306);
  nand n1521(x1521, x1520, x1519);
  nand n1522(x1522, x71202, x1300);
  nand n1523(x1523, x1448, x1294);
  nand n1524(x1524, x1523, x1522);
  nand n1525(x1525, x71202, x1288);
  nand n1526(x1526, x1448, x1282);
  nand n1527(x1527, x1526, x1525);
  nand n1528(x1528, x71205, x1518);
  nand n1529(x1529, x1461, x1521);
  nand n1530(x1530, x1529, x1528);
  nand n1531(x1531, x71205, x1524);
  nand n1532(x1532, x1461, x1527);
  nand n1533(x1533, x1532, x1531);
  nand n1534(x1534, x71210, x1530);
  nand n1535(x1535, x1468, x1533);
  nand n1536(x1536, x1535, x1534);
  nand n1537(x1537, x71275, x1324);
  nand n1538(x1538, x1472, x1318);
  nand n1539(x1539, x1538, x1537);
  nand n1540(x1540, x71275, x1312);
  nand n1541(x1541, x1472, x1306);
  nand n1542(x1542, x1541, x1540);
  nand n1543(x1543, x71275, x1300);
  nand n1544(x1544, x1472, x1294);
  nand n1545(x1545, x1544, x1543);
  nand n1546(x1546, x71275, x1288);
  nand n1547(x1547, x1472, x1282);
  nand n1548(x1548, x1547, x1546);
  nand n1549(x1549, x71277, x1539);
  nand n1550(x1550, x1485, x1542);
  nand n1551(x1551, x1550, x1549);
  nand n1552(x1552, x71277, x1545);
  nand n1553(x1553, x1485, x1548);
  nand n1554(x1554, x1553, x1552);
  nand n1555(x1555, x71279, x1551);
  nand n1556(x1556, x1492, x1554);
  nand n1557(x1557, x1556, x1555);
  nand n1558(x1558, x71215, x1372);
  nand n1559(x1559, x1424, x1366);
  nand n1560(x1560, x1559, x1558);
  nand n1561(x1561, x71215, x1360);
  nand n1562(x1562, x1424, x1354);
  nand n1563(x1563, x1562, x1561);
  nand n1564(x1564, x71215, x1348);
  nand n1565(x1565, x1424, x1342);
  nand n1566(x1566, x1565, x1564);
  nand n1567(x1567, x71215, x1336);
  nand n1568(x1568, x1424, x1330);
  nand n1569(x1569, x1568, x1567);
  nand n1570(x1570, x71220, x1560);
  nand n1571(x1571, x1437, x1563);
  nand n1572(x1572, x1571, x1570);
  nand n1573(x1573, x71220, x1566);
  nand n1574(x1574, x1437, x1569);
  nand n1575(x1575, x1574, x1573);
  nand n1576(x1576, x71225, x1572);
  nand n1577(x1577, x1444, x1575);
  nand n1578(x1578, x1577, x1576);
  nand n1579(x1579, x71202, x1372);
  nand n1580(x1580, x1448, x1366);
  nand n1581(x1581, x1580, x1579);
  nand n1582(x1582, x71202, x1360);
  nand n1583(x1583, x1448, x1354);
  nand n1584(x1584, x1583, x1582);
  nand n1585(x1585, x71202, x1348);
  nand n1586(x1586, x1448, x1342);
  nand n1587(x1587, x1586, x1585);
  nand n1588(x1588, x71202, x1336);
  nand n1589(x1589, x1448, x1330);
  nand n1590(x1590, x1589, x1588);
  nand n1591(x1591, x71205, x1581);
  nand n1592(x1592, x1461, x1584);
  nand n1593(x1593, x1592, x1591);
  nand n1594(x1594, x71205, x1587);
  nand n1595(x1595, x1461, x1590);
  nand n1596(x1596, x1595, x1594);
  nand n1597(x1597, x71210, x1593);
  nand n1598(x1598, x1468, x1596);
  nand n1599(x1599, x1598, x1597);
  nand n1600(x1600, x71275, x1372);
  nand n1601(x1601, x1472, x1366);
  nand n1602(x1602, x1601, x1600);
  nand n1603(x1603, x71275, x1360);
  nand n1604(x1604, x1472, x1354);
  nand n1605(x1605, x1604, x1603);
  nand n1606(x1606, x71275, x1348);
  nand n1607(x1607, x1472, x1342);
  nand n1608(x1608, x1607, x1606);
  nand n1609(x1609, x71275, x1336);
  nand n1610(x1610, x1472, x1330);
  nand n1611(x1611, x1610, x1609);
  nand n1612(x1612, x71277, x1602);
  nand n1613(x1613, x1485, x1605);
  nand n1614(x1614, x1613, x1612);
  nand n1615(x1615, x71277, x1608);
  nand n1616(x1616, x1485, x1611);
  nand n1617(x1617, x1616, x1615);
  nand n1618(x1618, x71279, x1614);
  nand n1619(x1619, x1492, x1617);
  nand n1620(x1620, x1619, x1618);
  nand n1621(x1621, x71215, x1422);
  nand n1622(x1622, x1424, x1416);
  nand n1623(x1623, x1622, x1621);
  nand n1624(x1624, x71215, x1410);
  nand n1625(x1625, x1424, x1404);
  nand n1626(x1626, x1625, x1624);
  nand n1627(x1627, x71215, x1398);
  nand n1628(x1628, x1424, x1392);
  nand n1629(x1629, x1628, x1627);
  nand n1630(x1630, x71215, x1386);
  nand n1631(x1631, x1424, x1380);
  nand n1632(x1632, x1631, x1630);
  nand n1633(x1633, x71220, x1623);
  nand n1634(x1634, x1437, x1626);
  nand n1635(x1635, x1634, x1633);
  nand n1636(x1636, x71220, x1629);
  nand n1637(x1637, x1437, x1632);
  nand n1638(x1638, x1637, x1636);
  nand n1639(x1639, x71225, x1635);
  nand n1640(x1640, x1444, x1638);
  nand n1641(x1641, x1640, x1639);
  nand n1642(x1642, x71202, x1422);
  nand n1643(x1643, x1448, x1416);
  nand n1644(x1644, x1643, x1642);
  nand n1645(x1645, x71202, x1410);
  nand n1646(x1646, x1448, x1404);
  nand n1647(x1647, x1646, x1645);
  nand n1648(x1648, x71202, x1398);
  nand n1649(x1649, x1448, x1392);
  nand n1650(x1650, x1649, x1648);
  nand n1651(x1651, x71202, x1386);
  nand n1652(x1652, x1448, x1380);
  nand n1653(x1653, x1652, x1651);
  nand n1654(x1654, x71205, x1644);
  nand n1655(x1655, x1461, x1647);
  nand n1656(x1656, x1655, x1654);
  nand n1657(x1657, x71205, x1650);
  nand n1658(x1658, x1461, x1653);
  nand n1659(x1659, x1658, x1657);
  nand n1660(x1660, x71210, x1656);
  nand n1661(x1661, x1468, x1659);
  nand n1662(x1662, x1661, x1660);
  nand n1663(x1663, x71275, x1422);
  nand n1664(x1664, x1472, x1416);
  nand n1665(x1665, x1664, x1663);
  nand n1666(x1666, x71275, x1410);
  nand n1667(x1667, x1472, x1404);
  nand n1668(x1668, x1667, x1666);
  nand n1669(x1669, x71275, x1398);
  nand n1670(x1670, x1472, x1392);
  nand n1671(x1671, x1670, x1669);
  nand n1672(x1672, x71275, x1386);
  nand n1673(x1673, x1472, x1380);
  nand n1674(x1674, x1673, x1672);
  nand n1675(x1675, x71277, x1665);
  nand n1676(x1676, x1485, x1668);
  nand n1677(x1677, x1676, x1675);
  nand n1678(x1678, x71277, x1671);
  nand n1679(x1679, x1485, x1674);
  nand n1680(x1680, x1679, x1678);
  nand n1681(x1681, x71279, x1677);
  nand n1682(x1682, x1492, x1680);
  nand n1683(x1683, x1682, x1681);
  nand n1685(x1685, x71284, x1684);
  nand n1687(x1687, x71284, x1686);
  nand n1689(x1689, x71284, x1688);
  nand n1691(x1691, x71284, x1690);
  nand n1692(x1692, x71449, x1685);
  nand n1694(x1694, x71449, x1687);
  nand n1696(x1696, x71449, x1689);
  nand n1698(x1698, x71449, x1691);
  nand n1700(x1700, x1186, x1189);
  nand n1702(x1702, x1173, x1184);
  nand n1704(x1704, x1703, x1701);
  nand n1706(x1706, x1705, x1184);
  nand n1708(x1708, x1707, x1701);
  nand n1710(x1710, x1173, x1709);
  nand n1712(x1712, x1711, x1701);
  nand n1713(x1713, x1712, x1708);
  nand n1715(x1715, x1714, x1704);
  nand n1716(x1716, x1715, x1);
  nand n1718(x1718, x1693, x1717);
  nand n1719(x1719, x1695, x1717);
  nand n1720(x1720, x1697, x1717);
  nand n1721(x1721, x1699, x1717);
  nand n1722(x1722, x1720, x1721);
  nand n1723(x1723, x1718, x1719);
  nand n1726(x1726, x1725, x1724);
  nand n1728(x1728, x1727, x1726);
  nand n1730(x1730, x71240, x1726);
  nand n1733(x1733, x1732, x1729);
  nand n1735(x1735, x71235, x1729);
  nand n1737(x1737, x1732, x1731);
  nand n1739(x1739, x71235, x1731);
  nand n1742(x1742, x1741, x1734);
  nand n1743(x1743, x71230, x1734);
  nand n1744(x1744, x1741, x1736);
  nand n1745(x1745, x71230, x1736);
  nand n1746(x1746, x1741, x1738);
  nand n1747(x1747, x71230, x1738);
  nand n1748(x1748, x1741, x1740);
  nand n1749(x1749, x71230, x1740);
  nand n1750(x1750, x1212, x1742);
  nand n1752(x1752, x1211, x1742);
  nand n1753(x1753, x1752, x1751);
  nand n1755(x1755, x1754, x1759);
  nand n1756(x1756, x1755, x1753);
  nand n1760(x1760, x1214, x1743);
  nand n1762(x1762, x1213, x1743);
  nand n1763(x1763, x1762, x1761);
  nand n1765(x1765, x1764, x1769);
  nand n1766(x1766, x1765, x1763);
  nand n1770(x1770, x1216, x1744);
  nand n1772(x1772, x1215, x1744);
  nand n1773(x1773, x1772, x1771);
  nand n1775(x1775, x1774, x1779);
  nand n1776(x1776, x1775, x1773);
  nand n1780(x1780, x1218, x1745);
  nand n1782(x1782, x1217, x1745);
  nand n1783(x1783, x1782, x1781);
  nand n1785(x1785, x1784, x1789);
  nand n1786(x1786, x1785, x1783);
  nand n1790(x1790, x1220, x1746);
  nand n1792(x1792, x1219, x1746);
  nand n1793(x1793, x1792, x1791);
  nand n1795(x1795, x1794, x1799);
  nand n1796(x1796, x1795, x1793);
  nand n1800(x1800, x1222, x1747);
  nand n1802(x1802, x1221, x1747);
  nand n1803(x1803, x1802, x1801);
  nand n1805(x1805, x1804, x1809);
  nand n1806(x1806, x1805, x1803);
  nand n1810(x1810, x1224, x1748);
  nand n1812(x1812, x1223, x1748);
  nand n1813(x1813, x1812, x1811);
  nand n1815(x1815, x1814, x1819);
  nand n1816(x1816, x1815, x1813);
  nand n1820(x1820, x1226, x1749);
  nand n1822(x1822, x1225, x1749);
  nand n1823(x1823, x1822, x1821);
  nand n1825(x1825, x1824, x1829);
  nand n1826(x1826, x1825, x1823);
  nand n1830(x1830, x71215, x1829);
  nand n1831(x1831, x1424, x1819);
  nand n1832(x1832, x1831, x1830);
  nand n1833(x1833, x71215, x1809);
  nand n1834(x1834, x1424, x1799);
  nand n1835(x1835, x1834, x1833);
  nand n1836(x1836, x71215, x1789);
  nand n1837(x1837, x1424, x1779);
  nand n1838(x1838, x1837, x1836);
  nand n1839(x1839, x71215, x1769);
  nand n1840(x1840, x1424, x1759);
  nand n1841(x1841, x1840, x1839);
  nand n1842(x1842, x71220, x1832);
  nand n1843(x1843, x1437, x1835);
  nand n1844(x1844, x1843, x1842);
  nand n1845(x1845, x71220, x1838);
  nand n1846(x1846, x1437, x1841);
  nand n1847(x1847, x1846, x1845);
  nand n1848(x1848, x71225, x1844);
  nand n1849(x1849, x1444, x1847);
  nand n1850(x1850, x1849, x1848);
  nand n1851(x1851, x71202, x1829);
  nand n1852(x1852, x1448, x1819);
  nand n1853(x1853, x1852, x1851);
  nand n1854(x1854, x71202, x1809);
  nand n1855(x1855, x1448, x1799);
  nand n1856(x1856, x1855, x1854);
  nand n1857(x1857, x71202, x1789);
  nand n1858(x1858, x1448, x1779);
  nand n1859(x1859, x1858, x1857);
  nand n1860(x1860, x71202, x1769);
  nand n1861(x1861, x1448, x1759);
  nand n1862(x1862, x1861, x1860);
  nand n1863(x1863, x71205, x1853);
  nand n1864(x1864, x1461, x1856);
  nand n1865(x1865, x1864, x1863);
  nand n1866(x1866, x71205, x1859);
  nand n1867(x1867, x1461, x1862);
  nand n1868(x1868, x1867, x1866);
  nand n1869(x1869, x71210, x1865);
  nand n1870(x1870, x1468, x1868);
  nand n1871(x1871, x1870, x1869);
  nand n1872(x1872, x71275, x1829);
  nand n1873(x1873, x1472, x1819);
  nand n1874(x1874, x1873, x1872);
  nand n1875(x1875, x71275, x1809);
  nand n1876(x1876, x1472, x1799);
  nand n1877(x1877, x1876, x1875);
  nand n1878(x1878, x71275, x1789);
  nand n1879(x1879, x1472, x1779);
  nand n1880(x1880, x1879, x1878);
  nand n1881(x1881, x71275, x1769);
  nand n1882(x1882, x1472, x1759);
  nand n1883(x1883, x1882, x1881);
  nand n1884(x1884, x71277, x1874);
  nand n1885(x1885, x1485, x1877);
  nand n1886(x1886, x1885, x1884);
  nand n1887(x1887, x71277, x1880);
  nand n1888(x1888, x1485, x1883);
  nand n1889(x1889, x1888, x1887);
  nand n1890(x1890, x71279, x1886);
  nand n1891(x1891, x1492, x1889);
  nand n1892(x1892, x1891, x1890);
  nand n1894(x1894, x1708, x1704);
  nand n1895(x1895, x1894, x1893);
  nand n1898(x1898, x1897, x1896);
  nand n1900(x1900, x71284, x1899);
  nand n1909(x1909, x1901, x1726);
  nand n1911(x1911, x1910, x71454);
  nand n1912(x1912, x1909, x1914);
  nand n1913(x1913, x1912, x1911);
  nand n1915(x1915, x1910, x71459);
  nand n1916(x1916, x1909, x1918);
  nand n1917(x1917, x1916, x1915);
  nand n1919(x1919, x1910, x71464);
  nand n1920(x1920, x1909, x1922);
  nand n1921(x1921, x1920, x1919);
  nand n1923(x1923, x1910, x71469);
  nand n1924(x1924, x1909, x1926);
  nand n1925(x1925, x1924, x1923);
  nand n1927(x1927, x1910, x71474);
  nand n1928(x1928, x1909, x1930);
  nand n1929(x1929, x1928, x1927);
  nand n1931(x1931, x1910, x71479);
  nand n1932(x1932, x1909, x1934);
  nand n1933(x1933, x1932, x1931);
  nand n1935(x1935, x1902, x1726);
  nand n1937(x1937, x1936, x71454);
  nand n1938(x1938, x1935, x1940);
  nand n1939(x1939, x1938, x1937);
  nand n1941(x1941, x1936, x71459);
  nand n1942(x1942, x1935, x1944);
  nand n1943(x1943, x1942, x1941);
  nand n1945(x1945, x1936, x71464);
  nand n1946(x1946, x1935, x1948);
  nand n1947(x1947, x1946, x1945);
  nand n1949(x1949, x1936, x71469);
  nand n1950(x1950, x1935, x1952);
  nand n1951(x1951, x1950, x1949);
  nand n1953(x1953, x1936, x71474);
  nand n1954(x1954, x1935, x1956);
  nand n1955(x1955, x1954, x1953);
  nand n1957(x1957, x1936, x71479);
  nand n1958(x1958, x1935, x1960);
  nand n1959(x1959, x1958, x1957);
  nand n1961(x1961, x1903, x1726);
  nand n1963(x1963, x1962, x71454);
  nand n1964(x1964, x1961, x1966);
  nand n1965(x1965, x1964, x1963);
  nand n1967(x1967, x1962, x71459);
  nand n1968(x1968, x1961, x1970);
  nand n1969(x1969, x1968, x1967);
  nand n1971(x1971, x1962, x71464);
  nand n1972(x1972, x1961, x1974);
  nand n1973(x1973, x1972, x1971);
  nand n1975(x1975, x1962, x71469);
  nand n1976(x1976, x1961, x1978);
  nand n1977(x1977, x1976, x1975);
  nand n1979(x1979, x1962, x71474);
  nand n1980(x1980, x1961, x1982);
  nand n1981(x1981, x1980, x1979);
  nand n1983(x1983, x1962, x71479);
  nand n1984(x1984, x1961, x1986);
  nand n1985(x1985, x1984, x1983);
  nand n1987(x1987, x1904, x1726);
  nand n1989(x1989, x1988, x71454);
  nand n1990(x1990, x1987, x1992);
  nand n1991(x1991, x1990, x1989);
  nand n1993(x1993, x1988, x71459);
  nand n1994(x1994, x1987, x1996);
  nand n1995(x1995, x1994, x1993);
  nand n1997(x1997, x1988, x71464);
  nand n1998(x1998, x1987, x2000);
  nand n1999(x1999, x1998, x1997);
  nand n2001(x2001, x1988, x71469);
  nand n2002(x2002, x1987, x2004);
  nand n2003(x2003, x2002, x2001);
  nand n2005(x2005, x1988, x71474);
  nand n2006(x2006, x1987, x2008);
  nand n2007(x2007, x2006, x2005);
  nand n2009(x2009, x1988, x71479);
  nand n2010(x2010, x1987, x2012);
  nand n2011(x2011, x2010, x2009);
  nand n2013(x2013, x1905, x1726);
  nand n2015(x2015, x2014, x71454);
  nand n2016(x2016, x2013, x2018);
  nand n2017(x2017, x2016, x2015);
  nand n2019(x2019, x2014, x71459);
  nand n2020(x2020, x2013, x2022);
  nand n2021(x2021, x2020, x2019);
  nand n2023(x2023, x2014, x71464);
  nand n2024(x2024, x2013, x2026);
  nand n2025(x2025, x2024, x2023);
  nand n2027(x2027, x2014, x71469);
  nand n2028(x2028, x2013, x2030);
  nand n2029(x2029, x2028, x2027);
  nand n2031(x2031, x2014, x71474);
  nand n2032(x2032, x2013, x2034);
  nand n2033(x2033, x2032, x2031);
  nand n2035(x2035, x2014, x71479);
  nand n2036(x2036, x2013, x2038);
  nand n2037(x2037, x2036, x2035);
  nand n2039(x2039, x1906, x1726);
  nand n2041(x2041, x2040, x71454);
  nand n2042(x2042, x2039, x2044);
  nand n2043(x2043, x2042, x2041);
  nand n2045(x2045, x2040, x71459);
  nand n2046(x2046, x2039, x2048);
  nand n2047(x2047, x2046, x2045);
  nand n2049(x2049, x2040, x71464);
  nand n2050(x2050, x2039, x2052);
  nand n2051(x2051, x2050, x2049);
  nand n2053(x2053, x2040, x71469);
  nand n2054(x2054, x2039, x2056);
  nand n2055(x2055, x2054, x2053);
  nand n2057(x2057, x2040, x71474);
  nand n2058(x2058, x2039, x2060);
  nand n2059(x2059, x2058, x2057);
  nand n2061(x2061, x2040, x71479);
  nand n2062(x2062, x2039, x2064);
  nand n2063(x2063, x2062, x2061);
  nand n2065(x2065, x1907, x1726);
  nand n2067(x2067, x2066, x71454);
  nand n2068(x2068, x2065, x2070);
  nand n2069(x2069, x2068, x2067);
  nand n2071(x2071, x2066, x71459);
  nand n2072(x2072, x2065, x2074);
  nand n2073(x2073, x2072, x2071);
  nand n2075(x2075, x2066, x71464);
  nand n2076(x2076, x2065, x2078);
  nand n2077(x2077, x2076, x2075);
  nand n2079(x2079, x2066, x71469);
  nand n2080(x2080, x2065, x2082);
  nand n2081(x2081, x2080, x2079);
  nand n2083(x2083, x2066, x71474);
  nand n2084(x2084, x2065, x2086);
  nand n2085(x2085, x2084, x2083);
  nand n2087(x2087, x2066, x71479);
  nand n2088(x2088, x2065, x2090);
  nand n2089(x2089, x2088, x2087);
  nand n2091(x2091, x1908, x1726);
  nand n2093(x2093, x2092, x71454);
  nand n2094(x2094, x2091, x2096);
  nand n2095(x2095, x2094, x2093);
  nand n2097(x2097, x2092, x71459);
  nand n2098(x2098, x2091, x2100);
  nand n2099(x2099, x2098, x2097);
  nand n2101(x2101, x2092, x71464);
  nand n2102(x2102, x2091, x2104);
  nand n2103(x2103, x2102, x2101);
  nand n2105(x2105, x2092, x71469);
  nand n2106(x2106, x2091, x2108);
  nand n2107(x2107, x2106, x2105);
  nand n2109(x2109, x2092, x71474);
  nand n2110(x2110, x2091, x2112);
  nand n2111(x2111, x2110, x2109);
  nand n2113(x2113, x2092, x71479);
  nand n2114(x2114, x2091, x2116);
  nand n2115(x2115, x2114, x2113);
  nand n2117(x2117, x70897, x2096);
  nand n2118(x2118, x1210, x2070);
  nand n2119(x2119, x2118, x2117);
  nand n2120(x2120, x70897, x2044);
  nand n2121(x2121, x1210, x2018);
  nand n2122(x2122, x2121, x2120);
  nand n2123(x2123, x70897, x1992);
  nand n2124(x2124, x1210, x1966);
  nand n2125(x2125, x2124, x2123);
  nand n2126(x2126, x70897, x1940);
  nand n2127(x2127, x1210, x1914);
  nand n2128(x2128, x2127, x2126);
  nand n2129(x2129, x70913, x2119);
  nand n2130(x2130, x1201, x2122);
  nand n2131(x2131, x2130, x2129);
  nand n2132(x2132, x70913, x2125);
  nand n2133(x2133, x1201, x2128);
  nand n2134(x2134, x2133, x2132);
  nand n2135(x2135, x70929, x2131);
  nand n2136(x2136, x1196, x2134);
  nand n2137(x2137, x2136, x2135);
  nand n2138(x2138, x70897, x2100);
  nand n2139(x2139, x1210, x2074);
  nand n2140(x2140, x2139, x2138);
  nand n2141(x2141, x70897, x2048);
  nand n2142(x2142, x1210, x2022);
  nand n2143(x2143, x2142, x2141);
  nand n2144(x2144, x70897, x1996);
  nand n2145(x2145, x1210, x1970);
  nand n2146(x2146, x2145, x2144);
  nand n2147(x2147, x70897, x1944);
  nand n2148(x2148, x1210, x1918);
  nand n2149(x2149, x2148, x2147);
  nand n2150(x2150, x70913, x2140);
  nand n2151(x2151, x1201, x2143);
  nand n2152(x2152, x2151, x2150);
  nand n2153(x2153, x70913, x2146);
  nand n2154(x2154, x1201, x2149);
  nand n2155(x2155, x2154, x2153);
  nand n2156(x2156, x70929, x2152);
  nand n2157(x2157, x1196, x2155);
  nand n2158(x2158, x2157, x2156);
  nand n2159(x2159, x70897, x2104);
  nand n2160(x2160, x1210, x2078);
  nand n2161(x2161, x2160, x2159);
  nand n2162(x2162, x70897, x2052);
  nand n2163(x2163, x1210, x2026);
  nand n2164(x2164, x2163, x2162);
  nand n2165(x2165, x70897, x2000);
  nand n2166(x2166, x1210, x1974);
  nand n2167(x2167, x2166, x2165);
  nand n2168(x2168, x70897, x1948);
  nand n2169(x2169, x1210, x1922);
  nand n2170(x2170, x2169, x2168);
  nand n2171(x2171, x70913, x2161);
  nand n2172(x2172, x1201, x2164);
  nand n2173(x2173, x2172, x2171);
  nand n2174(x2174, x70913, x2167);
  nand n2175(x2175, x1201, x2170);
  nand n2176(x2176, x2175, x2174);
  nand n2177(x2177, x70929, x2173);
  nand n2178(x2178, x1196, x2176);
  nand n2179(x2179, x2178, x2177);
  nand n2180(x2180, x70897, x2108);
  nand n2181(x2181, x1210, x2082);
  nand n2182(x2182, x2181, x2180);
  nand n2183(x2183, x70897, x2056);
  nand n2184(x2184, x1210, x2030);
  nand n2185(x2185, x2184, x2183);
  nand n2186(x2186, x70897, x2004);
  nand n2187(x2187, x1210, x1978);
  nand n2188(x2188, x2187, x2186);
  nand n2189(x2189, x70897, x1952);
  nand n2190(x2190, x1210, x1926);
  nand n2191(x2191, x2190, x2189);
  nand n2192(x2192, x70913, x2182);
  nand n2193(x2193, x1201, x2185);
  nand n2194(x2194, x2193, x2192);
  nand n2195(x2195, x70913, x2188);
  nand n2196(x2196, x1201, x2191);
  nand n2197(x2197, x2196, x2195);
  nand n2198(x2198, x70929, x2194);
  nand n2199(x2199, x1196, x2197);
  nand n2200(x2200, x2199, x2198);
  nand n2201(x2201, x70897, x2112);
  nand n2202(x2202, x1210, x2086);
  nand n2203(x2203, x2202, x2201);
  nand n2204(x2204, x70897, x2060);
  nand n2205(x2205, x1210, x2034);
  nand n2206(x2206, x2205, x2204);
  nand n2207(x2207, x70897, x2008);
  nand n2208(x2208, x1210, x1982);
  nand n2209(x2209, x2208, x2207);
  nand n2210(x2210, x70897, x1956);
  nand n2211(x2211, x1210, x1930);
  nand n2212(x2212, x2211, x2210);
  nand n2213(x2213, x70913, x2203);
  nand n2214(x2214, x1201, x2206);
  nand n2215(x2215, x2214, x2213);
  nand n2216(x2216, x70913, x2209);
  nand n2217(x2217, x1201, x2212);
  nand n2218(x2218, x2217, x2216);
  nand n2219(x2219, x70929, x2215);
  nand n2220(x2220, x1196, x2218);
  nand n2221(x2221, x2220, x2219);
  nand n2222(x2222, x70897, x2116);
  nand n2223(x2223, x1210, x2090);
  nand n2224(x2224, x2223, x2222);
  nand n2225(x2225, x70897, x2064);
  nand n2226(x2226, x1210, x2038);
  nand n2227(x2227, x2226, x2225);
  nand n2228(x2228, x70897, x2012);
  nand n2229(x2229, x1210, x1986);
  nand n2230(x2230, x2229, x2228);
  nand n2231(x2231, x70897, x1960);
  nand n2232(x2232, x1210, x1934);
  nand n2233(x2233, x2232, x2231);
  nand n2234(x2234, x70913, x2224);
  nand n2235(x2235, x1201, x2227);
  nand n2236(x2236, x2235, x2234);
  nand n2237(x2237, x70913, x2230);
  nand n2238(x2238, x1201, x2233);
  nand n2239(x2239, x2238, x2237);
  nand n2240(x2240, x70929, x2236);
  nand n2241(x2241, x1196, x2239);
  nand n2242(x2242, x2241, x2240);
  nand n2243(x2243, x1705, x1709);
  nand n2245(x2245, x2244, x1701);
  nand n2246(x2246, x1185, x1190);
  nand n2248(x2248, x2244, x2247);
  nand n2249(x2249, x1186, x1190);
  nand n2251(x2251, x1711, x2250);
  nand n2252(x2252, x2251, x2248);
  nand n2254(x2254, x2253, x2245);
  nand n2255(x2255, x2254, x71230);
  nand n2257(x2257, x2256, x71215);
  nand n2258(x2258, x2257, x2255);
  nand n2259(x2259, x2254, x71235);
  nand n2260(x2260, x2256, x71220);
  nand n2261(x2261, x2260, x2259);
  nand n2262(x2262, x2254, x71240);
  nand n2263(x2263, x2256, x71225);
  nand n2264(x2264, x2263, x2262);
  nand n2265(x2265, x2248, x2245);
  nand n2266(x2266, x2265, x71215);
  nand n2268(x2268, x2267, x71202);
  nand n2269(x2269, x2268, x2266);
  nand n2270(x2270, x2265, x71220);
  nand n2271(x2271, x2267, x71205);
  nand n2272(x2272, x2271, x2270);
  nand n2273(x2273, x2265, x71225);
  nand n2274(x2274, x2267, x71210);
  nand n2275(x2275, x2274, x2273);
  nand n2276(x2276, x71072, x71074);
  nand n2277(x2277, x71068, x71070);
  nand n2280(x2280, x2279, x2278);
  nand n2282(x2282, x2281, x2280);
  nand n2284(x2284, x70721, x2280);
  nand n2287(x2287, x2286, x2283);
  nand n2289(x2289, x70705, x2283);
  nand n2291(x2291, x2286, x2285);
  nand n2293(x2293, x70705, x2285);
  nand n2296(x2296, x2295, x2288);
  nand n2298(x2298, x70689, x2288);
  nand n2300(x2300, x2295, x2290);
  nand n2302(x2302, x70689, x2290);
  nand n2304(x2304, x2295, x2292);
  nand n2306(x2306, x70689, x2292);
  nand n2308(x2308, x2295, x2294);
  nand n2310(x2310, x70689, x2294);
  nand n2312(x2312, x2297, x71069);
  nand n2314(x2314, x2313, x68889);
  nand n2315(x2315, x2312, x2317);
  nand n2316(x2316, x2315, x2314);
  nand n2318(x2318, x2313, x68903);
  nand n2319(x2319, x2312, x2321);
  nand n2320(x2320, x2319, x2318);
  nand n2322(x2322, x2313, x68917);
  nand n2323(x2323, x2312, x2325);
  nand n2324(x2324, x2323, x2322);
  nand n2326(x2326, x2313, x68931);
  nand n2327(x2327, x2312, x2329);
  nand n2328(x2328, x2327, x2326);
  nand n2330(x2330, x2313, x68945);
  nand n2331(x2331, x2312, x2333);
  nand n2332(x2332, x2331, x2330);
  nand n2334(x2334, x2313, x68959);
  nand n2335(x2335, x2312, x2337);
  nand n2336(x2336, x2335, x2334);
  nand n2338(x2338, x2313, x68973);
  nand n2339(x2339, x2312, x2341);
  nand n2340(x2340, x2339, x2338);
  nand n2342(x2342, x2313, x68987);
  nand n2343(x2343, x2312, x2345);
  nand n2344(x2344, x2343, x2342);
  nand n2346(x2346, x2313, x69001);
  nand n2347(x2347, x2312, x2349);
  nand n2348(x2348, x2347, x2346);
  nand n2350(x2350, x2313, x69015);
  nand n2351(x2351, x2312, x2353);
  nand n2352(x2352, x2351, x2350);
  nand n2354(x2354, x2313, x69029);
  nand n2355(x2355, x2312, x2357);
  nand n2356(x2356, x2355, x2354);
  nand n2358(x2358, x2313, x69043);
  nand n2359(x2359, x2312, x2361);
  nand n2360(x2360, x2359, x2358);
  nand n2362(x2362, x2313, x69057);
  nand n2363(x2363, x2312, x2365);
  nand n2364(x2364, x2363, x2362);
  nand n2366(x2366, x2313, x69071);
  nand n2367(x2367, x2312, x2369);
  nand n2368(x2368, x2367, x2366);
  nand n2370(x2370, x2313, x69085);
  nand n2371(x2371, x2312, x2373);
  nand n2372(x2372, x2371, x2370);
  nand n2374(x2374, x2313, x69099);
  nand n2375(x2375, x2312, x2377);
  nand n2376(x2376, x2375, x2374);
  nand n2378(x2378, x2313, x69113);
  nand n2379(x2379, x2312, x2381);
  nand n2380(x2380, x2379, x2378);
  nand n2382(x2382, x2313, x69127);
  nand n2383(x2383, x2312, x2385);
  nand n2384(x2384, x2383, x2382);
  nand n2386(x2386, x2313, x69141);
  nand n2387(x2387, x2312, x2389);
  nand n2388(x2388, x2387, x2386);
  nand n2390(x2390, x2313, x69155);
  nand n2391(x2391, x2312, x2393);
  nand n2392(x2392, x2391, x2390);
  nand n2394(x2394, x2313, x69169);
  nand n2395(x2395, x2312, x2397);
  nand n2396(x2396, x2395, x2394);
  nand n2398(x2398, x2313, x69183);
  nand n2399(x2399, x2312, x2401);
  nand n2400(x2400, x2399, x2398);
  nand n2402(x2402, x2313, x69197);
  nand n2403(x2403, x2312, x2405);
  nand n2404(x2404, x2403, x2402);
  nand n2406(x2406, x2313, x69211);
  nand n2407(x2407, x2312, x2409);
  nand n2408(x2408, x2407, x2406);
  nand n2410(x2410, x2313, x69225);
  nand n2411(x2411, x2312, x2413);
  nand n2412(x2412, x2411, x2410);
  nand n2414(x2414, x2313, x69239);
  nand n2415(x2415, x2312, x2417);
  nand n2416(x2416, x2415, x2414);
  nand n2418(x2418, x2313, x69253);
  nand n2419(x2419, x2312, x2421);
  nand n2420(x2420, x2419, x2418);
  nand n2422(x2422, x2313, x69267);
  nand n2423(x2423, x2312, x2425);
  nand n2424(x2424, x2423, x2422);
  nand n2426(x2426, x2313, x69281);
  nand n2427(x2427, x2312, x2429);
  nand n2428(x2428, x2427, x2426);
  nand n2430(x2430, x2313, x69295);
  nand n2431(x2431, x2312, x2433);
  nand n2432(x2432, x2431, x2430);
  nand n2434(x2434, x2313, x69309);
  nand n2435(x2435, x2312, x2437);
  nand n2436(x2436, x2435, x2434);
  nand n2438(x2438, x2313, x69323);
  nand n2439(x2439, x2312, x2441);
  nand n2440(x2440, x2439, x2438);
  nand n2442(x2442, x2299, x71069);
  nand n2444(x2444, x2443, x68889);
  nand n2445(x2445, x2442, x2447);
  nand n2446(x2446, x2445, x2444);
  nand n2448(x2448, x2443, x68903);
  nand n2449(x2449, x2442, x2451);
  nand n2450(x2450, x2449, x2448);
  nand n2452(x2452, x2443, x68917);
  nand n2453(x2453, x2442, x2455);
  nand n2454(x2454, x2453, x2452);
  nand n2456(x2456, x2443, x68931);
  nand n2457(x2457, x2442, x2459);
  nand n2458(x2458, x2457, x2456);
  nand n2460(x2460, x2443, x68945);
  nand n2461(x2461, x2442, x2463);
  nand n2462(x2462, x2461, x2460);
  nand n2464(x2464, x2443, x68959);
  nand n2465(x2465, x2442, x2467);
  nand n2466(x2466, x2465, x2464);
  nand n2468(x2468, x2443, x68973);
  nand n2469(x2469, x2442, x2471);
  nand n2470(x2470, x2469, x2468);
  nand n2472(x2472, x2443, x68987);
  nand n2473(x2473, x2442, x2475);
  nand n2474(x2474, x2473, x2472);
  nand n2476(x2476, x2443, x69001);
  nand n2477(x2477, x2442, x2479);
  nand n2478(x2478, x2477, x2476);
  nand n2480(x2480, x2443, x69015);
  nand n2481(x2481, x2442, x2483);
  nand n2482(x2482, x2481, x2480);
  nand n2484(x2484, x2443, x69029);
  nand n2485(x2485, x2442, x2487);
  nand n2486(x2486, x2485, x2484);
  nand n2488(x2488, x2443, x69043);
  nand n2489(x2489, x2442, x2491);
  nand n2490(x2490, x2489, x2488);
  nand n2492(x2492, x2443, x69057);
  nand n2493(x2493, x2442, x2495);
  nand n2494(x2494, x2493, x2492);
  nand n2496(x2496, x2443, x69071);
  nand n2497(x2497, x2442, x2499);
  nand n2498(x2498, x2497, x2496);
  nand n2500(x2500, x2443, x69085);
  nand n2501(x2501, x2442, x2503);
  nand n2502(x2502, x2501, x2500);
  nand n2504(x2504, x2443, x69099);
  nand n2505(x2505, x2442, x2507);
  nand n2506(x2506, x2505, x2504);
  nand n2508(x2508, x2443, x69113);
  nand n2509(x2509, x2442, x2511);
  nand n2510(x2510, x2509, x2508);
  nand n2512(x2512, x2443, x69127);
  nand n2513(x2513, x2442, x2515);
  nand n2514(x2514, x2513, x2512);
  nand n2516(x2516, x2443, x69141);
  nand n2517(x2517, x2442, x2519);
  nand n2518(x2518, x2517, x2516);
  nand n2520(x2520, x2443, x69155);
  nand n2521(x2521, x2442, x2523);
  nand n2522(x2522, x2521, x2520);
  nand n2524(x2524, x2443, x69169);
  nand n2525(x2525, x2442, x2527);
  nand n2526(x2526, x2525, x2524);
  nand n2528(x2528, x2443, x69183);
  nand n2529(x2529, x2442, x2531);
  nand n2530(x2530, x2529, x2528);
  nand n2532(x2532, x2443, x69197);
  nand n2533(x2533, x2442, x2535);
  nand n2534(x2534, x2533, x2532);
  nand n2536(x2536, x2443, x69211);
  nand n2537(x2537, x2442, x2539);
  nand n2538(x2538, x2537, x2536);
  nand n2540(x2540, x2443, x69225);
  nand n2541(x2541, x2442, x2543);
  nand n2542(x2542, x2541, x2540);
  nand n2544(x2544, x2443, x69239);
  nand n2545(x2545, x2442, x2547);
  nand n2546(x2546, x2545, x2544);
  nand n2548(x2548, x2443, x69253);
  nand n2549(x2549, x2442, x2551);
  nand n2550(x2550, x2549, x2548);
  nand n2552(x2552, x2443, x69267);
  nand n2553(x2553, x2442, x2555);
  nand n2554(x2554, x2553, x2552);
  nand n2556(x2556, x2443, x69281);
  nand n2557(x2557, x2442, x2559);
  nand n2558(x2558, x2557, x2556);
  nand n2560(x2560, x2443, x69295);
  nand n2561(x2561, x2442, x2563);
  nand n2562(x2562, x2561, x2560);
  nand n2564(x2564, x2443, x69309);
  nand n2565(x2565, x2442, x2567);
  nand n2566(x2566, x2565, x2564);
  nand n2568(x2568, x2443, x69323);
  nand n2569(x2569, x2442, x2571);
  nand n2570(x2570, x2569, x2568);
  nand n2572(x2572, x2301, x71069);
  nand n2574(x2574, x2573, x68889);
  nand n2575(x2575, x2572, x2577);
  nand n2576(x2576, x2575, x2574);
  nand n2578(x2578, x2573, x68903);
  nand n2579(x2579, x2572, x2581);
  nand n2580(x2580, x2579, x2578);
  nand n2582(x2582, x2573, x68917);
  nand n2583(x2583, x2572, x2585);
  nand n2584(x2584, x2583, x2582);
  nand n2586(x2586, x2573, x68931);
  nand n2587(x2587, x2572, x2589);
  nand n2588(x2588, x2587, x2586);
  nand n2590(x2590, x2573, x68945);
  nand n2591(x2591, x2572, x2593);
  nand n2592(x2592, x2591, x2590);
  nand n2594(x2594, x2573, x68959);
  nand n2595(x2595, x2572, x2597);
  nand n2596(x2596, x2595, x2594);
  nand n2598(x2598, x2573, x68973);
  nand n2599(x2599, x2572, x2601);
  nand n2600(x2600, x2599, x2598);
  nand n2602(x2602, x2573, x68987);
  nand n2603(x2603, x2572, x2605);
  nand n2604(x2604, x2603, x2602);
  nand n2606(x2606, x2573, x69001);
  nand n2607(x2607, x2572, x2609);
  nand n2608(x2608, x2607, x2606);
  nand n2610(x2610, x2573, x69015);
  nand n2611(x2611, x2572, x2613);
  nand n2612(x2612, x2611, x2610);
  nand n2614(x2614, x2573, x69029);
  nand n2615(x2615, x2572, x2617);
  nand n2616(x2616, x2615, x2614);
  nand n2618(x2618, x2573, x69043);
  nand n2619(x2619, x2572, x2621);
  nand n2620(x2620, x2619, x2618);
  nand n2622(x2622, x2573, x69057);
  nand n2623(x2623, x2572, x2625);
  nand n2624(x2624, x2623, x2622);
  nand n2626(x2626, x2573, x69071);
  nand n2627(x2627, x2572, x2629);
  nand n2628(x2628, x2627, x2626);
  nand n2630(x2630, x2573, x69085);
  nand n2631(x2631, x2572, x2633);
  nand n2632(x2632, x2631, x2630);
  nand n2634(x2634, x2573, x69099);
  nand n2635(x2635, x2572, x2637);
  nand n2636(x2636, x2635, x2634);
  nand n2638(x2638, x2573, x69113);
  nand n2639(x2639, x2572, x2641);
  nand n2640(x2640, x2639, x2638);
  nand n2642(x2642, x2573, x69127);
  nand n2643(x2643, x2572, x2645);
  nand n2644(x2644, x2643, x2642);
  nand n2646(x2646, x2573, x69141);
  nand n2647(x2647, x2572, x2649);
  nand n2648(x2648, x2647, x2646);
  nand n2650(x2650, x2573, x69155);
  nand n2651(x2651, x2572, x2653);
  nand n2652(x2652, x2651, x2650);
  nand n2654(x2654, x2573, x69169);
  nand n2655(x2655, x2572, x2657);
  nand n2656(x2656, x2655, x2654);
  nand n2658(x2658, x2573, x69183);
  nand n2659(x2659, x2572, x2661);
  nand n2660(x2660, x2659, x2658);
  nand n2662(x2662, x2573, x69197);
  nand n2663(x2663, x2572, x2665);
  nand n2664(x2664, x2663, x2662);
  nand n2666(x2666, x2573, x69211);
  nand n2667(x2667, x2572, x2669);
  nand n2668(x2668, x2667, x2666);
  nand n2670(x2670, x2573, x69225);
  nand n2671(x2671, x2572, x2673);
  nand n2672(x2672, x2671, x2670);
  nand n2674(x2674, x2573, x69239);
  nand n2675(x2675, x2572, x2677);
  nand n2676(x2676, x2675, x2674);
  nand n2678(x2678, x2573, x69253);
  nand n2679(x2679, x2572, x2681);
  nand n2680(x2680, x2679, x2678);
  nand n2682(x2682, x2573, x69267);
  nand n2683(x2683, x2572, x2685);
  nand n2684(x2684, x2683, x2682);
  nand n2686(x2686, x2573, x69281);
  nand n2687(x2687, x2572, x2689);
  nand n2688(x2688, x2687, x2686);
  nand n2690(x2690, x2573, x69295);
  nand n2691(x2691, x2572, x2693);
  nand n2692(x2692, x2691, x2690);
  nand n2694(x2694, x2573, x69309);
  nand n2695(x2695, x2572, x2697);
  nand n2696(x2696, x2695, x2694);
  nand n2698(x2698, x2573, x69323);
  nand n2699(x2699, x2572, x2701);
  nand n2700(x2700, x2699, x2698);
  nand n2702(x2702, x2303, x71069);
  nand n2704(x2704, x2703, x68889);
  nand n2705(x2705, x2702, x2707);
  nand n2706(x2706, x2705, x2704);
  nand n2708(x2708, x2703, x68903);
  nand n2709(x2709, x2702, x2711);
  nand n2710(x2710, x2709, x2708);
  nand n2712(x2712, x2703, x68917);
  nand n2713(x2713, x2702, x2715);
  nand n2714(x2714, x2713, x2712);
  nand n2716(x2716, x2703, x68931);
  nand n2717(x2717, x2702, x2719);
  nand n2718(x2718, x2717, x2716);
  nand n2720(x2720, x2703, x68945);
  nand n2721(x2721, x2702, x2723);
  nand n2722(x2722, x2721, x2720);
  nand n2724(x2724, x2703, x68959);
  nand n2725(x2725, x2702, x2727);
  nand n2726(x2726, x2725, x2724);
  nand n2728(x2728, x2703, x68973);
  nand n2729(x2729, x2702, x2731);
  nand n2730(x2730, x2729, x2728);
  nand n2732(x2732, x2703, x68987);
  nand n2733(x2733, x2702, x2735);
  nand n2734(x2734, x2733, x2732);
  nand n2736(x2736, x2703, x69001);
  nand n2737(x2737, x2702, x2739);
  nand n2738(x2738, x2737, x2736);
  nand n2740(x2740, x2703, x69015);
  nand n2741(x2741, x2702, x2743);
  nand n2742(x2742, x2741, x2740);
  nand n2744(x2744, x2703, x69029);
  nand n2745(x2745, x2702, x2747);
  nand n2746(x2746, x2745, x2744);
  nand n2748(x2748, x2703, x69043);
  nand n2749(x2749, x2702, x2751);
  nand n2750(x2750, x2749, x2748);
  nand n2752(x2752, x2703, x69057);
  nand n2753(x2753, x2702, x2755);
  nand n2754(x2754, x2753, x2752);
  nand n2756(x2756, x2703, x69071);
  nand n2757(x2757, x2702, x2759);
  nand n2758(x2758, x2757, x2756);
  nand n2760(x2760, x2703, x69085);
  nand n2761(x2761, x2702, x2763);
  nand n2762(x2762, x2761, x2760);
  nand n2764(x2764, x2703, x69099);
  nand n2765(x2765, x2702, x2767);
  nand n2766(x2766, x2765, x2764);
  nand n2768(x2768, x2703, x69113);
  nand n2769(x2769, x2702, x2771);
  nand n2770(x2770, x2769, x2768);
  nand n2772(x2772, x2703, x69127);
  nand n2773(x2773, x2702, x2775);
  nand n2774(x2774, x2773, x2772);
  nand n2776(x2776, x2703, x69141);
  nand n2777(x2777, x2702, x2779);
  nand n2778(x2778, x2777, x2776);
  nand n2780(x2780, x2703, x69155);
  nand n2781(x2781, x2702, x2783);
  nand n2782(x2782, x2781, x2780);
  nand n2784(x2784, x2703, x69169);
  nand n2785(x2785, x2702, x2787);
  nand n2786(x2786, x2785, x2784);
  nand n2788(x2788, x2703, x69183);
  nand n2789(x2789, x2702, x2791);
  nand n2790(x2790, x2789, x2788);
  nand n2792(x2792, x2703, x69197);
  nand n2793(x2793, x2702, x2795);
  nand n2794(x2794, x2793, x2792);
  nand n2796(x2796, x2703, x69211);
  nand n2797(x2797, x2702, x2799);
  nand n2798(x2798, x2797, x2796);
  nand n2800(x2800, x2703, x69225);
  nand n2801(x2801, x2702, x2803);
  nand n2802(x2802, x2801, x2800);
  nand n2804(x2804, x2703, x69239);
  nand n2805(x2805, x2702, x2807);
  nand n2806(x2806, x2805, x2804);
  nand n2808(x2808, x2703, x69253);
  nand n2809(x2809, x2702, x2811);
  nand n2810(x2810, x2809, x2808);
  nand n2812(x2812, x2703, x69267);
  nand n2813(x2813, x2702, x2815);
  nand n2814(x2814, x2813, x2812);
  nand n2816(x2816, x2703, x69281);
  nand n2817(x2817, x2702, x2819);
  nand n2818(x2818, x2817, x2816);
  nand n2820(x2820, x2703, x69295);
  nand n2821(x2821, x2702, x2823);
  nand n2822(x2822, x2821, x2820);
  nand n2824(x2824, x2703, x69309);
  nand n2825(x2825, x2702, x2827);
  nand n2826(x2826, x2825, x2824);
  nand n2828(x2828, x2703, x69323);
  nand n2829(x2829, x2702, x2831);
  nand n2830(x2830, x2829, x2828);
  nand n2832(x2832, x2305, x71069);
  nand n2834(x2834, x2833, x68889);
  nand n2835(x2835, x2832, x2837);
  nand n2836(x2836, x2835, x2834);
  nand n2838(x2838, x2833, x68903);
  nand n2839(x2839, x2832, x2841);
  nand n2840(x2840, x2839, x2838);
  nand n2842(x2842, x2833, x68917);
  nand n2843(x2843, x2832, x2845);
  nand n2844(x2844, x2843, x2842);
  nand n2846(x2846, x2833, x68931);
  nand n2847(x2847, x2832, x2849);
  nand n2848(x2848, x2847, x2846);
  nand n2850(x2850, x2833, x68945);
  nand n2851(x2851, x2832, x2853);
  nand n2852(x2852, x2851, x2850);
  nand n2854(x2854, x2833, x68959);
  nand n2855(x2855, x2832, x2857);
  nand n2856(x2856, x2855, x2854);
  nand n2858(x2858, x2833, x68973);
  nand n2859(x2859, x2832, x2861);
  nand n2860(x2860, x2859, x2858);
  nand n2862(x2862, x2833, x68987);
  nand n2863(x2863, x2832, x2865);
  nand n2864(x2864, x2863, x2862);
  nand n2866(x2866, x2833, x69001);
  nand n2867(x2867, x2832, x2869);
  nand n2868(x2868, x2867, x2866);
  nand n2870(x2870, x2833, x69015);
  nand n2871(x2871, x2832, x2873);
  nand n2872(x2872, x2871, x2870);
  nand n2874(x2874, x2833, x69029);
  nand n2875(x2875, x2832, x2877);
  nand n2876(x2876, x2875, x2874);
  nand n2878(x2878, x2833, x69043);
  nand n2879(x2879, x2832, x2881);
  nand n2880(x2880, x2879, x2878);
  nand n2882(x2882, x2833, x69057);
  nand n2883(x2883, x2832, x2885);
  nand n2884(x2884, x2883, x2882);
  nand n2886(x2886, x2833, x69071);
  nand n2887(x2887, x2832, x2889);
  nand n2888(x2888, x2887, x2886);
  nand n2890(x2890, x2833, x69085);
  nand n2891(x2891, x2832, x2893);
  nand n2892(x2892, x2891, x2890);
  nand n2894(x2894, x2833, x69099);
  nand n2895(x2895, x2832, x2897);
  nand n2896(x2896, x2895, x2894);
  nand n2898(x2898, x2833, x69113);
  nand n2899(x2899, x2832, x2901);
  nand n2900(x2900, x2899, x2898);
  nand n2902(x2902, x2833, x69127);
  nand n2903(x2903, x2832, x2905);
  nand n2904(x2904, x2903, x2902);
  nand n2906(x2906, x2833, x69141);
  nand n2907(x2907, x2832, x2909);
  nand n2908(x2908, x2907, x2906);
  nand n2910(x2910, x2833, x69155);
  nand n2911(x2911, x2832, x2913);
  nand n2912(x2912, x2911, x2910);
  nand n2914(x2914, x2833, x69169);
  nand n2915(x2915, x2832, x2917);
  nand n2916(x2916, x2915, x2914);
  nand n2918(x2918, x2833, x69183);
  nand n2919(x2919, x2832, x2921);
  nand n2920(x2920, x2919, x2918);
  nand n2922(x2922, x2833, x69197);
  nand n2923(x2923, x2832, x2925);
  nand n2924(x2924, x2923, x2922);
  nand n2926(x2926, x2833, x69211);
  nand n2927(x2927, x2832, x2929);
  nand n2928(x2928, x2927, x2926);
  nand n2930(x2930, x2833, x69225);
  nand n2931(x2931, x2832, x2933);
  nand n2932(x2932, x2931, x2930);
  nand n2934(x2934, x2833, x69239);
  nand n2935(x2935, x2832, x2937);
  nand n2936(x2936, x2935, x2934);
  nand n2938(x2938, x2833, x69253);
  nand n2939(x2939, x2832, x2941);
  nand n2940(x2940, x2939, x2938);
  nand n2942(x2942, x2833, x69267);
  nand n2943(x2943, x2832, x2945);
  nand n2944(x2944, x2943, x2942);
  nand n2946(x2946, x2833, x69281);
  nand n2947(x2947, x2832, x2949);
  nand n2948(x2948, x2947, x2946);
  nand n2950(x2950, x2833, x69295);
  nand n2951(x2951, x2832, x2953);
  nand n2952(x2952, x2951, x2950);
  nand n2954(x2954, x2833, x69309);
  nand n2955(x2955, x2832, x2957);
  nand n2956(x2956, x2955, x2954);
  nand n2958(x2958, x2833, x69323);
  nand n2959(x2959, x2832, x2961);
  nand n2960(x2960, x2959, x2958);
  nand n2962(x2962, x2307, x71069);
  nand n2964(x2964, x2963, x68889);
  nand n2965(x2965, x2962, x2967);
  nand n2966(x2966, x2965, x2964);
  nand n2968(x2968, x2963, x68903);
  nand n2969(x2969, x2962, x2971);
  nand n2970(x2970, x2969, x2968);
  nand n2972(x2972, x2963, x68917);
  nand n2973(x2973, x2962, x2975);
  nand n2974(x2974, x2973, x2972);
  nand n2976(x2976, x2963, x68931);
  nand n2977(x2977, x2962, x2979);
  nand n2978(x2978, x2977, x2976);
  nand n2980(x2980, x2963, x68945);
  nand n2981(x2981, x2962, x2983);
  nand n2982(x2982, x2981, x2980);
  nand n2984(x2984, x2963, x68959);
  nand n2985(x2985, x2962, x2987);
  nand n2986(x2986, x2985, x2984);
  nand n2988(x2988, x2963, x68973);
  nand n2989(x2989, x2962, x2991);
  nand n2990(x2990, x2989, x2988);
  nand n2992(x2992, x2963, x68987);
  nand n2993(x2993, x2962, x2995);
  nand n2994(x2994, x2993, x2992);
  nand n2996(x2996, x2963, x69001);
  nand n2997(x2997, x2962, x2999);
  nand n2998(x2998, x2997, x2996);
  nand n3000(x3000, x2963, x69015);
  nand n3001(x3001, x2962, x3003);
  nand n3002(x3002, x3001, x3000);
  nand n3004(x3004, x2963, x69029);
  nand n3005(x3005, x2962, x3007);
  nand n3006(x3006, x3005, x3004);
  nand n3008(x3008, x2963, x69043);
  nand n3009(x3009, x2962, x3011);
  nand n3010(x3010, x3009, x3008);
  nand n3012(x3012, x2963, x69057);
  nand n3013(x3013, x2962, x3015);
  nand n3014(x3014, x3013, x3012);
  nand n3016(x3016, x2963, x69071);
  nand n3017(x3017, x2962, x3019);
  nand n3018(x3018, x3017, x3016);
  nand n3020(x3020, x2963, x69085);
  nand n3021(x3021, x2962, x3023);
  nand n3022(x3022, x3021, x3020);
  nand n3024(x3024, x2963, x69099);
  nand n3025(x3025, x2962, x3027);
  nand n3026(x3026, x3025, x3024);
  nand n3028(x3028, x2963, x69113);
  nand n3029(x3029, x2962, x3031);
  nand n3030(x3030, x3029, x3028);
  nand n3032(x3032, x2963, x69127);
  nand n3033(x3033, x2962, x3035);
  nand n3034(x3034, x3033, x3032);
  nand n3036(x3036, x2963, x69141);
  nand n3037(x3037, x2962, x3039);
  nand n3038(x3038, x3037, x3036);
  nand n3040(x3040, x2963, x69155);
  nand n3041(x3041, x2962, x3043);
  nand n3042(x3042, x3041, x3040);
  nand n3044(x3044, x2963, x69169);
  nand n3045(x3045, x2962, x3047);
  nand n3046(x3046, x3045, x3044);
  nand n3048(x3048, x2963, x69183);
  nand n3049(x3049, x2962, x3051);
  nand n3050(x3050, x3049, x3048);
  nand n3052(x3052, x2963, x69197);
  nand n3053(x3053, x2962, x3055);
  nand n3054(x3054, x3053, x3052);
  nand n3056(x3056, x2963, x69211);
  nand n3057(x3057, x2962, x3059);
  nand n3058(x3058, x3057, x3056);
  nand n3060(x3060, x2963, x69225);
  nand n3061(x3061, x2962, x3063);
  nand n3062(x3062, x3061, x3060);
  nand n3064(x3064, x2963, x69239);
  nand n3065(x3065, x2962, x3067);
  nand n3066(x3066, x3065, x3064);
  nand n3068(x3068, x2963, x69253);
  nand n3069(x3069, x2962, x3071);
  nand n3070(x3070, x3069, x3068);
  nand n3072(x3072, x2963, x69267);
  nand n3073(x3073, x2962, x3075);
  nand n3074(x3074, x3073, x3072);
  nand n3076(x3076, x2963, x69281);
  nand n3077(x3077, x2962, x3079);
  nand n3078(x3078, x3077, x3076);
  nand n3080(x3080, x2963, x69295);
  nand n3081(x3081, x2962, x3083);
  nand n3082(x3082, x3081, x3080);
  nand n3084(x3084, x2963, x69309);
  nand n3085(x3085, x2962, x3087);
  nand n3086(x3086, x3085, x3084);
  nand n3088(x3088, x2963, x69323);
  nand n3089(x3089, x2962, x3091);
  nand n3090(x3090, x3089, x3088);
  nand n3092(x3092, x2309, x71069);
  nand n3094(x3094, x3093, x68889);
  nand n3095(x3095, x3092, x3097);
  nand n3096(x3096, x3095, x3094);
  nand n3098(x3098, x3093, x68903);
  nand n3099(x3099, x3092, x3101);
  nand n3100(x3100, x3099, x3098);
  nand n3102(x3102, x3093, x68917);
  nand n3103(x3103, x3092, x3105);
  nand n3104(x3104, x3103, x3102);
  nand n3106(x3106, x3093, x68931);
  nand n3107(x3107, x3092, x3109);
  nand n3108(x3108, x3107, x3106);
  nand n3110(x3110, x3093, x68945);
  nand n3111(x3111, x3092, x3113);
  nand n3112(x3112, x3111, x3110);
  nand n3114(x3114, x3093, x68959);
  nand n3115(x3115, x3092, x3117);
  nand n3116(x3116, x3115, x3114);
  nand n3118(x3118, x3093, x68973);
  nand n3119(x3119, x3092, x3121);
  nand n3120(x3120, x3119, x3118);
  nand n3122(x3122, x3093, x68987);
  nand n3123(x3123, x3092, x3125);
  nand n3124(x3124, x3123, x3122);
  nand n3126(x3126, x3093, x69001);
  nand n3127(x3127, x3092, x3129);
  nand n3128(x3128, x3127, x3126);
  nand n3130(x3130, x3093, x69015);
  nand n3131(x3131, x3092, x3133);
  nand n3132(x3132, x3131, x3130);
  nand n3134(x3134, x3093, x69029);
  nand n3135(x3135, x3092, x3137);
  nand n3136(x3136, x3135, x3134);
  nand n3138(x3138, x3093, x69043);
  nand n3139(x3139, x3092, x3141);
  nand n3140(x3140, x3139, x3138);
  nand n3142(x3142, x3093, x69057);
  nand n3143(x3143, x3092, x3145);
  nand n3144(x3144, x3143, x3142);
  nand n3146(x3146, x3093, x69071);
  nand n3147(x3147, x3092, x3149);
  nand n3148(x3148, x3147, x3146);
  nand n3150(x3150, x3093, x69085);
  nand n3151(x3151, x3092, x3153);
  nand n3152(x3152, x3151, x3150);
  nand n3154(x3154, x3093, x69099);
  nand n3155(x3155, x3092, x3157);
  nand n3156(x3156, x3155, x3154);
  nand n3158(x3158, x3093, x69113);
  nand n3159(x3159, x3092, x3161);
  nand n3160(x3160, x3159, x3158);
  nand n3162(x3162, x3093, x69127);
  nand n3163(x3163, x3092, x3165);
  nand n3164(x3164, x3163, x3162);
  nand n3166(x3166, x3093, x69141);
  nand n3167(x3167, x3092, x3169);
  nand n3168(x3168, x3167, x3166);
  nand n3170(x3170, x3093, x69155);
  nand n3171(x3171, x3092, x3173);
  nand n3172(x3172, x3171, x3170);
  nand n3174(x3174, x3093, x69169);
  nand n3175(x3175, x3092, x3177);
  nand n3176(x3176, x3175, x3174);
  nand n3178(x3178, x3093, x69183);
  nand n3179(x3179, x3092, x3181);
  nand n3180(x3180, x3179, x3178);
  nand n3182(x3182, x3093, x69197);
  nand n3183(x3183, x3092, x3185);
  nand n3184(x3184, x3183, x3182);
  nand n3186(x3186, x3093, x69211);
  nand n3187(x3187, x3092, x3189);
  nand n3188(x3188, x3187, x3186);
  nand n3190(x3190, x3093, x69225);
  nand n3191(x3191, x3092, x3193);
  nand n3192(x3192, x3191, x3190);
  nand n3194(x3194, x3093, x69239);
  nand n3195(x3195, x3092, x3197);
  nand n3196(x3196, x3195, x3194);
  nand n3198(x3198, x3093, x69253);
  nand n3199(x3199, x3092, x3201);
  nand n3200(x3200, x3199, x3198);
  nand n3202(x3202, x3093, x69267);
  nand n3203(x3203, x3092, x3205);
  nand n3204(x3204, x3203, x3202);
  nand n3206(x3206, x3093, x69281);
  nand n3207(x3207, x3092, x3209);
  nand n3208(x3208, x3207, x3206);
  nand n3210(x3210, x3093, x69295);
  nand n3211(x3211, x3092, x3213);
  nand n3212(x3212, x3211, x3210);
  nand n3214(x3214, x3093, x69309);
  nand n3215(x3215, x3092, x3217);
  nand n3216(x3216, x3215, x3214);
  nand n3218(x3218, x3093, x69323);
  nand n3219(x3219, x3092, x3221);
  nand n3220(x3220, x3219, x3218);
  nand n3222(x3222, x2311, x71069);
  nand n3224(x3224, x3223, x68889);
  nand n3225(x3225, x3222, x3227);
  nand n3226(x3226, x3225, x3224);
  nand n3228(x3228, x3223, x68903);
  nand n3229(x3229, x3222, x3231);
  nand n3230(x3230, x3229, x3228);
  nand n3232(x3232, x3223, x68917);
  nand n3233(x3233, x3222, x3235);
  nand n3234(x3234, x3233, x3232);
  nand n3236(x3236, x3223, x68931);
  nand n3237(x3237, x3222, x3239);
  nand n3238(x3238, x3237, x3236);
  nand n3240(x3240, x3223, x68945);
  nand n3241(x3241, x3222, x3243);
  nand n3242(x3242, x3241, x3240);
  nand n3244(x3244, x3223, x68959);
  nand n3245(x3245, x3222, x3247);
  nand n3246(x3246, x3245, x3244);
  nand n3248(x3248, x3223, x68973);
  nand n3249(x3249, x3222, x3251);
  nand n3250(x3250, x3249, x3248);
  nand n3252(x3252, x3223, x68987);
  nand n3253(x3253, x3222, x3255);
  nand n3254(x3254, x3253, x3252);
  nand n3256(x3256, x3223, x69001);
  nand n3257(x3257, x3222, x3259);
  nand n3258(x3258, x3257, x3256);
  nand n3260(x3260, x3223, x69015);
  nand n3261(x3261, x3222, x3263);
  nand n3262(x3262, x3261, x3260);
  nand n3264(x3264, x3223, x69029);
  nand n3265(x3265, x3222, x3267);
  nand n3266(x3266, x3265, x3264);
  nand n3268(x3268, x3223, x69043);
  nand n3269(x3269, x3222, x3271);
  nand n3270(x3270, x3269, x3268);
  nand n3272(x3272, x3223, x69057);
  nand n3273(x3273, x3222, x3275);
  nand n3274(x3274, x3273, x3272);
  nand n3276(x3276, x3223, x69071);
  nand n3277(x3277, x3222, x3279);
  nand n3278(x3278, x3277, x3276);
  nand n3280(x3280, x3223, x69085);
  nand n3281(x3281, x3222, x3283);
  nand n3282(x3282, x3281, x3280);
  nand n3284(x3284, x3223, x69099);
  nand n3285(x3285, x3222, x3287);
  nand n3286(x3286, x3285, x3284);
  nand n3288(x3288, x3223, x69113);
  nand n3289(x3289, x3222, x3291);
  nand n3290(x3290, x3289, x3288);
  nand n3292(x3292, x3223, x69127);
  nand n3293(x3293, x3222, x3295);
  nand n3294(x3294, x3293, x3292);
  nand n3296(x3296, x3223, x69141);
  nand n3297(x3297, x3222, x3299);
  nand n3298(x3298, x3297, x3296);
  nand n3300(x3300, x3223, x69155);
  nand n3301(x3301, x3222, x3303);
  nand n3302(x3302, x3301, x3300);
  nand n3304(x3304, x3223, x69169);
  nand n3305(x3305, x3222, x3307);
  nand n3306(x3306, x3305, x3304);
  nand n3308(x3308, x3223, x69183);
  nand n3309(x3309, x3222, x3311);
  nand n3310(x3310, x3309, x3308);
  nand n3312(x3312, x3223, x69197);
  nand n3313(x3313, x3222, x3315);
  nand n3314(x3314, x3313, x3312);
  nand n3316(x3316, x3223, x69211);
  nand n3317(x3317, x3222, x3319);
  nand n3318(x3318, x3317, x3316);
  nand n3320(x3320, x3223, x69225);
  nand n3321(x3321, x3222, x3323);
  nand n3322(x3322, x3321, x3320);
  nand n3324(x3324, x3223, x69239);
  nand n3325(x3325, x3222, x3327);
  nand n3326(x3326, x3325, x3324);
  nand n3328(x3328, x3223, x69253);
  nand n3329(x3329, x3222, x3331);
  nand n3330(x3330, x3329, x3328);
  nand n3332(x3332, x3223, x69267);
  nand n3333(x3333, x3222, x3335);
  nand n3334(x3334, x3333, x3332);
  nand n3336(x3336, x3223, x69281);
  nand n3337(x3337, x3222, x3339);
  nand n3338(x3338, x3337, x3336);
  nand n3340(x3340, x3223, x69295);
  nand n3341(x3341, x3222, x3343);
  nand n3342(x3342, x3341, x3340);
  nand n3344(x3344, x3223, x69309);
  nand n3345(x3345, x3222, x3347);
  nand n3346(x3346, x3345, x3344);
  nand n3348(x3348, x3223, x69323);
  nand n3349(x3349, x3222, x3351);
  nand n3350(x3350, x3349, x3348);
  nand n3352(x3352, x2297, x71071);
  nand n3354(x3354, x3353, x69339);
  nand n3355(x3355, x3352, x3359);
  nand n3356(x3356, x3355, x3354);
  nand n3360(x3360, x3353, x69353);
  nand n3361(x3361, x3352, x3363);
  nand n3362(x3362, x3361, x3360);
  nand n3364(x3364, x3353, x69367);
  nand n3365(x3365, x3352, x3367);
  nand n3366(x3366, x3365, x3364);
  nand n3368(x3368, x3353, x69381);
  nand n3369(x3369, x3352, x3371);
  nand n3370(x3370, x3369, x3368);
  nand n3372(x3372, x3353, x69395);
  nand n3373(x3373, x3352, x3375);
  nand n3374(x3374, x3373, x3372);
  nand n3376(x3376, x3353, x69409);
  nand n3377(x3377, x3352, x3379);
  nand n3378(x3378, x3377, x3376);
  nand n3380(x3380, x3353, x69423);
  nand n3381(x3381, x3352, x3383);
  nand n3382(x3382, x3381, x3380);
  nand n3384(x3384, x3353, x69437);
  nand n3385(x3385, x3352, x3387);
  nand n3386(x3386, x3385, x3384);
  nand n3388(x3388, x3353, x69451);
  nand n3389(x3389, x3352, x3391);
  nand n3390(x3390, x3389, x3388);
  nand n3392(x3392, x3353, x69465);
  nand n3393(x3393, x3352, x3395);
  nand n3394(x3394, x3393, x3392);
  nand n3396(x3396, x3353, x69479);
  nand n3397(x3397, x3352, x3399);
  nand n3398(x3398, x3397, x3396);
  nand n3400(x3400, x3353, x69493);
  nand n3401(x3401, x3352, x3403);
  nand n3402(x3402, x3401, x3400);
  nand n3404(x3404, x3353, x69507);
  nand n3405(x3405, x3352, x3407);
  nand n3406(x3406, x3405, x3404);
  nand n3408(x3408, x3353, x69521);
  nand n3409(x3409, x3352, x3411);
  nand n3410(x3410, x3409, x3408);
  nand n3412(x3412, x3353, x69535);
  nand n3413(x3413, x3352, x3415);
  nand n3414(x3414, x3413, x3412);
  nand n3416(x3416, x3353, x69549);
  nand n3417(x3417, x3352, x3419);
  nand n3418(x3418, x3417, x3416);
  nand n3420(x3420, x3353, x69563);
  nand n3421(x3421, x3352, x3423);
  nand n3422(x3422, x3421, x3420);
  nand n3424(x3424, x3353, x69577);
  nand n3425(x3425, x3352, x3427);
  nand n3426(x3426, x3425, x3424);
  nand n3428(x3428, x3353, x69591);
  nand n3429(x3429, x3352, x3431);
  nand n3430(x3430, x3429, x3428);
  nand n3432(x3432, x3353, x69605);
  nand n3433(x3433, x3352, x3435);
  nand n3434(x3434, x3433, x3432);
  nand n3436(x3436, x3353, x69619);
  nand n3437(x3437, x3352, x3439);
  nand n3438(x3438, x3437, x3436);
  nand n3440(x3440, x3353, x69633);
  nand n3441(x3441, x3352, x3443);
  nand n3442(x3442, x3441, x3440);
  nand n3444(x3444, x3353, x69647);
  nand n3445(x3445, x3352, x3447);
  nand n3446(x3446, x3445, x3444);
  nand n3448(x3448, x3353, x69661);
  nand n3449(x3449, x3352, x3451);
  nand n3450(x3450, x3449, x3448);
  nand n3452(x3452, x3353, x69675);
  nand n3453(x3453, x3352, x3455);
  nand n3454(x3454, x3453, x3452);
  nand n3456(x3456, x3353, x69689);
  nand n3457(x3457, x3352, x3459);
  nand n3458(x3458, x3457, x3456);
  nand n3460(x3460, x3353, x69703);
  nand n3461(x3461, x3352, x3463);
  nand n3462(x3462, x3461, x3460);
  nand n3464(x3464, x3353, x69717);
  nand n3465(x3465, x3352, x3467);
  nand n3466(x3466, x3465, x3464);
  nand n3468(x3468, x3353, x69731);
  nand n3469(x3469, x3352, x3471);
  nand n3470(x3470, x3469, x3468);
  nand n3472(x3472, x3353, x69745);
  nand n3473(x3473, x3352, x3475);
  nand n3474(x3474, x3473, x3472);
  nand n3476(x3476, x3353, x69759);
  nand n3477(x3477, x3352, x3479);
  nand n3478(x3478, x3477, x3476);
  nand n3480(x3480, x3353, x69773);
  nand n3481(x3481, x3352, x3483);
  nand n3482(x3482, x3481, x3480);
  nand n3484(x3484, x2299, x71071);
  nand n3486(x3486, x3485, x69339);
  nand n3487(x3487, x3484, x3489);
  nand n3488(x3488, x3487, x3486);
  nand n3490(x3490, x3485, x69353);
  nand n3491(x3491, x3484, x3493);
  nand n3492(x3492, x3491, x3490);
  nand n3494(x3494, x3485, x69367);
  nand n3495(x3495, x3484, x3497);
  nand n3496(x3496, x3495, x3494);
  nand n3498(x3498, x3485, x69381);
  nand n3499(x3499, x3484, x3501);
  nand n3500(x3500, x3499, x3498);
  nand n3502(x3502, x3485, x69395);
  nand n3503(x3503, x3484, x3505);
  nand n3504(x3504, x3503, x3502);
  nand n3506(x3506, x3485, x69409);
  nand n3507(x3507, x3484, x3509);
  nand n3508(x3508, x3507, x3506);
  nand n3510(x3510, x3485, x69423);
  nand n3511(x3511, x3484, x3513);
  nand n3512(x3512, x3511, x3510);
  nand n3514(x3514, x3485, x69437);
  nand n3515(x3515, x3484, x3517);
  nand n3516(x3516, x3515, x3514);
  nand n3518(x3518, x3485, x69451);
  nand n3519(x3519, x3484, x3521);
  nand n3520(x3520, x3519, x3518);
  nand n3522(x3522, x3485, x69465);
  nand n3523(x3523, x3484, x3525);
  nand n3524(x3524, x3523, x3522);
  nand n3526(x3526, x3485, x69479);
  nand n3527(x3527, x3484, x3529);
  nand n3528(x3528, x3527, x3526);
  nand n3530(x3530, x3485, x69493);
  nand n3531(x3531, x3484, x3533);
  nand n3532(x3532, x3531, x3530);
  nand n3534(x3534, x3485, x69507);
  nand n3535(x3535, x3484, x3537);
  nand n3536(x3536, x3535, x3534);
  nand n3538(x3538, x3485, x69521);
  nand n3539(x3539, x3484, x3541);
  nand n3540(x3540, x3539, x3538);
  nand n3542(x3542, x3485, x69535);
  nand n3543(x3543, x3484, x3545);
  nand n3544(x3544, x3543, x3542);
  nand n3546(x3546, x3485, x69549);
  nand n3547(x3547, x3484, x3549);
  nand n3548(x3548, x3547, x3546);
  nand n3550(x3550, x3485, x69563);
  nand n3551(x3551, x3484, x3553);
  nand n3552(x3552, x3551, x3550);
  nand n3554(x3554, x3485, x69577);
  nand n3555(x3555, x3484, x3557);
  nand n3556(x3556, x3555, x3554);
  nand n3558(x3558, x3485, x69591);
  nand n3559(x3559, x3484, x3561);
  nand n3560(x3560, x3559, x3558);
  nand n3562(x3562, x3485, x69605);
  nand n3563(x3563, x3484, x3565);
  nand n3564(x3564, x3563, x3562);
  nand n3566(x3566, x3485, x69619);
  nand n3567(x3567, x3484, x3569);
  nand n3568(x3568, x3567, x3566);
  nand n3570(x3570, x3485, x69633);
  nand n3571(x3571, x3484, x3573);
  nand n3572(x3572, x3571, x3570);
  nand n3574(x3574, x3485, x69647);
  nand n3575(x3575, x3484, x3577);
  nand n3576(x3576, x3575, x3574);
  nand n3578(x3578, x3485, x69661);
  nand n3579(x3579, x3484, x3581);
  nand n3580(x3580, x3579, x3578);
  nand n3582(x3582, x3485, x69675);
  nand n3583(x3583, x3484, x3585);
  nand n3584(x3584, x3583, x3582);
  nand n3586(x3586, x3485, x69689);
  nand n3587(x3587, x3484, x3589);
  nand n3588(x3588, x3587, x3586);
  nand n3590(x3590, x3485, x69703);
  nand n3591(x3591, x3484, x3593);
  nand n3592(x3592, x3591, x3590);
  nand n3594(x3594, x3485, x69717);
  nand n3595(x3595, x3484, x3597);
  nand n3596(x3596, x3595, x3594);
  nand n3598(x3598, x3485, x69731);
  nand n3599(x3599, x3484, x3601);
  nand n3600(x3600, x3599, x3598);
  nand n3602(x3602, x3485, x69745);
  nand n3603(x3603, x3484, x3605);
  nand n3604(x3604, x3603, x3602);
  nand n3606(x3606, x3485, x69759);
  nand n3607(x3607, x3484, x3609);
  nand n3608(x3608, x3607, x3606);
  nand n3610(x3610, x3485, x69773);
  nand n3611(x3611, x3484, x3613);
  nand n3612(x3612, x3611, x3610);
  nand n3614(x3614, x2301, x71071);
  nand n3616(x3616, x3615, x69339);
  nand n3617(x3617, x3614, x3619);
  nand n3618(x3618, x3617, x3616);
  nand n3620(x3620, x3615, x69353);
  nand n3621(x3621, x3614, x3623);
  nand n3622(x3622, x3621, x3620);
  nand n3624(x3624, x3615, x69367);
  nand n3625(x3625, x3614, x3627);
  nand n3626(x3626, x3625, x3624);
  nand n3628(x3628, x3615, x69381);
  nand n3629(x3629, x3614, x3631);
  nand n3630(x3630, x3629, x3628);
  nand n3632(x3632, x3615, x69395);
  nand n3633(x3633, x3614, x3635);
  nand n3634(x3634, x3633, x3632);
  nand n3636(x3636, x3615, x69409);
  nand n3637(x3637, x3614, x3639);
  nand n3638(x3638, x3637, x3636);
  nand n3640(x3640, x3615, x69423);
  nand n3641(x3641, x3614, x3643);
  nand n3642(x3642, x3641, x3640);
  nand n3644(x3644, x3615, x69437);
  nand n3645(x3645, x3614, x3647);
  nand n3646(x3646, x3645, x3644);
  nand n3648(x3648, x3615, x69451);
  nand n3649(x3649, x3614, x3651);
  nand n3650(x3650, x3649, x3648);
  nand n3652(x3652, x3615, x69465);
  nand n3653(x3653, x3614, x3655);
  nand n3654(x3654, x3653, x3652);
  nand n3656(x3656, x3615, x69479);
  nand n3657(x3657, x3614, x3659);
  nand n3658(x3658, x3657, x3656);
  nand n3660(x3660, x3615, x69493);
  nand n3661(x3661, x3614, x3663);
  nand n3662(x3662, x3661, x3660);
  nand n3664(x3664, x3615, x69507);
  nand n3665(x3665, x3614, x3667);
  nand n3666(x3666, x3665, x3664);
  nand n3668(x3668, x3615, x69521);
  nand n3669(x3669, x3614, x3671);
  nand n3670(x3670, x3669, x3668);
  nand n3672(x3672, x3615, x69535);
  nand n3673(x3673, x3614, x3675);
  nand n3674(x3674, x3673, x3672);
  nand n3676(x3676, x3615, x69549);
  nand n3677(x3677, x3614, x3679);
  nand n3678(x3678, x3677, x3676);
  nand n3680(x3680, x3615, x69563);
  nand n3681(x3681, x3614, x3683);
  nand n3682(x3682, x3681, x3680);
  nand n3684(x3684, x3615, x69577);
  nand n3685(x3685, x3614, x3687);
  nand n3686(x3686, x3685, x3684);
  nand n3688(x3688, x3615, x69591);
  nand n3689(x3689, x3614, x3691);
  nand n3690(x3690, x3689, x3688);
  nand n3692(x3692, x3615, x69605);
  nand n3693(x3693, x3614, x3695);
  nand n3694(x3694, x3693, x3692);
  nand n3696(x3696, x3615, x69619);
  nand n3697(x3697, x3614, x3699);
  nand n3698(x3698, x3697, x3696);
  nand n3700(x3700, x3615, x69633);
  nand n3701(x3701, x3614, x3703);
  nand n3702(x3702, x3701, x3700);
  nand n3704(x3704, x3615, x69647);
  nand n3705(x3705, x3614, x3707);
  nand n3706(x3706, x3705, x3704);
  nand n3708(x3708, x3615, x69661);
  nand n3709(x3709, x3614, x3711);
  nand n3710(x3710, x3709, x3708);
  nand n3712(x3712, x3615, x69675);
  nand n3713(x3713, x3614, x3715);
  nand n3714(x3714, x3713, x3712);
  nand n3716(x3716, x3615, x69689);
  nand n3717(x3717, x3614, x3719);
  nand n3718(x3718, x3717, x3716);
  nand n3720(x3720, x3615, x69703);
  nand n3721(x3721, x3614, x3723);
  nand n3722(x3722, x3721, x3720);
  nand n3724(x3724, x3615, x69717);
  nand n3725(x3725, x3614, x3727);
  nand n3726(x3726, x3725, x3724);
  nand n3728(x3728, x3615, x69731);
  nand n3729(x3729, x3614, x3731);
  nand n3730(x3730, x3729, x3728);
  nand n3732(x3732, x3615, x69745);
  nand n3733(x3733, x3614, x3735);
  nand n3734(x3734, x3733, x3732);
  nand n3736(x3736, x3615, x69759);
  nand n3737(x3737, x3614, x3739);
  nand n3738(x3738, x3737, x3736);
  nand n3740(x3740, x3615, x69773);
  nand n3741(x3741, x3614, x3743);
  nand n3742(x3742, x3741, x3740);
  nand n3744(x3744, x2303, x71071);
  nand n3746(x3746, x3745, x69339);
  nand n3747(x3747, x3744, x3749);
  nand n3748(x3748, x3747, x3746);
  nand n3750(x3750, x3745, x69353);
  nand n3751(x3751, x3744, x3753);
  nand n3752(x3752, x3751, x3750);
  nand n3754(x3754, x3745, x69367);
  nand n3755(x3755, x3744, x3757);
  nand n3756(x3756, x3755, x3754);
  nand n3758(x3758, x3745, x69381);
  nand n3759(x3759, x3744, x3761);
  nand n3760(x3760, x3759, x3758);
  nand n3762(x3762, x3745, x69395);
  nand n3763(x3763, x3744, x3765);
  nand n3764(x3764, x3763, x3762);
  nand n3766(x3766, x3745, x69409);
  nand n3767(x3767, x3744, x3769);
  nand n3768(x3768, x3767, x3766);
  nand n3770(x3770, x3745, x69423);
  nand n3771(x3771, x3744, x3773);
  nand n3772(x3772, x3771, x3770);
  nand n3774(x3774, x3745, x69437);
  nand n3775(x3775, x3744, x3777);
  nand n3776(x3776, x3775, x3774);
  nand n3778(x3778, x3745, x69451);
  nand n3779(x3779, x3744, x3781);
  nand n3780(x3780, x3779, x3778);
  nand n3782(x3782, x3745, x69465);
  nand n3783(x3783, x3744, x3785);
  nand n3784(x3784, x3783, x3782);
  nand n3786(x3786, x3745, x69479);
  nand n3787(x3787, x3744, x3789);
  nand n3788(x3788, x3787, x3786);
  nand n3790(x3790, x3745, x69493);
  nand n3791(x3791, x3744, x3793);
  nand n3792(x3792, x3791, x3790);
  nand n3794(x3794, x3745, x69507);
  nand n3795(x3795, x3744, x3797);
  nand n3796(x3796, x3795, x3794);
  nand n3798(x3798, x3745, x69521);
  nand n3799(x3799, x3744, x3801);
  nand n3800(x3800, x3799, x3798);
  nand n3802(x3802, x3745, x69535);
  nand n3803(x3803, x3744, x3805);
  nand n3804(x3804, x3803, x3802);
  nand n3806(x3806, x3745, x69549);
  nand n3807(x3807, x3744, x3809);
  nand n3808(x3808, x3807, x3806);
  nand n3810(x3810, x3745, x69563);
  nand n3811(x3811, x3744, x3813);
  nand n3812(x3812, x3811, x3810);
  nand n3814(x3814, x3745, x69577);
  nand n3815(x3815, x3744, x3817);
  nand n3816(x3816, x3815, x3814);
  nand n3818(x3818, x3745, x69591);
  nand n3819(x3819, x3744, x3821);
  nand n3820(x3820, x3819, x3818);
  nand n3822(x3822, x3745, x69605);
  nand n3823(x3823, x3744, x3825);
  nand n3824(x3824, x3823, x3822);
  nand n3826(x3826, x3745, x69619);
  nand n3827(x3827, x3744, x3829);
  nand n3828(x3828, x3827, x3826);
  nand n3830(x3830, x3745, x69633);
  nand n3831(x3831, x3744, x3833);
  nand n3832(x3832, x3831, x3830);
  nand n3834(x3834, x3745, x69647);
  nand n3835(x3835, x3744, x3837);
  nand n3836(x3836, x3835, x3834);
  nand n3838(x3838, x3745, x69661);
  nand n3839(x3839, x3744, x3841);
  nand n3840(x3840, x3839, x3838);
  nand n3842(x3842, x3745, x69675);
  nand n3843(x3843, x3744, x3845);
  nand n3844(x3844, x3843, x3842);
  nand n3846(x3846, x3745, x69689);
  nand n3847(x3847, x3744, x3849);
  nand n3848(x3848, x3847, x3846);
  nand n3850(x3850, x3745, x69703);
  nand n3851(x3851, x3744, x3853);
  nand n3852(x3852, x3851, x3850);
  nand n3854(x3854, x3745, x69717);
  nand n3855(x3855, x3744, x3857);
  nand n3856(x3856, x3855, x3854);
  nand n3858(x3858, x3745, x69731);
  nand n3859(x3859, x3744, x3861);
  nand n3860(x3860, x3859, x3858);
  nand n3862(x3862, x3745, x69745);
  nand n3863(x3863, x3744, x3865);
  nand n3864(x3864, x3863, x3862);
  nand n3866(x3866, x3745, x69759);
  nand n3867(x3867, x3744, x3869);
  nand n3868(x3868, x3867, x3866);
  nand n3870(x3870, x3745, x69773);
  nand n3871(x3871, x3744, x3873);
  nand n3872(x3872, x3871, x3870);
  nand n3874(x3874, x2305, x71071);
  nand n3876(x3876, x3875, x69339);
  nand n3877(x3877, x3874, x3879);
  nand n3878(x3878, x3877, x3876);
  nand n3880(x3880, x3875, x69353);
  nand n3881(x3881, x3874, x3883);
  nand n3882(x3882, x3881, x3880);
  nand n3884(x3884, x3875, x69367);
  nand n3885(x3885, x3874, x3887);
  nand n3886(x3886, x3885, x3884);
  nand n3888(x3888, x3875, x69381);
  nand n3889(x3889, x3874, x3891);
  nand n3890(x3890, x3889, x3888);
  nand n3892(x3892, x3875, x69395);
  nand n3893(x3893, x3874, x3895);
  nand n3894(x3894, x3893, x3892);
  nand n3896(x3896, x3875, x69409);
  nand n3897(x3897, x3874, x3899);
  nand n3898(x3898, x3897, x3896);
  nand n3900(x3900, x3875, x69423);
  nand n3901(x3901, x3874, x3903);
  nand n3902(x3902, x3901, x3900);
  nand n3904(x3904, x3875, x69437);
  nand n3905(x3905, x3874, x3907);
  nand n3906(x3906, x3905, x3904);
  nand n3908(x3908, x3875, x69451);
  nand n3909(x3909, x3874, x3911);
  nand n3910(x3910, x3909, x3908);
  nand n3912(x3912, x3875, x69465);
  nand n3913(x3913, x3874, x3915);
  nand n3914(x3914, x3913, x3912);
  nand n3916(x3916, x3875, x69479);
  nand n3917(x3917, x3874, x3919);
  nand n3918(x3918, x3917, x3916);
  nand n3920(x3920, x3875, x69493);
  nand n3921(x3921, x3874, x3923);
  nand n3922(x3922, x3921, x3920);
  nand n3924(x3924, x3875, x69507);
  nand n3925(x3925, x3874, x3927);
  nand n3926(x3926, x3925, x3924);
  nand n3928(x3928, x3875, x69521);
  nand n3929(x3929, x3874, x3931);
  nand n3930(x3930, x3929, x3928);
  nand n3932(x3932, x3875, x69535);
  nand n3933(x3933, x3874, x3935);
  nand n3934(x3934, x3933, x3932);
  nand n3936(x3936, x3875, x69549);
  nand n3937(x3937, x3874, x3939);
  nand n3938(x3938, x3937, x3936);
  nand n3940(x3940, x3875, x69563);
  nand n3941(x3941, x3874, x3943);
  nand n3942(x3942, x3941, x3940);
  nand n3944(x3944, x3875, x69577);
  nand n3945(x3945, x3874, x3947);
  nand n3946(x3946, x3945, x3944);
  nand n3948(x3948, x3875, x69591);
  nand n3949(x3949, x3874, x3951);
  nand n3950(x3950, x3949, x3948);
  nand n3952(x3952, x3875, x69605);
  nand n3953(x3953, x3874, x3955);
  nand n3954(x3954, x3953, x3952);
  nand n3956(x3956, x3875, x69619);
  nand n3957(x3957, x3874, x3959);
  nand n3958(x3958, x3957, x3956);
  nand n3960(x3960, x3875, x69633);
  nand n3961(x3961, x3874, x3963);
  nand n3962(x3962, x3961, x3960);
  nand n3964(x3964, x3875, x69647);
  nand n3965(x3965, x3874, x3967);
  nand n3966(x3966, x3965, x3964);
  nand n3968(x3968, x3875, x69661);
  nand n3969(x3969, x3874, x3971);
  nand n3970(x3970, x3969, x3968);
  nand n3972(x3972, x3875, x69675);
  nand n3973(x3973, x3874, x3975);
  nand n3974(x3974, x3973, x3972);
  nand n3976(x3976, x3875, x69689);
  nand n3977(x3977, x3874, x3979);
  nand n3978(x3978, x3977, x3976);
  nand n3980(x3980, x3875, x69703);
  nand n3981(x3981, x3874, x3983);
  nand n3982(x3982, x3981, x3980);
  nand n3984(x3984, x3875, x69717);
  nand n3985(x3985, x3874, x3987);
  nand n3986(x3986, x3985, x3984);
  nand n3988(x3988, x3875, x69731);
  nand n3989(x3989, x3874, x3991);
  nand n3990(x3990, x3989, x3988);
  nand n3992(x3992, x3875, x69745);
  nand n3993(x3993, x3874, x3995);
  nand n3994(x3994, x3993, x3992);
  nand n3996(x3996, x3875, x69759);
  nand n3997(x3997, x3874, x3999);
  nand n3998(x3998, x3997, x3996);
  nand n4000(x4000, x3875, x69773);
  nand n4001(x4001, x3874, x4003);
  nand n4002(x4002, x4001, x4000);
  nand n4004(x4004, x2307, x71071);
  nand n4006(x4006, x4005, x69339);
  nand n4007(x4007, x4004, x4009);
  nand n4008(x4008, x4007, x4006);
  nand n4010(x4010, x4005, x69353);
  nand n4011(x4011, x4004, x4013);
  nand n4012(x4012, x4011, x4010);
  nand n4014(x4014, x4005, x69367);
  nand n4015(x4015, x4004, x4017);
  nand n4016(x4016, x4015, x4014);
  nand n4018(x4018, x4005, x69381);
  nand n4019(x4019, x4004, x4021);
  nand n4020(x4020, x4019, x4018);
  nand n4022(x4022, x4005, x69395);
  nand n4023(x4023, x4004, x4025);
  nand n4024(x4024, x4023, x4022);
  nand n4026(x4026, x4005, x69409);
  nand n4027(x4027, x4004, x4029);
  nand n4028(x4028, x4027, x4026);
  nand n4030(x4030, x4005, x69423);
  nand n4031(x4031, x4004, x4033);
  nand n4032(x4032, x4031, x4030);
  nand n4034(x4034, x4005, x69437);
  nand n4035(x4035, x4004, x4037);
  nand n4036(x4036, x4035, x4034);
  nand n4038(x4038, x4005, x69451);
  nand n4039(x4039, x4004, x4041);
  nand n4040(x4040, x4039, x4038);
  nand n4042(x4042, x4005, x69465);
  nand n4043(x4043, x4004, x4045);
  nand n4044(x4044, x4043, x4042);
  nand n4046(x4046, x4005, x69479);
  nand n4047(x4047, x4004, x4049);
  nand n4048(x4048, x4047, x4046);
  nand n4050(x4050, x4005, x69493);
  nand n4051(x4051, x4004, x4053);
  nand n4052(x4052, x4051, x4050);
  nand n4054(x4054, x4005, x69507);
  nand n4055(x4055, x4004, x4057);
  nand n4056(x4056, x4055, x4054);
  nand n4058(x4058, x4005, x69521);
  nand n4059(x4059, x4004, x4061);
  nand n4060(x4060, x4059, x4058);
  nand n4062(x4062, x4005, x69535);
  nand n4063(x4063, x4004, x4065);
  nand n4064(x4064, x4063, x4062);
  nand n4066(x4066, x4005, x69549);
  nand n4067(x4067, x4004, x4069);
  nand n4068(x4068, x4067, x4066);
  nand n4070(x4070, x4005, x69563);
  nand n4071(x4071, x4004, x4073);
  nand n4072(x4072, x4071, x4070);
  nand n4074(x4074, x4005, x69577);
  nand n4075(x4075, x4004, x4077);
  nand n4076(x4076, x4075, x4074);
  nand n4078(x4078, x4005, x69591);
  nand n4079(x4079, x4004, x4081);
  nand n4080(x4080, x4079, x4078);
  nand n4082(x4082, x4005, x69605);
  nand n4083(x4083, x4004, x4085);
  nand n4084(x4084, x4083, x4082);
  nand n4086(x4086, x4005, x69619);
  nand n4087(x4087, x4004, x4089);
  nand n4088(x4088, x4087, x4086);
  nand n4090(x4090, x4005, x69633);
  nand n4091(x4091, x4004, x4093);
  nand n4092(x4092, x4091, x4090);
  nand n4094(x4094, x4005, x69647);
  nand n4095(x4095, x4004, x4097);
  nand n4096(x4096, x4095, x4094);
  nand n4098(x4098, x4005, x69661);
  nand n4099(x4099, x4004, x4101);
  nand n4100(x4100, x4099, x4098);
  nand n4102(x4102, x4005, x69675);
  nand n4103(x4103, x4004, x4105);
  nand n4104(x4104, x4103, x4102);
  nand n4106(x4106, x4005, x69689);
  nand n4107(x4107, x4004, x4109);
  nand n4108(x4108, x4107, x4106);
  nand n4110(x4110, x4005, x69703);
  nand n4111(x4111, x4004, x4113);
  nand n4112(x4112, x4111, x4110);
  nand n4114(x4114, x4005, x69717);
  nand n4115(x4115, x4004, x4117);
  nand n4116(x4116, x4115, x4114);
  nand n4118(x4118, x4005, x69731);
  nand n4119(x4119, x4004, x4121);
  nand n4120(x4120, x4119, x4118);
  nand n4122(x4122, x4005, x69745);
  nand n4123(x4123, x4004, x4125);
  nand n4124(x4124, x4123, x4122);
  nand n4126(x4126, x4005, x69759);
  nand n4127(x4127, x4004, x4129);
  nand n4128(x4128, x4127, x4126);
  nand n4130(x4130, x4005, x69773);
  nand n4131(x4131, x4004, x4133);
  nand n4132(x4132, x4131, x4130);
  nand n4134(x4134, x2309, x71071);
  nand n4136(x4136, x4135, x69339);
  nand n4137(x4137, x4134, x4139);
  nand n4138(x4138, x4137, x4136);
  nand n4140(x4140, x4135, x69353);
  nand n4141(x4141, x4134, x4143);
  nand n4142(x4142, x4141, x4140);
  nand n4144(x4144, x4135, x69367);
  nand n4145(x4145, x4134, x4147);
  nand n4146(x4146, x4145, x4144);
  nand n4148(x4148, x4135, x69381);
  nand n4149(x4149, x4134, x4151);
  nand n4150(x4150, x4149, x4148);
  nand n4152(x4152, x4135, x69395);
  nand n4153(x4153, x4134, x4155);
  nand n4154(x4154, x4153, x4152);
  nand n4156(x4156, x4135, x69409);
  nand n4157(x4157, x4134, x4159);
  nand n4158(x4158, x4157, x4156);
  nand n4160(x4160, x4135, x69423);
  nand n4161(x4161, x4134, x4163);
  nand n4162(x4162, x4161, x4160);
  nand n4164(x4164, x4135, x69437);
  nand n4165(x4165, x4134, x4167);
  nand n4166(x4166, x4165, x4164);
  nand n4168(x4168, x4135, x69451);
  nand n4169(x4169, x4134, x4171);
  nand n4170(x4170, x4169, x4168);
  nand n4172(x4172, x4135, x69465);
  nand n4173(x4173, x4134, x4175);
  nand n4174(x4174, x4173, x4172);
  nand n4176(x4176, x4135, x69479);
  nand n4177(x4177, x4134, x4179);
  nand n4178(x4178, x4177, x4176);
  nand n4180(x4180, x4135, x69493);
  nand n4181(x4181, x4134, x4183);
  nand n4182(x4182, x4181, x4180);
  nand n4184(x4184, x4135, x69507);
  nand n4185(x4185, x4134, x4187);
  nand n4186(x4186, x4185, x4184);
  nand n4188(x4188, x4135, x69521);
  nand n4189(x4189, x4134, x4191);
  nand n4190(x4190, x4189, x4188);
  nand n4192(x4192, x4135, x69535);
  nand n4193(x4193, x4134, x4195);
  nand n4194(x4194, x4193, x4192);
  nand n4196(x4196, x4135, x69549);
  nand n4197(x4197, x4134, x4199);
  nand n4198(x4198, x4197, x4196);
  nand n4200(x4200, x4135, x69563);
  nand n4201(x4201, x4134, x4203);
  nand n4202(x4202, x4201, x4200);
  nand n4204(x4204, x4135, x69577);
  nand n4205(x4205, x4134, x4207);
  nand n4206(x4206, x4205, x4204);
  nand n4208(x4208, x4135, x69591);
  nand n4209(x4209, x4134, x4211);
  nand n4210(x4210, x4209, x4208);
  nand n4212(x4212, x4135, x69605);
  nand n4213(x4213, x4134, x4215);
  nand n4214(x4214, x4213, x4212);
  nand n4216(x4216, x4135, x69619);
  nand n4217(x4217, x4134, x4219);
  nand n4218(x4218, x4217, x4216);
  nand n4220(x4220, x4135, x69633);
  nand n4221(x4221, x4134, x4223);
  nand n4222(x4222, x4221, x4220);
  nand n4224(x4224, x4135, x69647);
  nand n4225(x4225, x4134, x4227);
  nand n4226(x4226, x4225, x4224);
  nand n4228(x4228, x4135, x69661);
  nand n4229(x4229, x4134, x4231);
  nand n4230(x4230, x4229, x4228);
  nand n4232(x4232, x4135, x69675);
  nand n4233(x4233, x4134, x4235);
  nand n4234(x4234, x4233, x4232);
  nand n4236(x4236, x4135, x69689);
  nand n4237(x4237, x4134, x4239);
  nand n4238(x4238, x4237, x4236);
  nand n4240(x4240, x4135, x69703);
  nand n4241(x4241, x4134, x4243);
  nand n4242(x4242, x4241, x4240);
  nand n4244(x4244, x4135, x69717);
  nand n4245(x4245, x4134, x4247);
  nand n4246(x4246, x4245, x4244);
  nand n4248(x4248, x4135, x69731);
  nand n4249(x4249, x4134, x4251);
  nand n4250(x4250, x4249, x4248);
  nand n4252(x4252, x4135, x69745);
  nand n4253(x4253, x4134, x4255);
  nand n4254(x4254, x4253, x4252);
  nand n4256(x4256, x4135, x69759);
  nand n4257(x4257, x4134, x4259);
  nand n4258(x4258, x4257, x4256);
  nand n4260(x4260, x4135, x69773);
  nand n4261(x4261, x4134, x4263);
  nand n4262(x4262, x4261, x4260);
  nand n4264(x4264, x2311, x71071);
  nand n4266(x4266, x4265, x69339);
  nand n4267(x4267, x4264, x4269);
  nand n4268(x4268, x4267, x4266);
  nand n4270(x4270, x4265, x69353);
  nand n4271(x4271, x4264, x4273);
  nand n4272(x4272, x4271, x4270);
  nand n4274(x4274, x4265, x69367);
  nand n4275(x4275, x4264, x4277);
  nand n4276(x4276, x4275, x4274);
  nand n4278(x4278, x4265, x69381);
  nand n4279(x4279, x4264, x4281);
  nand n4280(x4280, x4279, x4278);
  nand n4282(x4282, x4265, x69395);
  nand n4283(x4283, x4264, x4285);
  nand n4284(x4284, x4283, x4282);
  nand n4286(x4286, x4265, x69409);
  nand n4287(x4287, x4264, x4289);
  nand n4288(x4288, x4287, x4286);
  nand n4290(x4290, x4265, x69423);
  nand n4291(x4291, x4264, x4293);
  nand n4292(x4292, x4291, x4290);
  nand n4294(x4294, x4265, x69437);
  nand n4295(x4295, x4264, x4297);
  nand n4296(x4296, x4295, x4294);
  nand n4298(x4298, x4265, x69451);
  nand n4299(x4299, x4264, x4301);
  nand n4300(x4300, x4299, x4298);
  nand n4302(x4302, x4265, x69465);
  nand n4303(x4303, x4264, x4305);
  nand n4304(x4304, x4303, x4302);
  nand n4306(x4306, x4265, x69479);
  nand n4307(x4307, x4264, x4309);
  nand n4308(x4308, x4307, x4306);
  nand n4310(x4310, x4265, x69493);
  nand n4311(x4311, x4264, x4313);
  nand n4312(x4312, x4311, x4310);
  nand n4314(x4314, x4265, x69507);
  nand n4315(x4315, x4264, x4317);
  nand n4316(x4316, x4315, x4314);
  nand n4318(x4318, x4265, x69521);
  nand n4319(x4319, x4264, x4321);
  nand n4320(x4320, x4319, x4318);
  nand n4322(x4322, x4265, x69535);
  nand n4323(x4323, x4264, x4325);
  nand n4324(x4324, x4323, x4322);
  nand n4326(x4326, x4265, x69549);
  nand n4327(x4327, x4264, x4329);
  nand n4328(x4328, x4327, x4326);
  nand n4330(x4330, x4265, x69563);
  nand n4331(x4331, x4264, x4333);
  nand n4332(x4332, x4331, x4330);
  nand n4334(x4334, x4265, x69577);
  nand n4335(x4335, x4264, x4337);
  nand n4336(x4336, x4335, x4334);
  nand n4338(x4338, x4265, x69591);
  nand n4339(x4339, x4264, x4341);
  nand n4340(x4340, x4339, x4338);
  nand n4342(x4342, x4265, x69605);
  nand n4343(x4343, x4264, x4345);
  nand n4344(x4344, x4343, x4342);
  nand n4346(x4346, x4265, x69619);
  nand n4347(x4347, x4264, x4349);
  nand n4348(x4348, x4347, x4346);
  nand n4350(x4350, x4265, x69633);
  nand n4351(x4351, x4264, x4353);
  nand n4352(x4352, x4351, x4350);
  nand n4354(x4354, x4265, x69647);
  nand n4355(x4355, x4264, x4357);
  nand n4356(x4356, x4355, x4354);
  nand n4358(x4358, x4265, x69661);
  nand n4359(x4359, x4264, x4361);
  nand n4360(x4360, x4359, x4358);
  nand n4362(x4362, x4265, x69675);
  nand n4363(x4363, x4264, x4365);
  nand n4364(x4364, x4363, x4362);
  nand n4366(x4366, x4265, x69689);
  nand n4367(x4367, x4264, x4369);
  nand n4368(x4368, x4367, x4366);
  nand n4370(x4370, x4265, x69703);
  nand n4371(x4371, x4264, x4373);
  nand n4372(x4372, x4371, x4370);
  nand n4374(x4374, x4265, x69717);
  nand n4375(x4375, x4264, x4377);
  nand n4376(x4376, x4375, x4374);
  nand n4378(x4378, x4265, x69731);
  nand n4379(x4379, x4264, x4381);
  nand n4380(x4380, x4379, x4378);
  nand n4382(x4382, x4265, x69745);
  nand n4383(x4383, x4264, x4385);
  nand n4384(x4384, x4383, x4382);
  nand n4386(x4386, x4265, x69759);
  nand n4387(x4387, x4264, x4389);
  nand n4388(x4388, x4387, x4386);
  nand n4390(x4390, x4265, x69773);
  nand n4391(x4391, x4264, x4393);
  nand n4392(x4392, x4391, x4390);
  nand n4394(x4394, x2297, x71073);
  nand n4396(x4396, x4395, x69789);
  nand n4397(x4397, x4394, x4399);
  nand n4398(x4398, x4397, x4396);
  nand n4400(x4400, x4395, x69803);
  nand n4401(x4401, x4394, x4405);
  nand n4402(x4402, x4401, x4400);
  nand n4406(x4406, x4395, x69817);
  nand n4407(x4407, x4394, x4409);
  nand n4408(x4408, x4407, x4406);
  nand n4410(x4410, x4395, x69831);
  nand n4411(x4411, x4394, x4413);
  nand n4412(x4412, x4411, x4410);
  nand n4414(x4414, x4395, x69845);
  nand n4415(x4415, x4394, x4417);
  nand n4416(x4416, x4415, x4414);
  nand n4418(x4418, x4395, x69859);
  nand n4419(x4419, x4394, x4421);
  nand n4420(x4420, x4419, x4418);
  nand n4422(x4422, x4395, x69873);
  nand n4423(x4423, x4394, x4425);
  nand n4424(x4424, x4423, x4422);
  nand n4426(x4426, x4395, x69887);
  nand n4427(x4427, x4394, x4429);
  nand n4428(x4428, x4427, x4426);
  nand n4430(x4430, x4395, x69901);
  nand n4431(x4431, x4394, x4433);
  nand n4432(x4432, x4431, x4430);
  nand n4434(x4434, x4395, x69915);
  nand n4435(x4435, x4394, x4437);
  nand n4436(x4436, x4435, x4434);
  nand n4438(x4438, x4395, x69929);
  nand n4439(x4439, x4394, x4441);
  nand n4440(x4440, x4439, x4438);
  nand n4442(x4442, x4395, x69943);
  nand n4443(x4443, x4394, x4445);
  nand n4444(x4444, x4443, x4442);
  nand n4446(x4446, x4395, x69957);
  nand n4447(x4447, x4394, x4449);
  nand n4448(x4448, x4447, x4446);
  nand n4450(x4450, x4395, x69971);
  nand n4451(x4451, x4394, x4453);
  nand n4452(x4452, x4451, x4450);
  nand n4454(x4454, x4395, x69985);
  nand n4455(x4455, x4394, x4457);
  nand n4456(x4456, x4455, x4454);
  nand n4458(x4458, x4395, x69999);
  nand n4459(x4459, x4394, x4461);
  nand n4460(x4460, x4459, x4458);
  nand n4462(x4462, x4395, x70013);
  nand n4463(x4463, x4394, x4465);
  nand n4464(x4464, x4463, x4462);
  nand n4466(x4466, x4395, x70027);
  nand n4467(x4467, x4394, x4469);
  nand n4468(x4468, x4467, x4466);
  nand n4470(x4470, x4395, x70041);
  nand n4471(x4471, x4394, x4473);
  nand n4472(x4472, x4471, x4470);
  nand n4474(x4474, x4395, x70055);
  nand n4475(x4475, x4394, x4477);
  nand n4476(x4476, x4475, x4474);
  nand n4478(x4478, x4395, x70069);
  nand n4479(x4479, x4394, x4481);
  nand n4480(x4480, x4479, x4478);
  nand n4482(x4482, x4395, x70083);
  nand n4483(x4483, x4394, x4485);
  nand n4484(x4484, x4483, x4482);
  nand n4486(x4486, x4395, x70097);
  nand n4487(x4487, x4394, x4489);
  nand n4488(x4488, x4487, x4486);
  nand n4490(x4490, x4395, x70111);
  nand n4491(x4491, x4394, x4493);
  nand n4492(x4492, x4491, x4490);
  nand n4494(x4494, x4395, x70125);
  nand n4495(x4495, x4394, x4497);
  nand n4496(x4496, x4495, x4494);
  nand n4498(x4498, x4395, x70139);
  nand n4499(x4499, x4394, x4501);
  nand n4500(x4500, x4499, x4498);
  nand n4502(x4502, x4395, x70153);
  nand n4503(x4503, x4394, x4505);
  nand n4504(x4504, x4503, x4502);
  nand n4506(x4506, x4395, x70167);
  nand n4507(x4507, x4394, x4509);
  nand n4508(x4508, x4507, x4506);
  nand n4510(x4510, x4395, x70181);
  nand n4511(x4511, x4394, x4513);
  nand n4512(x4512, x4511, x4510);
  nand n4514(x4514, x4395, x70195);
  nand n4515(x4515, x4394, x4517);
  nand n4516(x4516, x4515, x4514);
  nand n4518(x4518, x4395, x70209);
  nand n4519(x4519, x4394, x4521);
  nand n4520(x4520, x4519, x4518);
  nand n4522(x4522, x4395, x70223);
  nand n4523(x4523, x4394, x4525);
  nand n4524(x4524, x4523, x4522);
  nand n4526(x4526, x2299, x71073);
  nand n4528(x4528, x4527, x69789);
  nand n4529(x4529, x4526, x4531);
  nand n4530(x4530, x4529, x4528);
  nand n4532(x4532, x4527, x69803);
  nand n4533(x4533, x4526, x4535);
  nand n4534(x4534, x4533, x4532);
  nand n4536(x4536, x4527, x69817);
  nand n4537(x4537, x4526, x4539);
  nand n4538(x4538, x4537, x4536);
  nand n4540(x4540, x4527, x69831);
  nand n4541(x4541, x4526, x4543);
  nand n4542(x4542, x4541, x4540);
  nand n4544(x4544, x4527, x69845);
  nand n4545(x4545, x4526, x4547);
  nand n4546(x4546, x4545, x4544);
  nand n4548(x4548, x4527, x69859);
  nand n4549(x4549, x4526, x4551);
  nand n4550(x4550, x4549, x4548);
  nand n4552(x4552, x4527, x69873);
  nand n4553(x4553, x4526, x4555);
  nand n4554(x4554, x4553, x4552);
  nand n4556(x4556, x4527, x69887);
  nand n4557(x4557, x4526, x4559);
  nand n4558(x4558, x4557, x4556);
  nand n4560(x4560, x4527, x69901);
  nand n4561(x4561, x4526, x4563);
  nand n4562(x4562, x4561, x4560);
  nand n4564(x4564, x4527, x69915);
  nand n4565(x4565, x4526, x4567);
  nand n4566(x4566, x4565, x4564);
  nand n4568(x4568, x4527, x69929);
  nand n4569(x4569, x4526, x4571);
  nand n4570(x4570, x4569, x4568);
  nand n4572(x4572, x4527, x69943);
  nand n4573(x4573, x4526, x4575);
  nand n4574(x4574, x4573, x4572);
  nand n4576(x4576, x4527, x69957);
  nand n4577(x4577, x4526, x4579);
  nand n4578(x4578, x4577, x4576);
  nand n4580(x4580, x4527, x69971);
  nand n4581(x4581, x4526, x4583);
  nand n4582(x4582, x4581, x4580);
  nand n4584(x4584, x4527, x69985);
  nand n4585(x4585, x4526, x4587);
  nand n4586(x4586, x4585, x4584);
  nand n4588(x4588, x4527, x69999);
  nand n4589(x4589, x4526, x4591);
  nand n4590(x4590, x4589, x4588);
  nand n4592(x4592, x4527, x70013);
  nand n4593(x4593, x4526, x4595);
  nand n4594(x4594, x4593, x4592);
  nand n4596(x4596, x4527, x70027);
  nand n4597(x4597, x4526, x4599);
  nand n4598(x4598, x4597, x4596);
  nand n4600(x4600, x4527, x70041);
  nand n4601(x4601, x4526, x4603);
  nand n4602(x4602, x4601, x4600);
  nand n4604(x4604, x4527, x70055);
  nand n4605(x4605, x4526, x4607);
  nand n4606(x4606, x4605, x4604);
  nand n4608(x4608, x4527, x70069);
  nand n4609(x4609, x4526, x4611);
  nand n4610(x4610, x4609, x4608);
  nand n4612(x4612, x4527, x70083);
  nand n4613(x4613, x4526, x4615);
  nand n4614(x4614, x4613, x4612);
  nand n4616(x4616, x4527, x70097);
  nand n4617(x4617, x4526, x4619);
  nand n4618(x4618, x4617, x4616);
  nand n4620(x4620, x4527, x70111);
  nand n4621(x4621, x4526, x4623);
  nand n4622(x4622, x4621, x4620);
  nand n4624(x4624, x4527, x70125);
  nand n4625(x4625, x4526, x4627);
  nand n4626(x4626, x4625, x4624);
  nand n4628(x4628, x4527, x70139);
  nand n4629(x4629, x4526, x4631);
  nand n4630(x4630, x4629, x4628);
  nand n4632(x4632, x4527, x70153);
  nand n4633(x4633, x4526, x4635);
  nand n4634(x4634, x4633, x4632);
  nand n4636(x4636, x4527, x70167);
  nand n4637(x4637, x4526, x4639);
  nand n4638(x4638, x4637, x4636);
  nand n4640(x4640, x4527, x70181);
  nand n4641(x4641, x4526, x4643);
  nand n4642(x4642, x4641, x4640);
  nand n4644(x4644, x4527, x70195);
  nand n4645(x4645, x4526, x4647);
  nand n4646(x4646, x4645, x4644);
  nand n4648(x4648, x4527, x70209);
  nand n4649(x4649, x4526, x4651);
  nand n4650(x4650, x4649, x4648);
  nand n4652(x4652, x4527, x70223);
  nand n4653(x4653, x4526, x4655);
  nand n4654(x4654, x4653, x4652);
  nand n4656(x4656, x2301, x71073);
  nand n4658(x4658, x4657, x69789);
  nand n4659(x4659, x4656, x4661);
  nand n4660(x4660, x4659, x4658);
  nand n4662(x4662, x4657, x69803);
  nand n4663(x4663, x4656, x4665);
  nand n4664(x4664, x4663, x4662);
  nand n4666(x4666, x4657, x69817);
  nand n4667(x4667, x4656, x4669);
  nand n4668(x4668, x4667, x4666);
  nand n4670(x4670, x4657, x69831);
  nand n4671(x4671, x4656, x4673);
  nand n4672(x4672, x4671, x4670);
  nand n4674(x4674, x4657, x69845);
  nand n4675(x4675, x4656, x4677);
  nand n4676(x4676, x4675, x4674);
  nand n4678(x4678, x4657, x69859);
  nand n4679(x4679, x4656, x4681);
  nand n4680(x4680, x4679, x4678);
  nand n4682(x4682, x4657, x69873);
  nand n4683(x4683, x4656, x4685);
  nand n4684(x4684, x4683, x4682);
  nand n4686(x4686, x4657, x69887);
  nand n4687(x4687, x4656, x4689);
  nand n4688(x4688, x4687, x4686);
  nand n4690(x4690, x4657, x69901);
  nand n4691(x4691, x4656, x4693);
  nand n4692(x4692, x4691, x4690);
  nand n4694(x4694, x4657, x69915);
  nand n4695(x4695, x4656, x4697);
  nand n4696(x4696, x4695, x4694);
  nand n4698(x4698, x4657, x69929);
  nand n4699(x4699, x4656, x4701);
  nand n4700(x4700, x4699, x4698);
  nand n4702(x4702, x4657, x69943);
  nand n4703(x4703, x4656, x4705);
  nand n4704(x4704, x4703, x4702);
  nand n4706(x4706, x4657, x69957);
  nand n4707(x4707, x4656, x4709);
  nand n4708(x4708, x4707, x4706);
  nand n4710(x4710, x4657, x69971);
  nand n4711(x4711, x4656, x4713);
  nand n4712(x4712, x4711, x4710);
  nand n4714(x4714, x4657, x69985);
  nand n4715(x4715, x4656, x4717);
  nand n4716(x4716, x4715, x4714);
  nand n4718(x4718, x4657, x69999);
  nand n4719(x4719, x4656, x4721);
  nand n4720(x4720, x4719, x4718);
  nand n4722(x4722, x4657, x70013);
  nand n4723(x4723, x4656, x4725);
  nand n4724(x4724, x4723, x4722);
  nand n4726(x4726, x4657, x70027);
  nand n4727(x4727, x4656, x4729);
  nand n4728(x4728, x4727, x4726);
  nand n4730(x4730, x4657, x70041);
  nand n4731(x4731, x4656, x4733);
  nand n4732(x4732, x4731, x4730);
  nand n4734(x4734, x4657, x70055);
  nand n4735(x4735, x4656, x4737);
  nand n4736(x4736, x4735, x4734);
  nand n4738(x4738, x4657, x70069);
  nand n4739(x4739, x4656, x4741);
  nand n4740(x4740, x4739, x4738);
  nand n4742(x4742, x4657, x70083);
  nand n4743(x4743, x4656, x4745);
  nand n4744(x4744, x4743, x4742);
  nand n4746(x4746, x4657, x70097);
  nand n4747(x4747, x4656, x4749);
  nand n4748(x4748, x4747, x4746);
  nand n4750(x4750, x4657, x70111);
  nand n4751(x4751, x4656, x4753);
  nand n4752(x4752, x4751, x4750);
  nand n4754(x4754, x4657, x70125);
  nand n4755(x4755, x4656, x4757);
  nand n4756(x4756, x4755, x4754);
  nand n4758(x4758, x4657, x70139);
  nand n4759(x4759, x4656, x4761);
  nand n4760(x4760, x4759, x4758);
  nand n4762(x4762, x4657, x70153);
  nand n4763(x4763, x4656, x4765);
  nand n4764(x4764, x4763, x4762);
  nand n4766(x4766, x4657, x70167);
  nand n4767(x4767, x4656, x4769);
  nand n4768(x4768, x4767, x4766);
  nand n4770(x4770, x4657, x70181);
  nand n4771(x4771, x4656, x4773);
  nand n4772(x4772, x4771, x4770);
  nand n4774(x4774, x4657, x70195);
  nand n4775(x4775, x4656, x4777);
  nand n4776(x4776, x4775, x4774);
  nand n4778(x4778, x4657, x70209);
  nand n4779(x4779, x4656, x4781);
  nand n4780(x4780, x4779, x4778);
  nand n4782(x4782, x4657, x70223);
  nand n4783(x4783, x4656, x4785);
  nand n4784(x4784, x4783, x4782);
  nand n4786(x4786, x2303, x71073);
  nand n4788(x4788, x4787, x69789);
  nand n4789(x4789, x4786, x4791);
  nand n4790(x4790, x4789, x4788);
  nand n4792(x4792, x4787, x69803);
  nand n4793(x4793, x4786, x4795);
  nand n4794(x4794, x4793, x4792);
  nand n4796(x4796, x4787, x69817);
  nand n4797(x4797, x4786, x4799);
  nand n4798(x4798, x4797, x4796);
  nand n4800(x4800, x4787, x69831);
  nand n4801(x4801, x4786, x4803);
  nand n4802(x4802, x4801, x4800);
  nand n4804(x4804, x4787, x69845);
  nand n4805(x4805, x4786, x4807);
  nand n4806(x4806, x4805, x4804);
  nand n4808(x4808, x4787, x69859);
  nand n4809(x4809, x4786, x4811);
  nand n4810(x4810, x4809, x4808);
  nand n4812(x4812, x4787, x69873);
  nand n4813(x4813, x4786, x4815);
  nand n4814(x4814, x4813, x4812);
  nand n4816(x4816, x4787, x69887);
  nand n4817(x4817, x4786, x4819);
  nand n4818(x4818, x4817, x4816);
  nand n4820(x4820, x4787, x69901);
  nand n4821(x4821, x4786, x4823);
  nand n4822(x4822, x4821, x4820);
  nand n4824(x4824, x4787, x69915);
  nand n4825(x4825, x4786, x4827);
  nand n4826(x4826, x4825, x4824);
  nand n4828(x4828, x4787, x69929);
  nand n4829(x4829, x4786, x4831);
  nand n4830(x4830, x4829, x4828);
  nand n4832(x4832, x4787, x69943);
  nand n4833(x4833, x4786, x4835);
  nand n4834(x4834, x4833, x4832);
  nand n4836(x4836, x4787, x69957);
  nand n4837(x4837, x4786, x4839);
  nand n4838(x4838, x4837, x4836);
  nand n4840(x4840, x4787, x69971);
  nand n4841(x4841, x4786, x4843);
  nand n4842(x4842, x4841, x4840);
  nand n4844(x4844, x4787, x69985);
  nand n4845(x4845, x4786, x4847);
  nand n4846(x4846, x4845, x4844);
  nand n4848(x4848, x4787, x69999);
  nand n4849(x4849, x4786, x4851);
  nand n4850(x4850, x4849, x4848);
  nand n4852(x4852, x4787, x70013);
  nand n4853(x4853, x4786, x4855);
  nand n4854(x4854, x4853, x4852);
  nand n4856(x4856, x4787, x70027);
  nand n4857(x4857, x4786, x4859);
  nand n4858(x4858, x4857, x4856);
  nand n4860(x4860, x4787, x70041);
  nand n4861(x4861, x4786, x4863);
  nand n4862(x4862, x4861, x4860);
  nand n4864(x4864, x4787, x70055);
  nand n4865(x4865, x4786, x4867);
  nand n4866(x4866, x4865, x4864);
  nand n4868(x4868, x4787, x70069);
  nand n4869(x4869, x4786, x4871);
  nand n4870(x4870, x4869, x4868);
  nand n4872(x4872, x4787, x70083);
  nand n4873(x4873, x4786, x4875);
  nand n4874(x4874, x4873, x4872);
  nand n4876(x4876, x4787, x70097);
  nand n4877(x4877, x4786, x4879);
  nand n4878(x4878, x4877, x4876);
  nand n4880(x4880, x4787, x70111);
  nand n4881(x4881, x4786, x4883);
  nand n4882(x4882, x4881, x4880);
  nand n4884(x4884, x4787, x70125);
  nand n4885(x4885, x4786, x4887);
  nand n4886(x4886, x4885, x4884);
  nand n4888(x4888, x4787, x70139);
  nand n4889(x4889, x4786, x4891);
  nand n4890(x4890, x4889, x4888);
  nand n4892(x4892, x4787, x70153);
  nand n4893(x4893, x4786, x4895);
  nand n4894(x4894, x4893, x4892);
  nand n4896(x4896, x4787, x70167);
  nand n4897(x4897, x4786, x4899);
  nand n4898(x4898, x4897, x4896);
  nand n4900(x4900, x4787, x70181);
  nand n4901(x4901, x4786, x4903);
  nand n4902(x4902, x4901, x4900);
  nand n4904(x4904, x4787, x70195);
  nand n4905(x4905, x4786, x4907);
  nand n4906(x4906, x4905, x4904);
  nand n4908(x4908, x4787, x70209);
  nand n4909(x4909, x4786, x4911);
  nand n4910(x4910, x4909, x4908);
  nand n4912(x4912, x4787, x70223);
  nand n4913(x4913, x4786, x4915);
  nand n4914(x4914, x4913, x4912);
  nand n4916(x4916, x2305, x71073);
  nand n4918(x4918, x4917, x69789);
  nand n4919(x4919, x4916, x4921);
  nand n4920(x4920, x4919, x4918);
  nand n4922(x4922, x4917, x69803);
  nand n4923(x4923, x4916, x4925);
  nand n4924(x4924, x4923, x4922);
  nand n4926(x4926, x4917, x69817);
  nand n4927(x4927, x4916, x4929);
  nand n4928(x4928, x4927, x4926);
  nand n4930(x4930, x4917, x69831);
  nand n4931(x4931, x4916, x4933);
  nand n4932(x4932, x4931, x4930);
  nand n4934(x4934, x4917, x69845);
  nand n4935(x4935, x4916, x4937);
  nand n4936(x4936, x4935, x4934);
  nand n4938(x4938, x4917, x69859);
  nand n4939(x4939, x4916, x4941);
  nand n4940(x4940, x4939, x4938);
  nand n4942(x4942, x4917, x69873);
  nand n4943(x4943, x4916, x4945);
  nand n4944(x4944, x4943, x4942);
  nand n4946(x4946, x4917, x69887);
  nand n4947(x4947, x4916, x4949);
  nand n4948(x4948, x4947, x4946);
  nand n4950(x4950, x4917, x69901);
  nand n4951(x4951, x4916, x4953);
  nand n4952(x4952, x4951, x4950);
  nand n4954(x4954, x4917, x69915);
  nand n4955(x4955, x4916, x4957);
  nand n4956(x4956, x4955, x4954);
  nand n4958(x4958, x4917, x69929);
  nand n4959(x4959, x4916, x4961);
  nand n4960(x4960, x4959, x4958);
  nand n4962(x4962, x4917, x69943);
  nand n4963(x4963, x4916, x4965);
  nand n4964(x4964, x4963, x4962);
  nand n4966(x4966, x4917, x69957);
  nand n4967(x4967, x4916, x4969);
  nand n4968(x4968, x4967, x4966);
  nand n4970(x4970, x4917, x69971);
  nand n4971(x4971, x4916, x4973);
  nand n4972(x4972, x4971, x4970);
  nand n4974(x4974, x4917, x69985);
  nand n4975(x4975, x4916, x4977);
  nand n4976(x4976, x4975, x4974);
  nand n4978(x4978, x4917, x69999);
  nand n4979(x4979, x4916, x4981);
  nand n4980(x4980, x4979, x4978);
  nand n4982(x4982, x4917, x70013);
  nand n4983(x4983, x4916, x4985);
  nand n4984(x4984, x4983, x4982);
  nand n4986(x4986, x4917, x70027);
  nand n4987(x4987, x4916, x4989);
  nand n4988(x4988, x4987, x4986);
  nand n4990(x4990, x4917, x70041);
  nand n4991(x4991, x4916, x4993);
  nand n4992(x4992, x4991, x4990);
  nand n4994(x4994, x4917, x70055);
  nand n4995(x4995, x4916, x4997);
  nand n4996(x4996, x4995, x4994);
  nand n4998(x4998, x4917, x70069);
  nand n4999(x4999, x4916, x5001);
  nand n5000(x5000, x4999, x4998);
  nand n5002(x5002, x4917, x70083);
  nand n5003(x5003, x4916, x5005);
  nand n5004(x5004, x5003, x5002);
  nand n5006(x5006, x4917, x70097);
  nand n5007(x5007, x4916, x5009);
  nand n5008(x5008, x5007, x5006);
  nand n5010(x5010, x4917, x70111);
  nand n5011(x5011, x4916, x5013);
  nand n5012(x5012, x5011, x5010);
  nand n5014(x5014, x4917, x70125);
  nand n5015(x5015, x4916, x5017);
  nand n5016(x5016, x5015, x5014);
  nand n5018(x5018, x4917, x70139);
  nand n5019(x5019, x4916, x5021);
  nand n5020(x5020, x5019, x5018);
  nand n5022(x5022, x4917, x70153);
  nand n5023(x5023, x4916, x5025);
  nand n5024(x5024, x5023, x5022);
  nand n5026(x5026, x4917, x70167);
  nand n5027(x5027, x4916, x5029);
  nand n5028(x5028, x5027, x5026);
  nand n5030(x5030, x4917, x70181);
  nand n5031(x5031, x4916, x5033);
  nand n5032(x5032, x5031, x5030);
  nand n5034(x5034, x4917, x70195);
  nand n5035(x5035, x4916, x5037);
  nand n5036(x5036, x5035, x5034);
  nand n5038(x5038, x4917, x70209);
  nand n5039(x5039, x4916, x5041);
  nand n5040(x5040, x5039, x5038);
  nand n5042(x5042, x4917, x70223);
  nand n5043(x5043, x4916, x5045);
  nand n5044(x5044, x5043, x5042);
  nand n5046(x5046, x2307, x71073);
  nand n5048(x5048, x5047, x69789);
  nand n5049(x5049, x5046, x5051);
  nand n5050(x5050, x5049, x5048);
  nand n5052(x5052, x5047, x69803);
  nand n5053(x5053, x5046, x5055);
  nand n5054(x5054, x5053, x5052);
  nand n5056(x5056, x5047, x69817);
  nand n5057(x5057, x5046, x5059);
  nand n5058(x5058, x5057, x5056);
  nand n5060(x5060, x5047, x69831);
  nand n5061(x5061, x5046, x5063);
  nand n5062(x5062, x5061, x5060);
  nand n5064(x5064, x5047, x69845);
  nand n5065(x5065, x5046, x5067);
  nand n5066(x5066, x5065, x5064);
  nand n5068(x5068, x5047, x69859);
  nand n5069(x5069, x5046, x5071);
  nand n5070(x5070, x5069, x5068);
  nand n5072(x5072, x5047, x69873);
  nand n5073(x5073, x5046, x5075);
  nand n5074(x5074, x5073, x5072);
  nand n5076(x5076, x5047, x69887);
  nand n5077(x5077, x5046, x5079);
  nand n5078(x5078, x5077, x5076);
  nand n5080(x5080, x5047, x69901);
  nand n5081(x5081, x5046, x5083);
  nand n5082(x5082, x5081, x5080);
  nand n5084(x5084, x5047, x69915);
  nand n5085(x5085, x5046, x5087);
  nand n5086(x5086, x5085, x5084);
  nand n5088(x5088, x5047, x69929);
  nand n5089(x5089, x5046, x5091);
  nand n5090(x5090, x5089, x5088);
  nand n5092(x5092, x5047, x69943);
  nand n5093(x5093, x5046, x5095);
  nand n5094(x5094, x5093, x5092);
  nand n5096(x5096, x5047, x69957);
  nand n5097(x5097, x5046, x5099);
  nand n5098(x5098, x5097, x5096);
  nand n5100(x5100, x5047, x69971);
  nand n5101(x5101, x5046, x5103);
  nand n5102(x5102, x5101, x5100);
  nand n5104(x5104, x5047, x69985);
  nand n5105(x5105, x5046, x5107);
  nand n5106(x5106, x5105, x5104);
  nand n5108(x5108, x5047, x69999);
  nand n5109(x5109, x5046, x5111);
  nand n5110(x5110, x5109, x5108);
  nand n5112(x5112, x5047, x70013);
  nand n5113(x5113, x5046, x5115);
  nand n5114(x5114, x5113, x5112);
  nand n5116(x5116, x5047, x70027);
  nand n5117(x5117, x5046, x5119);
  nand n5118(x5118, x5117, x5116);
  nand n5120(x5120, x5047, x70041);
  nand n5121(x5121, x5046, x5123);
  nand n5122(x5122, x5121, x5120);
  nand n5124(x5124, x5047, x70055);
  nand n5125(x5125, x5046, x5127);
  nand n5126(x5126, x5125, x5124);
  nand n5128(x5128, x5047, x70069);
  nand n5129(x5129, x5046, x5131);
  nand n5130(x5130, x5129, x5128);
  nand n5132(x5132, x5047, x70083);
  nand n5133(x5133, x5046, x5135);
  nand n5134(x5134, x5133, x5132);
  nand n5136(x5136, x5047, x70097);
  nand n5137(x5137, x5046, x5139);
  nand n5138(x5138, x5137, x5136);
  nand n5140(x5140, x5047, x70111);
  nand n5141(x5141, x5046, x5143);
  nand n5142(x5142, x5141, x5140);
  nand n5144(x5144, x5047, x70125);
  nand n5145(x5145, x5046, x5147);
  nand n5146(x5146, x5145, x5144);
  nand n5148(x5148, x5047, x70139);
  nand n5149(x5149, x5046, x5151);
  nand n5150(x5150, x5149, x5148);
  nand n5152(x5152, x5047, x70153);
  nand n5153(x5153, x5046, x5155);
  nand n5154(x5154, x5153, x5152);
  nand n5156(x5156, x5047, x70167);
  nand n5157(x5157, x5046, x5159);
  nand n5158(x5158, x5157, x5156);
  nand n5160(x5160, x5047, x70181);
  nand n5161(x5161, x5046, x5163);
  nand n5162(x5162, x5161, x5160);
  nand n5164(x5164, x5047, x70195);
  nand n5165(x5165, x5046, x5167);
  nand n5166(x5166, x5165, x5164);
  nand n5168(x5168, x5047, x70209);
  nand n5169(x5169, x5046, x5171);
  nand n5170(x5170, x5169, x5168);
  nand n5172(x5172, x5047, x70223);
  nand n5173(x5173, x5046, x5175);
  nand n5174(x5174, x5173, x5172);
  nand n5176(x5176, x2309, x71073);
  nand n5178(x5178, x5177, x69789);
  nand n5179(x5179, x5176, x5181);
  nand n5180(x5180, x5179, x5178);
  nand n5182(x5182, x5177, x69803);
  nand n5183(x5183, x5176, x5185);
  nand n5184(x5184, x5183, x5182);
  nand n5186(x5186, x5177, x69817);
  nand n5187(x5187, x5176, x5189);
  nand n5188(x5188, x5187, x5186);
  nand n5190(x5190, x5177, x69831);
  nand n5191(x5191, x5176, x5193);
  nand n5192(x5192, x5191, x5190);
  nand n5194(x5194, x5177, x69845);
  nand n5195(x5195, x5176, x5197);
  nand n5196(x5196, x5195, x5194);
  nand n5198(x5198, x5177, x69859);
  nand n5199(x5199, x5176, x5201);
  nand n5200(x5200, x5199, x5198);
  nand n5202(x5202, x5177, x69873);
  nand n5203(x5203, x5176, x5205);
  nand n5204(x5204, x5203, x5202);
  nand n5206(x5206, x5177, x69887);
  nand n5207(x5207, x5176, x5209);
  nand n5208(x5208, x5207, x5206);
  nand n5210(x5210, x5177, x69901);
  nand n5211(x5211, x5176, x5213);
  nand n5212(x5212, x5211, x5210);
  nand n5214(x5214, x5177, x69915);
  nand n5215(x5215, x5176, x5217);
  nand n5216(x5216, x5215, x5214);
  nand n5218(x5218, x5177, x69929);
  nand n5219(x5219, x5176, x5221);
  nand n5220(x5220, x5219, x5218);
  nand n5222(x5222, x5177, x69943);
  nand n5223(x5223, x5176, x5225);
  nand n5224(x5224, x5223, x5222);
  nand n5226(x5226, x5177, x69957);
  nand n5227(x5227, x5176, x5229);
  nand n5228(x5228, x5227, x5226);
  nand n5230(x5230, x5177, x69971);
  nand n5231(x5231, x5176, x5233);
  nand n5232(x5232, x5231, x5230);
  nand n5234(x5234, x5177, x69985);
  nand n5235(x5235, x5176, x5237);
  nand n5236(x5236, x5235, x5234);
  nand n5238(x5238, x5177, x69999);
  nand n5239(x5239, x5176, x5241);
  nand n5240(x5240, x5239, x5238);
  nand n5242(x5242, x5177, x70013);
  nand n5243(x5243, x5176, x5245);
  nand n5244(x5244, x5243, x5242);
  nand n5246(x5246, x5177, x70027);
  nand n5247(x5247, x5176, x5249);
  nand n5248(x5248, x5247, x5246);
  nand n5250(x5250, x5177, x70041);
  nand n5251(x5251, x5176, x5253);
  nand n5252(x5252, x5251, x5250);
  nand n5254(x5254, x5177, x70055);
  nand n5255(x5255, x5176, x5257);
  nand n5256(x5256, x5255, x5254);
  nand n5258(x5258, x5177, x70069);
  nand n5259(x5259, x5176, x5261);
  nand n5260(x5260, x5259, x5258);
  nand n5262(x5262, x5177, x70083);
  nand n5263(x5263, x5176, x5265);
  nand n5264(x5264, x5263, x5262);
  nand n5266(x5266, x5177, x70097);
  nand n5267(x5267, x5176, x5269);
  nand n5268(x5268, x5267, x5266);
  nand n5270(x5270, x5177, x70111);
  nand n5271(x5271, x5176, x5273);
  nand n5272(x5272, x5271, x5270);
  nand n5274(x5274, x5177, x70125);
  nand n5275(x5275, x5176, x5277);
  nand n5276(x5276, x5275, x5274);
  nand n5278(x5278, x5177, x70139);
  nand n5279(x5279, x5176, x5281);
  nand n5280(x5280, x5279, x5278);
  nand n5282(x5282, x5177, x70153);
  nand n5283(x5283, x5176, x5285);
  nand n5284(x5284, x5283, x5282);
  nand n5286(x5286, x5177, x70167);
  nand n5287(x5287, x5176, x5289);
  nand n5288(x5288, x5287, x5286);
  nand n5290(x5290, x5177, x70181);
  nand n5291(x5291, x5176, x5293);
  nand n5292(x5292, x5291, x5290);
  nand n5294(x5294, x5177, x70195);
  nand n5295(x5295, x5176, x5297);
  nand n5296(x5296, x5295, x5294);
  nand n5298(x5298, x5177, x70209);
  nand n5299(x5299, x5176, x5301);
  nand n5300(x5300, x5299, x5298);
  nand n5302(x5302, x5177, x70223);
  nand n5303(x5303, x5176, x5305);
  nand n5304(x5304, x5303, x5302);
  nand n5306(x5306, x2311, x71073);
  nand n5308(x5308, x5307, x69789);
  nand n5309(x5309, x5306, x5311);
  nand n5310(x5310, x5309, x5308);
  nand n5312(x5312, x5307, x69803);
  nand n5313(x5313, x5306, x5315);
  nand n5314(x5314, x5313, x5312);
  nand n5316(x5316, x5307, x69817);
  nand n5317(x5317, x5306, x5319);
  nand n5318(x5318, x5317, x5316);
  nand n5320(x5320, x5307, x69831);
  nand n5321(x5321, x5306, x5323);
  nand n5322(x5322, x5321, x5320);
  nand n5324(x5324, x5307, x69845);
  nand n5325(x5325, x5306, x5327);
  nand n5326(x5326, x5325, x5324);
  nand n5328(x5328, x5307, x69859);
  nand n5329(x5329, x5306, x5331);
  nand n5330(x5330, x5329, x5328);
  nand n5332(x5332, x5307, x69873);
  nand n5333(x5333, x5306, x5335);
  nand n5334(x5334, x5333, x5332);
  nand n5336(x5336, x5307, x69887);
  nand n5337(x5337, x5306, x5339);
  nand n5338(x5338, x5337, x5336);
  nand n5340(x5340, x5307, x69901);
  nand n5341(x5341, x5306, x5343);
  nand n5342(x5342, x5341, x5340);
  nand n5344(x5344, x5307, x69915);
  nand n5345(x5345, x5306, x5347);
  nand n5346(x5346, x5345, x5344);
  nand n5348(x5348, x5307, x69929);
  nand n5349(x5349, x5306, x5351);
  nand n5350(x5350, x5349, x5348);
  nand n5352(x5352, x5307, x69943);
  nand n5353(x5353, x5306, x5355);
  nand n5354(x5354, x5353, x5352);
  nand n5356(x5356, x5307, x69957);
  nand n5357(x5357, x5306, x5359);
  nand n5358(x5358, x5357, x5356);
  nand n5360(x5360, x5307, x69971);
  nand n5361(x5361, x5306, x5363);
  nand n5362(x5362, x5361, x5360);
  nand n5364(x5364, x5307, x69985);
  nand n5365(x5365, x5306, x5367);
  nand n5366(x5366, x5365, x5364);
  nand n5368(x5368, x5307, x69999);
  nand n5369(x5369, x5306, x5371);
  nand n5370(x5370, x5369, x5368);
  nand n5372(x5372, x5307, x70013);
  nand n5373(x5373, x5306, x5375);
  nand n5374(x5374, x5373, x5372);
  nand n5376(x5376, x5307, x70027);
  nand n5377(x5377, x5306, x5379);
  nand n5378(x5378, x5377, x5376);
  nand n5380(x5380, x5307, x70041);
  nand n5381(x5381, x5306, x5383);
  nand n5382(x5382, x5381, x5380);
  nand n5384(x5384, x5307, x70055);
  nand n5385(x5385, x5306, x5387);
  nand n5386(x5386, x5385, x5384);
  nand n5388(x5388, x5307, x70069);
  nand n5389(x5389, x5306, x5391);
  nand n5390(x5390, x5389, x5388);
  nand n5392(x5392, x5307, x70083);
  nand n5393(x5393, x5306, x5395);
  nand n5394(x5394, x5393, x5392);
  nand n5396(x5396, x5307, x70097);
  nand n5397(x5397, x5306, x5399);
  nand n5398(x5398, x5397, x5396);
  nand n5400(x5400, x5307, x70111);
  nand n5401(x5401, x5306, x5403);
  nand n5402(x5402, x5401, x5400);
  nand n5404(x5404, x5307, x70125);
  nand n5405(x5405, x5306, x5407);
  nand n5406(x5406, x5405, x5404);
  nand n5408(x5408, x5307, x70139);
  nand n5409(x5409, x5306, x5411);
  nand n5410(x5410, x5409, x5408);
  nand n5412(x5412, x5307, x70153);
  nand n5413(x5413, x5306, x5415);
  nand n5414(x5414, x5413, x5412);
  nand n5416(x5416, x5307, x70167);
  nand n5417(x5417, x5306, x5419);
  nand n5418(x5418, x5417, x5416);
  nand n5420(x5420, x5307, x70181);
  nand n5421(x5421, x5306, x5423);
  nand n5422(x5422, x5421, x5420);
  nand n5424(x5424, x5307, x70195);
  nand n5425(x5425, x5306, x5427);
  nand n5426(x5426, x5425, x5424);
  nand n5428(x5428, x5307, x70209);
  nand n5429(x5429, x5306, x5431);
  nand n5430(x5430, x5429, x5428);
  nand n5432(x5432, x5307, x70223);
  nand n5433(x5433, x5306, x5435);
  nand n5434(x5434, x5433, x5432);
  nand n5436(x5436, x2297, x71075);
  nand n5438(x5438, x5437, x70239);
  nand n5439(x5439, x5436, x5443);
  nand n5440(x5440, x5439, x5438);
  nand n5444(x5444, x5437, x70253);
  nand n5445(x5445, x5436, x5449);
  nand n5446(x5446, x5445, x5444);
  nand n5450(x5450, x5437, x70267);
  nand n5451(x5451, x5436, x5453);
  nand n5452(x5452, x5451, x5450);
  nand n5454(x5454, x5437, x70281);
  nand n5455(x5455, x5436, x5457);
  nand n5456(x5456, x5455, x5454);
  nand n5458(x5458, x5437, x70295);
  nand n5459(x5459, x5436, x5461);
  nand n5460(x5460, x5459, x5458);
  nand n5462(x5462, x5437, x70309);
  nand n5463(x5463, x5436, x5465);
  nand n5464(x5464, x5463, x5462);
  nand n5466(x5466, x5437, x70323);
  nand n5467(x5467, x5436, x5469);
  nand n5468(x5468, x5467, x5466);
  nand n5470(x5470, x5437, x70337);
  nand n5471(x5471, x5436, x5473);
  nand n5472(x5472, x5471, x5470);
  nand n5474(x5474, x5437, x70351);
  nand n5475(x5475, x5436, x5477);
  nand n5476(x5476, x5475, x5474);
  nand n5478(x5478, x5437, x70365);
  nand n5479(x5479, x5436, x5481);
  nand n5480(x5480, x5479, x5478);
  nand n5482(x5482, x5437, x70379);
  nand n5483(x5483, x5436, x5485);
  nand n5484(x5484, x5483, x5482);
  nand n5486(x5486, x5437, x70393);
  nand n5487(x5487, x5436, x5489);
  nand n5488(x5488, x5487, x5486);
  nand n5490(x5490, x5437, x70407);
  nand n5491(x5491, x5436, x5493);
  nand n5492(x5492, x5491, x5490);
  nand n5494(x5494, x5437, x70421);
  nand n5495(x5495, x5436, x5497);
  nand n5496(x5496, x5495, x5494);
  nand n5498(x5498, x5437, x70435);
  nand n5499(x5499, x5436, x5501);
  nand n5500(x5500, x5499, x5498);
  nand n5502(x5502, x5437, x70449);
  nand n5503(x5503, x5436, x5505);
  nand n5504(x5504, x5503, x5502);
  nand n5506(x5506, x5437, x70463);
  nand n5507(x5507, x5436, x5509);
  nand n5508(x5508, x5507, x5506);
  nand n5510(x5510, x5437, x70477);
  nand n5511(x5511, x5436, x5513);
  nand n5512(x5512, x5511, x5510);
  nand n5514(x5514, x5437, x70491);
  nand n5515(x5515, x5436, x5517);
  nand n5516(x5516, x5515, x5514);
  nand n5518(x5518, x5437, x70505);
  nand n5519(x5519, x5436, x5521);
  nand n5520(x5520, x5519, x5518);
  nand n5522(x5522, x5437, x70519);
  nand n5523(x5523, x5436, x5525);
  nand n5524(x5524, x5523, x5522);
  nand n5526(x5526, x5437, x70533);
  nand n5527(x5527, x5436, x5529);
  nand n5528(x5528, x5527, x5526);
  nand n5530(x5530, x5437, x70547);
  nand n5531(x5531, x5436, x5533);
  nand n5532(x5532, x5531, x5530);
  nand n5534(x5534, x5437, x70561);
  nand n5535(x5535, x5436, x5537);
  nand n5536(x5536, x5535, x5534);
  nand n5538(x5538, x5437, x70575);
  nand n5539(x5539, x5436, x5541);
  nand n5540(x5540, x5539, x5538);
  nand n5542(x5542, x5437, x70589);
  nand n5543(x5543, x5436, x5545);
  nand n5544(x5544, x5543, x5542);
  nand n5546(x5546, x5437, x70603);
  nand n5547(x5547, x5436, x5549);
  nand n5548(x5548, x5547, x5546);
  nand n5550(x5550, x5437, x70617);
  nand n5551(x5551, x5436, x5553);
  nand n5552(x5552, x5551, x5550);
  nand n5554(x5554, x5437, x70631);
  nand n5555(x5555, x5436, x5557);
  nand n5556(x5556, x5555, x5554);
  nand n5558(x5558, x5437, x70645);
  nand n5559(x5559, x5436, x5561);
  nand n5560(x5560, x5559, x5558);
  nand n5562(x5562, x5437, x70659);
  nand n5563(x5563, x5436, x5565);
  nand n5564(x5564, x5563, x5562);
  nand n5566(x5566, x5437, x70673);
  nand n5567(x5567, x5436, x5569);
  nand n5568(x5568, x5567, x5566);
  nand n5570(x5570, x2299, x71075);
  nand n5572(x5572, x5571, x70239);
  nand n5573(x5573, x5570, x5575);
  nand n5574(x5574, x5573, x5572);
  nand n5576(x5576, x5571, x70253);
  nand n5577(x5577, x5570, x5579);
  nand n5578(x5578, x5577, x5576);
  nand n5580(x5580, x5571, x70267);
  nand n5581(x5581, x5570, x5583);
  nand n5582(x5582, x5581, x5580);
  nand n5584(x5584, x5571, x70281);
  nand n5585(x5585, x5570, x5587);
  nand n5586(x5586, x5585, x5584);
  nand n5588(x5588, x5571, x70295);
  nand n5589(x5589, x5570, x5591);
  nand n5590(x5590, x5589, x5588);
  nand n5592(x5592, x5571, x70309);
  nand n5593(x5593, x5570, x5595);
  nand n5594(x5594, x5593, x5592);
  nand n5596(x5596, x5571, x70323);
  nand n5597(x5597, x5570, x5599);
  nand n5598(x5598, x5597, x5596);
  nand n5600(x5600, x5571, x70337);
  nand n5601(x5601, x5570, x5603);
  nand n5602(x5602, x5601, x5600);
  nand n5604(x5604, x5571, x70351);
  nand n5605(x5605, x5570, x5607);
  nand n5606(x5606, x5605, x5604);
  nand n5608(x5608, x5571, x70365);
  nand n5609(x5609, x5570, x5611);
  nand n5610(x5610, x5609, x5608);
  nand n5612(x5612, x5571, x70379);
  nand n5613(x5613, x5570, x5615);
  nand n5614(x5614, x5613, x5612);
  nand n5616(x5616, x5571, x70393);
  nand n5617(x5617, x5570, x5619);
  nand n5618(x5618, x5617, x5616);
  nand n5620(x5620, x5571, x70407);
  nand n5621(x5621, x5570, x5623);
  nand n5622(x5622, x5621, x5620);
  nand n5624(x5624, x5571, x70421);
  nand n5625(x5625, x5570, x5627);
  nand n5626(x5626, x5625, x5624);
  nand n5628(x5628, x5571, x70435);
  nand n5629(x5629, x5570, x5631);
  nand n5630(x5630, x5629, x5628);
  nand n5632(x5632, x5571, x70449);
  nand n5633(x5633, x5570, x5635);
  nand n5634(x5634, x5633, x5632);
  nand n5636(x5636, x5571, x70463);
  nand n5637(x5637, x5570, x5639);
  nand n5638(x5638, x5637, x5636);
  nand n5640(x5640, x5571, x70477);
  nand n5641(x5641, x5570, x5643);
  nand n5642(x5642, x5641, x5640);
  nand n5644(x5644, x5571, x70491);
  nand n5645(x5645, x5570, x5647);
  nand n5646(x5646, x5645, x5644);
  nand n5648(x5648, x5571, x70505);
  nand n5649(x5649, x5570, x5651);
  nand n5650(x5650, x5649, x5648);
  nand n5652(x5652, x5571, x70519);
  nand n5653(x5653, x5570, x5655);
  nand n5654(x5654, x5653, x5652);
  nand n5656(x5656, x5571, x70533);
  nand n5657(x5657, x5570, x5659);
  nand n5658(x5658, x5657, x5656);
  nand n5660(x5660, x5571, x70547);
  nand n5661(x5661, x5570, x5663);
  nand n5662(x5662, x5661, x5660);
  nand n5664(x5664, x5571, x70561);
  nand n5665(x5665, x5570, x5667);
  nand n5666(x5666, x5665, x5664);
  nand n5668(x5668, x5571, x70575);
  nand n5669(x5669, x5570, x5671);
  nand n5670(x5670, x5669, x5668);
  nand n5672(x5672, x5571, x70589);
  nand n5673(x5673, x5570, x5675);
  nand n5674(x5674, x5673, x5672);
  nand n5676(x5676, x5571, x70603);
  nand n5677(x5677, x5570, x5679);
  nand n5678(x5678, x5677, x5676);
  nand n5680(x5680, x5571, x70617);
  nand n5681(x5681, x5570, x5683);
  nand n5682(x5682, x5681, x5680);
  nand n5684(x5684, x5571, x70631);
  nand n5685(x5685, x5570, x5687);
  nand n5686(x5686, x5685, x5684);
  nand n5688(x5688, x5571, x70645);
  nand n5689(x5689, x5570, x5691);
  nand n5690(x5690, x5689, x5688);
  nand n5692(x5692, x5571, x70659);
  nand n5693(x5693, x5570, x5695);
  nand n5694(x5694, x5693, x5692);
  nand n5696(x5696, x5571, x70673);
  nand n5697(x5697, x5570, x5699);
  nand n5698(x5698, x5697, x5696);
  nand n5700(x5700, x2301, x71075);
  nand n5702(x5702, x5701, x70239);
  nand n5703(x5703, x5700, x5705);
  nand n5704(x5704, x5703, x5702);
  nand n5706(x5706, x5701, x70253);
  nand n5707(x5707, x5700, x5709);
  nand n5708(x5708, x5707, x5706);
  nand n5710(x5710, x5701, x70267);
  nand n5711(x5711, x5700, x5713);
  nand n5712(x5712, x5711, x5710);
  nand n5714(x5714, x5701, x70281);
  nand n5715(x5715, x5700, x5717);
  nand n5716(x5716, x5715, x5714);
  nand n5718(x5718, x5701, x70295);
  nand n5719(x5719, x5700, x5721);
  nand n5720(x5720, x5719, x5718);
  nand n5722(x5722, x5701, x70309);
  nand n5723(x5723, x5700, x5725);
  nand n5724(x5724, x5723, x5722);
  nand n5726(x5726, x5701, x70323);
  nand n5727(x5727, x5700, x5729);
  nand n5728(x5728, x5727, x5726);
  nand n5730(x5730, x5701, x70337);
  nand n5731(x5731, x5700, x5733);
  nand n5732(x5732, x5731, x5730);
  nand n5734(x5734, x5701, x70351);
  nand n5735(x5735, x5700, x5737);
  nand n5736(x5736, x5735, x5734);
  nand n5738(x5738, x5701, x70365);
  nand n5739(x5739, x5700, x5741);
  nand n5740(x5740, x5739, x5738);
  nand n5742(x5742, x5701, x70379);
  nand n5743(x5743, x5700, x5745);
  nand n5744(x5744, x5743, x5742);
  nand n5746(x5746, x5701, x70393);
  nand n5747(x5747, x5700, x5749);
  nand n5748(x5748, x5747, x5746);
  nand n5750(x5750, x5701, x70407);
  nand n5751(x5751, x5700, x5753);
  nand n5752(x5752, x5751, x5750);
  nand n5754(x5754, x5701, x70421);
  nand n5755(x5755, x5700, x5757);
  nand n5756(x5756, x5755, x5754);
  nand n5758(x5758, x5701, x70435);
  nand n5759(x5759, x5700, x5761);
  nand n5760(x5760, x5759, x5758);
  nand n5762(x5762, x5701, x70449);
  nand n5763(x5763, x5700, x5765);
  nand n5764(x5764, x5763, x5762);
  nand n5766(x5766, x5701, x70463);
  nand n5767(x5767, x5700, x5769);
  nand n5768(x5768, x5767, x5766);
  nand n5770(x5770, x5701, x70477);
  nand n5771(x5771, x5700, x5773);
  nand n5772(x5772, x5771, x5770);
  nand n5774(x5774, x5701, x70491);
  nand n5775(x5775, x5700, x5777);
  nand n5776(x5776, x5775, x5774);
  nand n5778(x5778, x5701, x70505);
  nand n5779(x5779, x5700, x5781);
  nand n5780(x5780, x5779, x5778);
  nand n5782(x5782, x5701, x70519);
  nand n5783(x5783, x5700, x5785);
  nand n5784(x5784, x5783, x5782);
  nand n5786(x5786, x5701, x70533);
  nand n5787(x5787, x5700, x5789);
  nand n5788(x5788, x5787, x5786);
  nand n5790(x5790, x5701, x70547);
  nand n5791(x5791, x5700, x5793);
  nand n5792(x5792, x5791, x5790);
  nand n5794(x5794, x5701, x70561);
  nand n5795(x5795, x5700, x5797);
  nand n5796(x5796, x5795, x5794);
  nand n5798(x5798, x5701, x70575);
  nand n5799(x5799, x5700, x5801);
  nand n5800(x5800, x5799, x5798);
  nand n5802(x5802, x5701, x70589);
  nand n5803(x5803, x5700, x5805);
  nand n5804(x5804, x5803, x5802);
  nand n5806(x5806, x5701, x70603);
  nand n5807(x5807, x5700, x5809);
  nand n5808(x5808, x5807, x5806);
  nand n5810(x5810, x5701, x70617);
  nand n5811(x5811, x5700, x5813);
  nand n5812(x5812, x5811, x5810);
  nand n5814(x5814, x5701, x70631);
  nand n5815(x5815, x5700, x5817);
  nand n5816(x5816, x5815, x5814);
  nand n5818(x5818, x5701, x70645);
  nand n5819(x5819, x5700, x5821);
  nand n5820(x5820, x5819, x5818);
  nand n5822(x5822, x5701, x70659);
  nand n5823(x5823, x5700, x5825);
  nand n5824(x5824, x5823, x5822);
  nand n5826(x5826, x5701, x70673);
  nand n5827(x5827, x5700, x5829);
  nand n5828(x5828, x5827, x5826);
  nand n5830(x5830, x2303, x71075);
  nand n5832(x5832, x5831, x70239);
  nand n5833(x5833, x5830, x5835);
  nand n5834(x5834, x5833, x5832);
  nand n5836(x5836, x5831, x70253);
  nand n5837(x5837, x5830, x5839);
  nand n5838(x5838, x5837, x5836);
  nand n5840(x5840, x5831, x70267);
  nand n5841(x5841, x5830, x5843);
  nand n5842(x5842, x5841, x5840);
  nand n5844(x5844, x5831, x70281);
  nand n5845(x5845, x5830, x5847);
  nand n5846(x5846, x5845, x5844);
  nand n5848(x5848, x5831, x70295);
  nand n5849(x5849, x5830, x5851);
  nand n5850(x5850, x5849, x5848);
  nand n5852(x5852, x5831, x70309);
  nand n5853(x5853, x5830, x5855);
  nand n5854(x5854, x5853, x5852);
  nand n5856(x5856, x5831, x70323);
  nand n5857(x5857, x5830, x5859);
  nand n5858(x5858, x5857, x5856);
  nand n5860(x5860, x5831, x70337);
  nand n5861(x5861, x5830, x5863);
  nand n5862(x5862, x5861, x5860);
  nand n5864(x5864, x5831, x70351);
  nand n5865(x5865, x5830, x5867);
  nand n5866(x5866, x5865, x5864);
  nand n5868(x5868, x5831, x70365);
  nand n5869(x5869, x5830, x5871);
  nand n5870(x5870, x5869, x5868);
  nand n5872(x5872, x5831, x70379);
  nand n5873(x5873, x5830, x5875);
  nand n5874(x5874, x5873, x5872);
  nand n5876(x5876, x5831, x70393);
  nand n5877(x5877, x5830, x5879);
  nand n5878(x5878, x5877, x5876);
  nand n5880(x5880, x5831, x70407);
  nand n5881(x5881, x5830, x5883);
  nand n5882(x5882, x5881, x5880);
  nand n5884(x5884, x5831, x70421);
  nand n5885(x5885, x5830, x5887);
  nand n5886(x5886, x5885, x5884);
  nand n5888(x5888, x5831, x70435);
  nand n5889(x5889, x5830, x5891);
  nand n5890(x5890, x5889, x5888);
  nand n5892(x5892, x5831, x70449);
  nand n5893(x5893, x5830, x5895);
  nand n5894(x5894, x5893, x5892);
  nand n5896(x5896, x5831, x70463);
  nand n5897(x5897, x5830, x5899);
  nand n5898(x5898, x5897, x5896);
  nand n5900(x5900, x5831, x70477);
  nand n5901(x5901, x5830, x5903);
  nand n5902(x5902, x5901, x5900);
  nand n5904(x5904, x5831, x70491);
  nand n5905(x5905, x5830, x5907);
  nand n5906(x5906, x5905, x5904);
  nand n5908(x5908, x5831, x70505);
  nand n5909(x5909, x5830, x5911);
  nand n5910(x5910, x5909, x5908);
  nand n5912(x5912, x5831, x70519);
  nand n5913(x5913, x5830, x5915);
  nand n5914(x5914, x5913, x5912);
  nand n5916(x5916, x5831, x70533);
  nand n5917(x5917, x5830, x5919);
  nand n5918(x5918, x5917, x5916);
  nand n5920(x5920, x5831, x70547);
  nand n5921(x5921, x5830, x5923);
  nand n5922(x5922, x5921, x5920);
  nand n5924(x5924, x5831, x70561);
  nand n5925(x5925, x5830, x5927);
  nand n5926(x5926, x5925, x5924);
  nand n5928(x5928, x5831, x70575);
  nand n5929(x5929, x5830, x5931);
  nand n5930(x5930, x5929, x5928);
  nand n5932(x5932, x5831, x70589);
  nand n5933(x5933, x5830, x5935);
  nand n5934(x5934, x5933, x5932);
  nand n5936(x5936, x5831, x70603);
  nand n5937(x5937, x5830, x5939);
  nand n5938(x5938, x5937, x5936);
  nand n5940(x5940, x5831, x70617);
  nand n5941(x5941, x5830, x5943);
  nand n5942(x5942, x5941, x5940);
  nand n5944(x5944, x5831, x70631);
  nand n5945(x5945, x5830, x5947);
  nand n5946(x5946, x5945, x5944);
  nand n5948(x5948, x5831, x70645);
  nand n5949(x5949, x5830, x5951);
  nand n5950(x5950, x5949, x5948);
  nand n5952(x5952, x5831, x70659);
  nand n5953(x5953, x5830, x5955);
  nand n5954(x5954, x5953, x5952);
  nand n5956(x5956, x5831, x70673);
  nand n5957(x5957, x5830, x5959);
  nand n5958(x5958, x5957, x5956);
  nand n5960(x5960, x2305, x71075);
  nand n5962(x5962, x5961, x70239);
  nand n5963(x5963, x5960, x5965);
  nand n5964(x5964, x5963, x5962);
  nand n5966(x5966, x5961, x70253);
  nand n5967(x5967, x5960, x5969);
  nand n5968(x5968, x5967, x5966);
  nand n5970(x5970, x5961, x70267);
  nand n5971(x5971, x5960, x5973);
  nand n5972(x5972, x5971, x5970);
  nand n5974(x5974, x5961, x70281);
  nand n5975(x5975, x5960, x5977);
  nand n5976(x5976, x5975, x5974);
  nand n5978(x5978, x5961, x70295);
  nand n5979(x5979, x5960, x5981);
  nand n5980(x5980, x5979, x5978);
  nand n5982(x5982, x5961, x70309);
  nand n5983(x5983, x5960, x5985);
  nand n5984(x5984, x5983, x5982);
  nand n5986(x5986, x5961, x70323);
  nand n5987(x5987, x5960, x5989);
  nand n5988(x5988, x5987, x5986);
  nand n5990(x5990, x5961, x70337);
  nand n5991(x5991, x5960, x5993);
  nand n5992(x5992, x5991, x5990);
  nand n5994(x5994, x5961, x70351);
  nand n5995(x5995, x5960, x5997);
  nand n5996(x5996, x5995, x5994);
  nand n5998(x5998, x5961, x70365);
  nand n5999(x5999, x5960, x6001);
  nand n6000(x6000, x5999, x5998);
  nand n6002(x6002, x5961, x70379);
  nand n6003(x6003, x5960, x6005);
  nand n6004(x6004, x6003, x6002);
  nand n6006(x6006, x5961, x70393);
  nand n6007(x6007, x5960, x6009);
  nand n6008(x6008, x6007, x6006);
  nand n6010(x6010, x5961, x70407);
  nand n6011(x6011, x5960, x6013);
  nand n6012(x6012, x6011, x6010);
  nand n6014(x6014, x5961, x70421);
  nand n6015(x6015, x5960, x6017);
  nand n6016(x6016, x6015, x6014);
  nand n6018(x6018, x5961, x70435);
  nand n6019(x6019, x5960, x6021);
  nand n6020(x6020, x6019, x6018);
  nand n6022(x6022, x5961, x70449);
  nand n6023(x6023, x5960, x6025);
  nand n6024(x6024, x6023, x6022);
  nand n6026(x6026, x5961, x70463);
  nand n6027(x6027, x5960, x6029);
  nand n6028(x6028, x6027, x6026);
  nand n6030(x6030, x5961, x70477);
  nand n6031(x6031, x5960, x6033);
  nand n6032(x6032, x6031, x6030);
  nand n6034(x6034, x5961, x70491);
  nand n6035(x6035, x5960, x6037);
  nand n6036(x6036, x6035, x6034);
  nand n6038(x6038, x5961, x70505);
  nand n6039(x6039, x5960, x6041);
  nand n6040(x6040, x6039, x6038);
  nand n6042(x6042, x5961, x70519);
  nand n6043(x6043, x5960, x6045);
  nand n6044(x6044, x6043, x6042);
  nand n6046(x6046, x5961, x70533);
  nand n6047(x6047, x5960, x6049);
  nand n6048(x6048, x6047, x6046);
  nand n6050(x6050, x5961, x70547);
  nand n6051(x6051, x5960, x6053);
  nand n6052(x6052, x6051, x6050);
  nand n6054(x6054, x5961, x70561);
  nand n6055(x6055, x5960, x6057);
  nand n6056(x6056, x6055, x6054);
  nand n6058(x6058, x5961, x70575);
  nand n6059(x6059, x5960, x6061);
  nand n6060(x6060, x6059, x6058);
  nand n6062(x6062, x5961, x70589);
  nand n6063(x6063, x5960, x6065);
  nand n6064(x6064, x6063, x6062);
  nand n6066(x6066, x5961, x70603);
  nand n6067(x6067, x5960, x6069);
  nand n6068(x6068, x6067, x6066);
  nand n6070(x6070, x5961, x70617);
  nand n6071(x6071, x5960, x6073);
  nand n6072(x6072, x6071, x6070);
  nand n6074(x6074, x5961, x70631);
  nand n6075(x6075, x5960, x6077);
  nand n6076(x6076, x6075, x6074);
  nand n6078(x6078, x5961, x70645);
  nand n6079(x6079, x5960, x6081);
  nand n6080(x6080, x6079, x6078);
  nand n6082(x6082, x5961, x70659);
  nand n6083(x6083, x5960, x6085);
  nand n6084(x6084, x6083, x6082);
  nand n6086(x6086, x5961, x70673);
  nand n6087(x6087, x5960, x6089);
  nand n6088(x6088, x6087, x6086);
  nand n6090(x6090, x2307, x71075);
  nand n6092(x6092, x6091, x70239);
  nand n6093(x6093, x6090, x6095);
  nand n6094(x6094, x6093, x6092);
  nand n6096(x6096, x6091, x70253);
  nand n6097(x6097, x6090, x6099);
  nand n6098(x6098, x6097, x6096);
  nand n6100(x6100, x6091, x70267);
  nand n6101(x6101, x6090, x6103);
  nand n6102(x6102, x6101, x6100);
  nand n6104(x6104, x6091, x70281);
  nand n6105(x6105, x6090, x6107);
  nand n6106(x6106, x6105, x6104);
  nand n6108(x6108, x6091, x70295);
  nand n6109(x6109, x6090, x6111);
  nand n6110(x6110, x6109, x6108);
  nand n6112(x6112, x6091, x70309);
  nand n6113(x6113, x6090, x6115);
  nand n6114(x6114, x6113, x6112);
  nand n6116(x6116, x6091, x70323);
  nand n6117(x6117, x6090, x6119);
  nand n6118(x6118, x6117, x6116);
  nand n6120(x6120, x6091, x70337);
  nand n6121(x6121, x6090, x6123);
  nand n6122(x6122, x6121, x6120);
  nand n6124(x6124, x6091, x70351);
  nand n6125(x6125, x6090, x6127);
  nand n6126(x6126, x6125, x6124);
  nand n6128(x6128, x6091, x70365);
  nand n6129(x6129, x6090, x6131);
  nand n6130(x6130, x6129, x6128);
  nand n6132(x6132, x6091, x70379);
  nand n6133(x6133, x6090, x6135);
  nand n6134(x6134, x6133, x6132);
  nand n6136(x6136, x6091, x70393);
  nand n6137(x6137, x6090, x6139);
  nand n6138(x6138, x6137, x6136);
  nand n6140(x6140, x6091, x70407);
  nand n6141(x6141, x6090, x6143);
  nand n6142(x6142, x6141, x6140);
  nand n6144(x6144, x6091, x70421);
  nand n6145(x6145, x6090, x6147);
  nand n6146(x6146, x6145, x6144);
  nand n6148(x6148, x6091, x70435);
  nand n6149(x6149, x6090, x6151);
  nand n6150(x6150, x6149, x6148);
  nand n6152(x6152, x6091, x70449);
  nand n6153(x6153, x6090, x6155);
  nand n6154(x6154, x6153, x6152);
  nand n6156(x6156, x6091, x70463);
  nand n6157(x6157, x6090, x6159);
  nand n6158(x6158, x6157, x6156);
  nand n6160(x6160, x6091, x70477);
  nand n6161(x6161, x6090, x6163);
  nand n6162(x6162, x6161, x6160);
  nand n6164(x6164, x6091, x70491);
  nand n6165(x6165, x6090, x6167);
  nand n6166(x6166, x6165, x6164);
  nand n6168(x6168, x6091, x70505);
  nand n6169(x6169, x6090, x6171);
  nand n6170(x6170, x6169, x6168);
  nand n6172(x6172, x6091, x70519);
  nand n6173(x6173, x6090, x6175);
  nand n6174(x6174, x6173, x6172);
  nand n6176(x6176, x6091, x70533);
  nand n6177(x6177, x6090, x6179);
  nand n6178(x6178, x6177, x6176);
  nand n6180(x6180, x6091, x70547);
  nand n6181(x6181, x6090, x6183);
  nand n6182(x6182, x6181, x6180);
  nand n6184(x6184, x6091, x70561);
  nand n6185(x6185, x6090, x6187);
  nand n6186(x6186, x6185, x6184);
  nand n6188(x6188, x6091, x70575);
  nand n6189(x6189, x6090, x6191);
  nand n6190(x6190, x6189, x6188);
  nand n6192(x6192, x6091, x70589);
  nand n6193(x6193, x6090, x6195);
  nand n6194(x6194, x6193, x6192);
  nand n6196(x6196, x6091, x70603);
  nand n6197(x6197, x6090, x6199);
  nand n6198(x6198, x6197, x6196);
  nand n6200(x6200, x6091, x70617);
  nand n6201(x6201, x6090, x6203);
  nand n6202(x6202, x6201, x6200);
  nand n6204(x6204, x6091, x70631);
  nand n6205(x6205, x6090, x6207);
  nand n6206(x6206, x6205, x6204);
  nand n6208(x6208, x6091, x70645);
  nand n6209(x6209, x6090, x6211);
  nand n6210(x6210, x6209, x6208);
  nand n6212(x6212, x6091, x70659);
  nand n6213(x6213, x6090, x6215);
  nand n6214(x6214, x6213, x6212);
  nand n6216(x6216, x6091, x70673);
  nand n6217(x6217, x6090, x6219);
  nand n6218(x6218, x6217, x6216);
  nand n6220(x6220, x2309, x71075);
  nand n6222(x6222, x6221, x70239);
  nand n6223(x6223, x6220, x6225);
  nand n6224(x6224, x6223, x6222);
  nand n6226(x6226, x6221, x70253);
  nand n6227(x6227, x6220, x6229);
  nand n6228(x6228, x6227, x6226);
  nand n6230(x6230, x6221, x70267);
  nand n6231(x6231, x6220, x6233);
  nand n6232(x6232, x6231, x6230);
  nand n6234(x6234, x6221, x70281);
  nand n6235(x6235, x6220, x6237);
  nand n6236(x6236, x6235, x6234);
  nand n6238(x6238, x6221, x70295);
  nand n6239(x6239, x6220, x6241);
  nand n6240(x6240, x6239, x6238);
  nand n6242(x6242, x6221, x70309);
  nand n6243(x6243, x6220, x6245);
  nand n6244(x6244, x6243, x6242);
  nand n6246(x6246, x6221, x70323);
  nand n6247(x6247, x6220, x6249);
  nand n6248(x6248, x6247, x6246);
  nand n6250(x6250, x6221, x70337);
  nand n6251(x6251, x6220, x6253);
  nand n6252(x6252, x6251, x6250);
  nand n6254(x6254, x6221, x70351);
  nand n6255(x6255, x6220, x6257);
  nand n6256(x6256, x6255, x6254);
  nand n6258(x6258, x6221, x70365);
  nand n6259(x6259, x6220, x6261);
  nand n6260(x6260, x6259, x6258);
  nand n6262(x6262, x6221, x70379);
  nand n6263(x6263, x6220, x6265);
  nand n6264(x6264, x6263, x6262);
  nand n6266(x6266, x6221, x70393);
  nand n6267(x6267, x6220, x6269);
  nand n6268(x6268, x6267, x6266);
  nand n6270(x6270, x6221, x70407);
  nand n6271(x6271, x6220, x6273);
  nand n6272(x6272, x6271, x6270);
  nand n6274(x6274, x6221, x70421);
  nand n6275(x6275, x6220, x6277);
  nand n6276(x6276, x6275, x6274);
  nand n6278(x6278, x6221, x70435);
  nand n6279(x6279, x6220, x6281);
  nand n6280(x6280, x6279, x6278);
  nand n6282(x6282, x6221, x70449);
  nand n6283(x6283, x6220, x6285);
  nand n6284(x6284, x6283, x6282);
  nand n6286(x6286, x6221, x70463);
  nand n6287(x6287, x6220, x6289);
  nand n6288(x6288, x6287, x6286);
  nand n6290(x6290, x6221, x70477);
  nand n6291(x6291, x6220, x6293);
  nand n6292(x6292, x6291, x6290);
  nand n6294(x6294, x6221, x70491);
  nand n6295(x6295, x6220, x6297);
  nand n6296(x6296, x6295, x6294);
  nand n6298(x6298, x6221, x70505);
  nand n6299(x6299, x6220, x6301);
  nand n6300(x6300, x6299, x6298);
  nand n6302(x6302, x6221, x70519);
  nand n6303(x6303, x6220, x6305);
  nand n6304(x6304, x6303, x6302);
  nand n6306(x6306, x6221, x70533);
  nand n6307(x6307, x6220, x6309);
  nand n6308(x6308, x6307, x6306);
  nand n6310(x6310, x6221, x70547);
  nand n6311(x6311, x6220, x6313);
  nand n6312(x6312, x6311, x6310);
  nand n6314(x6314, x6221, x70561);
  nand n6315(x6315, x6220, x6317);
  nand n6316(x6316, x6315, x6314);
  nand n6318(x6318, x6221, x70575);
  nand n6319(x6319, x6220, x6321);
  nand n6320(x6320, x6319, x6318);
  nand n6322(x6322, x6221, x70589);
  nand n6323(x6323, x6220, x6325);
  nand n6324(x6324, x6323, x6322);
  nand n6326(x6326, x6221, x70603);
  nand n6327(x6327, x6220, x6329);
  nand n6328(x6328, x6327, x6326);
  nand n6330(x6330, x6221, x70617);
  nand n6331(x6331, x6220, x6333);
  nand n6332(x6332, x6331, x6330);
  nand n6334(x6334, x6221, x70631);
  nand n6335(x6335, x6220, x6337);
  nand n6336(x6336, x6335, x6334);
  nand n6338(x6338, x6221, x70645);
  nand n6339(x6339, x6220, x6341);
  nand n6340(x6340, x6339, x6338);
  nand n6342(x6342, x6221, x70659);
  nand n6343(x6343, x6220, x6345);
  nand n6344(x6344, x6343, x6342);
  nand n6346(x6346, x6221, x70673);
  nand n6347(x6347, x6220, x6349);
  nand n6348(x6348, x6347, x6346);
  nand n6350(x6350, x2311, x71075);
  nand n6352(x6352, x6351, x70239);
  nand n6353(x6353, x6350, x6355);
  nand n6354(x6354, x6353, x6352);
  nand n6356(x6356, x6351, x70253);
  nand n6357(x6357, x6350, x6359);
  nand n6358(x6358, x6357, x6356);
  nand n6360(x6360, x6351, x70267);
  nand n6361(x6361, x6350, x6363);
  nand n6362(x6362, x6361, x6360);
  nand n6364(x6364, x6351, x70281);
  nand n6365(x6365, x6350, x6367);
  nand n6366(x6366, x6365, x6364);
  nand n6368(x6368, x6351, x70295);
  nand n6369(x6369, x6350, x6371);
  nand n6370(x6370, x6369, x6368);
  nand n6372(x6372, x6351, x70309);
  nand n6373(x6373, x6350, x6375);
  nand n6374(x6374, x6373, x6372);
  nand n6376(x6376, x6351, x70323);
  nand n6377(x6377, x6350, x6379);
  nand n6378(x6378, x6377, x6376);
  nand n6380(x6380, x6351, x70337);
  nand n6381(x6381, x6350, x6383);
  nand n6382(x6382, x6381, x6380);
  nand n6384(x6384, x6351, x70351);
  nand n6385(x6385, x6350, x6387);
  nand n6386(x6386, x6385, x6384);
  nand n6388(x6388, x6351, x70365);
  nand n6389(x6389, x6350, x6391);
  nand n6390(x6390, x6389, x6388);
  nand n6392(x6392, x6351, x70379);
  nand n6393(x6393, x6350, x6395);
  nand n6394(x6394, x6393, x6392);
  nand n6396(x6396, x6351, x70393);
  nand n6397(x6397, x6350, x6399);
  nand n6398(x6398, x6397, x6396);
  nand n6400(x6400, x6351, x70407);
  nand n6401(x6401, x6350, x6403);
  nand n6402(x6402, x6401, x6400);
  nand n6404(x6404, x6351, x70421);
  nand n6405(x6405, x6350, x6407);
  nand n6406(x6406, x6405, x6404);
  nand n6408(x6408, x6351, x70435);
  nand n6409(x6409, x6350, x6411);
  nand n6410(x6410, x6409, x6408);
  nand n6412(x6412, x6351, x70449);
  nand n6413(x6413, x6350, x6415);
  nand n6414(x6414, x6413, x6412);
  nand n6416(x6416, x6351, x70463);
  nand n6417(x6417, x6350, x6419);
  nand n6418(x6418, x6417, x6416);
  nand n6420(x6420, x6351, x70477);
  nand n6421(x6421, x6350, x6423);
  nand n6422(x6422, x6421, x6420);
  nand n6424(x6424, x6351, x70491);
  nand n6425(x6425, x6350, x6427);
  nand n6426(x6426, x6425, x6424);
  nand n6428(x6428, x6351, x70505);
  nand n6429(x6429, x6350, x6431);
  nand n6430(x6430, x6429, x6428);
  nand n6432(x6432, x6351, x70519);
  nand n6433(x6433, x6350, x6435);
  nand n6434(x6434, x6433, x6432);
  nand n6436(x6436, x6351, x70533);
  nand n6437(x6437, x6350, x6439);
  nand n6438(x6438, x6437, x6436);
  nand n6440(x6440, x6351, x70547);
  nand n6441(x6441, x6350, x6443);
  nand n6442(x6442, x6441, x6440);
  nand n6444(x6444, x6351, x70561);
  nand n6445(x6445, x6350, x6447);
  nand n6446(x6446, x6445, x6444);
  nand n6448(x6448, x6351, x70575);
  nand n6449(x6449, x6350, x6451);
  nand n6450(x6450, x6449, x6448);
  nand n6452(x6452, x6351, x70589);
  nand n6453(x6453, x6350, x6455);
  nand n6454(x6454, x6453, x6452);
  nand n6456(x6456, x6351, x70603);
  nand n6457(x6457, x6350, x6459);
  nand n6458(x6458, x6457, x6456);
  nand n6460(x6460, x6351, x70617);
  nand n6461(x6461, x6350, x6463);
  nand n6462(x6462, x6461, x6460);
  nand n6464(x6464, x6351, x70631);
  nand n6465(x6465, x6350, x6467);
  nand n6466(x6466, x6465, x6464);
  nand n6468(x6468, x6351, x70645);
  nand n6469(x6469, x6350, x6471);
  nand n6470(x6470, x6469, x6468);
  nand n6472(x6472, x6351, x70659);
  nand n6473(x6473, x6350, x6475);
  nand n6474(x6474, x6473, x6472);
  nand n6476(x6476, x6351, x70673);
  nand n6477(x6477, x6350, x6479);
  nand n6478(x6478, x6477, x6476);
  nand n6480(x6480, x2258, x3227);
  nand n6482(x6482, x6481, x3097);
  nand n6483(x6483, x6482, x6480);
  nand n6484(x6484, x2258, x2967);
  nand n6485(x6485, x6481, x2837);
  nand n6486(x6486, x6485, x6484);
  nand n6487(x6487, x2258, x2707);
  nand n6488(x6488, x6481, x2577);
  nand n6489(x6489, x6488, x6487);
  nand n6490(x6490, x2258, x2447);
  nand n6491(x6491, x6481, x2317);
  nand n6492(x6492, x6491, x6490);
  nand n6493(x6493, x2261, x6483);
  nand n6495(x6495, x6494, x6486);
  nand n6496(x6496, x6495, x6493);
  nand n6497(x6497, x2261, x6489);
  nand n6498(x6498, x6494, x6492);
  nand n6499(x6499, x6498, x6497);
  nand n6500(x6500, x2264, x6496);
  nand n6502(x6502, x6501, x6499);
  nand n6503(x6503, x6502, x6500);
  nand n6504(x6504, x2258, x3231);
  nand n6505(x6505, x6481, x3101);
  nand n6506(x6506, x6505, x6504);
  nand n6507(x6507, x2258, x2971);
  nand n6508(x6508, x6481, x2841);
  nand n6509(x6509, x6508, x6507);
  nand n6510(x6510, x2258, x2711);
  nand n6511(x6511, x6481, x2581);
  nand n6512(x6512, x6511, x6510);
  nand n6513(x6513, x2258, x2451);
  nand n6514(x6514, x6481, x2321);
  nand n6515(x6515, x6514, x6513);
  nand n6516(x6516, x2261, x6506);
  nand n6517(x6517, x6494, x6509);
  nand n6518(x6518, x6517, x6516);
  nand n6519(x6519, x2261, x6512);
  nand n6520(x6520, x6494, x6515);
  nand n6521(x6521, x6520, x6519);
  nand n6522(x6522, x2264, x6518);
  nand n6523(x6523, x6501, x6521);
  nand n6524(x6524, x6523, x6522);
  nand n6525(x6525, x2258, x3235);
  nand n6526(x6526, x6481, x3105);
  nand n6527(x6527, x6526, x6525);
  nand n6528(x6528, x2258, x2975);
  nand n6529(x6529, x6481, x2845);
  nand n6530(x6530, x6529, x6528);
  nand n6531(x6531, x2258, x2715);
  nand n6532(x6532, x6481, x2585);
  nand n6533(x6533, x6532, x6531);
  nand n6534(x6534, x2258, x2455);
  nand n6535(x6535, x6481, x2325);
  nand n6536(x6536, x6535, x6534);
  nand n6537(x6537, x2261, x6527);
  nand n6538(x6538, x6494, x6530);
  nand n6539(x6539, x6538, x6537);
  nand n6540(x6540, x2261, x6533);
  nand n6541(x6541, x6494, x6536);
  nand n6542(x6542, x6541, x6540);
  nand n6543(x6543, x2264, x6539);
  nand n6544(x6544, x6501, x6542);
  nand n6545(x6545, x6544, x6543);
  nand n6546(x6546, x2258, x3239);
  nand n6547(x6547, x6481, x3109);
  nand n6548(x6548, x6547, x6546);
  nand n6549(x6549, x2258, x2979);
  nand n6550(x6550, x6481, x2849);
  nand n6551(x6551, x6550, x6549);
  nand n6552(x6552, x2258, x2719);
  nand n6553(x6553, x6481, x2589);
  nand n6554(x6554, x6553, x6552);
  nand n6555(x6555, x2258, x2459);
  nand n6556(x6556, x6481, x2329);
  nand n6557(x6557, x6556, x6555);
  nand n6558(x6558, x2261, x6548);
  nand n6559(x6559, x6494, x6551);
  nand n6560(x6560, x6559, x6558);
  nand n6561(x6561, x2261, x6554);
  nand n6562(x6562, x6494, x6557);
  nand n6563(x6563, x6562, x6561);
  nand n6564(x6564, x2264, x6560);
  nand n6565(x6565, x6501, x6563);
  nand n6566(x6566, x6565, x6564);
  nand n6567(x6567, x2258, x3243);
  nand n6568(x6568, x6481, x3113);
  nand n6569(x6569, x6568, x6567);
  nand n6570(x6570, x2258, x2983);
  nand n6571(x6571, x6481, x2853);
  nand n6572(x6572, x6571, x6570);
  nand n6573(x6573, x2258, x2723);
  nand n6574(x6574, x6481, x2593);
  nand n6575(x6575, x6574, x6573);
  nand n6576(x6576, x2258, x2463);
  nand n6577(x6577, x6481, x2333);
  nand n6578(x6578, x6577, x6576);
  nand n6579(x6579, x2261, x6569);
  nand n6580(x6580, x6494, x6572);
  nand n6581(x6581, x6580, x6579);
  nand n6582(x6582, x2261, x6575);
  nand n6583(x6583, x6494, x6578);
  nand n6584(x6584, x6583, x6582);
  nand n6585(x6585, x2264, x6581);
  nand n6586(x6586, x6501, x6584);
  nand n6587(x6587, x6586, x6585);
  nand n6588(x6588, x2258, x3247);
  nand n6589(x6589, x6481, x3117);
  nand n6590(x6590, x6589, x6588);
  nand n6591(x6591, x2258, x2987);
  nand n6592(x6592, x6481, x2857);
  nand n6593(x6593, x6592, x6591);
  nand n6594(x6594, x2258, x2727);
  nand n6595(x6595, x6481, x2597);
  nand n6596(x6596, x6595, x6594);
  nand n6597(x6597, x2258, x2467);
  nand n6598(x6598, x6481, x2337);
  nand n6599(x6599, x6598, x6597);
  nand n6600(x6600, x2261, x6590);
  nand n6601(x6601, x6494, x6593);
  nand n6602(x6602, x6601, x6600);
  nand n6603(x6603, x2261, x6596);
  nand n6604(x6604, x6494, x6599);
  nand n6605(x6605, x6604, x6603);
  nand n6606(x6606, x2264, x6602);
  nand n6607(x6607, x6501, x6605);
  nand n6608(x6608, x6607, x6606);
  nand n6609(x6609, x2258, x3251);
  nand n6610(x6610, x6481, x3121);
  nand n6611(x6611, x6610, x6609);
  nand n6612(x6612, x2258, x2991);
  nand n6613(x6613, x6481, x2861);
  nand n6614(x6614, x6613, x6612);
  nand n6615(x6615, x2258, x2731);
  nand n6616(x6616, x6481, x2601);
  nand n6617(x6617, x6616, x6615);
  nand n6618(x6618, x2258, x2471);
  nand n6619(x6619, x6481, x2341);
  nand n6620(x6620, x6619, x6618);
  nand n6621(x6621, x2261, x6611);
  nand n6622(x6622, x6494, x6614);
  nand n6623(x6623, x6622, x6621);
  nand n6624(x6624, x2261, x6617);
  nand n6625(x6625, x6494, x6620);
  nand n6626(x6626, x6625, x6624);
  nand n6627(x6627, x2264, x6623);
  nand n6628(x6628, x6501, x6626);
  nand n6629(x6629, x6628, x6627);
  nand n6630(x6630, x2258, x3255);
  nand n6631(x6631, x6481, x3125);
  nand n6632(x6632, x6631, x6630);
  nand n6633(x6633, x2258, x2995);
  nand n6634(x6634, x6481, x2865);
  nand n6635(x6635, x6634, x6633);
  nand n6636(x6636, x2258, x2735);
  nand n6637(x6637, x6481, x2605);
  nand n6638(x6638, x6637, x6636);
  nand n6639(x6639, x2258, x2475);
  nand n6640(x6640, x6481, x2345);
  nand n6641(x6641, x6640, x6639);
  nand n6642(x6642, x2261, x6632);
  nand n6643(x6643, x6494, x6635);
  nand n6644(x6644, x6643, x6642);
  nand n6645(x6645, x2261, x6638);
  nand n6646(x6646, x6494, x6641);
  nand n6647(x6647, x6646, x6645);
  nand n6648(x6648, x2264, x6644);
  nand n6649(x6649, x6501, x6647);
  nand n6650(x6650, x6649, x6648);
  nand n6651(x6651, x2258, x3259);
  nand n6652(x6652, x6481, x3129);
  nand n6653(x6653, x6652, x6651);
  nand n6654(x6654, x2258, x2999);
  nand n6655(x6655, x6481, x2869);
  nand n6656(x6656, x6655, x6654);
  nand n6657(x6657, x2258, x2739);
  nand n6658(x6658, x6481, x2609);
  nand n6659(x6659, x6658, x6657);
  nand n6660(x6660, x2258, x2479);
  nand n6661(x6661, x6481, x2349);
  nand n6662(x6662, x6661, x6660);
  nand n6663(x6663, x2261, x6653);
  nand n6664(x6664, x6494, x6656);
  nand n6665(x6665, x6664, x6663);
  nand n6666(x6666, x2261, x6659);
  nand n6667(x6667, x6494, x6662);
  nand n6668(x6668, x6667, x6666);
  nand n6669(x6669, x2264, x6665);
  nand n6670(x6670, x6501, x6668);
  nand n6671(x6671, x6670, x6669);
  nand n6672(x6672, x2258, x3263);
  nand n6673(x6673, x6481, x3133);
  nand n6674(x6674, x6673, x6672);
  nand n6675(x6675, x2258, x3003);
  nand n6676(x6676, x6481, x2873);
  nand n6677(x6677, x6676, x6675);
  nand n6678(x6678, x2258, x2743);
  nand n6679(x6679, x6481, x2613);
  nand n6680(x6680, x6679, x6678);
  nand n6681(x6681, x2258, x2483);
  nand n6682(x6682, x6481, x2353);
  nand n6683(x6683, x6682, x6681);
  nand n6684(x6684, x2261, x6674);
  nand n6685(x6685, x6494, x6677);
  nand n6686(x6686, x6685, x6684);
  nand n6687(x6687, x2261, x6680);
  nand n6688(x6688, x6494, x6683);
  nand n6689(x6689, x6688, x6687);
  nand n6690(x6690, x2264, x6686);
  nand n6691(x6691, x6501, x6689);
  nand n6692(x6692, x6691, x6690);
  nand n6693(x6693, x2258, x3267);
  nand n6694(x6694, x6481, x3137);
  nand n6695(x6695, x6694, x6693);
  nand n6696(x6696, x2258, x3007);
  nand n6697(x6697, x6481, x2877);
  nand n6698(x6698, x6697, x6696);
  nand n6699(x6699, x2258, x2747);
  nand n6700(x6700, x6481, x2617);
  nand n6701(x6701, x6700, x6699);
  nand n6702(x6702, x2258, x2487);
  nand n6703(x6703, x6481, x2357);
  nand n6704(x6704, x6703, x6702);
  nand n6705(x6705, x2261, x6695);
  nand n6706(x6706, x6494, x6698);
  nand n6707(x6707, x6706, x6705);
  nand n6708(x6708, x2261, x6701);
  nand n6709(x6709, x6494, x6704);
  nand n6710(x6710, x6709, x6708);
  nand n6711(x6711, x2264, x6707);
  nand n6712(x6712, x6501, x6710);
  nand n6713(x6713, x6712, x6711);
  nand n6714(x6714, x2258, x3271);
  nand n6715(x6715, x6481, x3141);
  nand n6716(x6716, x6715, x6714);
  nand n6717(x6717, x2258, x3011);
  nand n6718(x6718, x6481, x2881);
  nand n6719(x6719, x6718, x6717);
  nand n6720(x6720, x2258, x2751);
  nand n6721(x6721, x6481, x2621);
  nand n6722(x6722, x6721, x6720);
  nand n6723(x6723, x2258, x2491);
  nand n6724(x6724, x6481, x2361);
  nand n6725(x6725, x6724, x6723);
  nand n6726(x6726, x2261, x6716);
  nand n6727(x6727, x6494, x6719);
  nand n6728(x6728, x6727, x6726);
  nand n6729(x6729, x2261, x6722);
  nand n6730(x6730, x6494, x6725);
  nand n6731(x6731, x6730, x6729);
  nand n6732(x6732, x2264, x6728);
  nand n6733(x6733, x6501, x6731);
  nand n6734(x6734, x6733, x6732);
  nand n6735(x6735, x2258, x3275);
  nand n6736(x6736, x6481, x3145);
  nand n6737(x6737, x6736, x6735);
  nand n6738(x6738, x2258, x3015);
  nand n6739(x6739, x6481, x2885);
  nand n6740(x6740, x6739, x6738);
  nand n6741(x6741, x2258, x2755);
  nand n6742(x6742, x6481, x2625);
  nand n6743(x6743, x6742, x6741);
  nand n6744(x6744, x2258, x2495);
  nand n6745(x6745, x6481, x2365);
  nand n6746(x6746, x6745, x6744);
  nand n6747(x6747, x2261, x6737);
  nand n6748(x6748, x6494, x6740);
  nand n6749(x6749, x6748, x6747);
  nand n6750(x6750, x2261, x6743);
  nand n6751(x6751, x6494, x6746);
  nand n6752(x6752, x6751, x6750);
  nand n6753(x6753, x2264, x6749);
  nand n6754(x6754, x6501, x6752);
  nand n6755(x6755, x6754, x6753);
  nand n6756(x6756, x2258, x3279);
  nand n6757(x6757, x6481, x3149);
  nand n6758(x6758, x6757, x6756);
  nand n6759(x6759, x2258, x3019);
  nand n6760(x6760, x6481, x2889);
  nand n6761(x6761, x6760, x6759);
  nand n6762(x6762, x2258, x2759);
  nand n6763(x6763, x6481, x2629);
  nand n6764(x6764, x6763, x6762);
  nand n6765(x6765, x2258, x2499);
  nand n6766(x6766, x6481, x2369);
  nand n6767(x6767, x6766, x6765);
  nand n6768(x6768, x2261, x6758);
  nand n6769(x6769, x6494, x6761);
  nand n6770(x6770, x6769, x6768);
  nand n6771(x6771, x2261, x6764);
  nand n6772(x6772, x6494, x6767);
  nand n6773(x6773, x6772, x6771);
  nand n6774(x6774, x2264, x6770);
  nand n6775(x6775, x6501, x6773);
  nand n6776(x6776, x6775, x6774);
  nand n6777(x6777, x2258, x3283);
  nand n6778(x6778, x6481, x3153);
  nand n6779(x6779, x6778, x6777);
  nand n6780(x6780, x2258, x3023);
  nand n6781(x6781, x6481, x2893);
  nand n6782(x6782, x6781, x6780);
  nand n6783(x6783, x2258, x2763);
  nand n6784(x6784, x6481, x2633);
  nand n6785(x6785, x6784, x6783);
  nand n6786(x6786, x2258, x2503);
  nand n6787(x6787, x6481, x2373);
  nand n6788(x6788, x6787, x6786);
  nand n6789(x6789, x2261, x6779);
  nand n6790(x6790, x6494, x6782);
  nand n6791(x6791, x6790, x6789);
  nand n6792(x6792, x2261, x6785);
  nand n6793(x6793, x6494, x6788);
  nand n6794(x6794, x6793, x6792);
  nand n6795(x6795, x2264, x6791);
  nand n6796(x6796, x6501, x6794);
  nand n6797(x6797, x6796, x6795);
  nand n6798(x6798, x2258, x3287);
  nand n6799(x6799, x6481, x3157);
  nand n6800(x6800, x6799, x6798);
  nand n6801(x6801, x2258, x3027);
  nand n6802(x6802, x6481, x2897);
  nand n6803(x6803, x6802, x6801);
  nand n6804(x6804, x2258, x2767);
  nand n6805(x6805, x6481, x2637);
  nand n6806(x6806, x6805, x6804);
  nand n6807(x6807, x2258, x2507);
  nand n6808(x6808, x6481, x2377);
  nand n6809(x6809, x6808, x6807);
  nand n6810(x6810, x2261, x6800);
  nand n6811(x6811, x6494, x6803);
  nand n6812(x6812, x6811, x6810);
  nand n6813(x6813, x2261, x6806);
  nand n6814(x6814, x6494, x6809);
  nand n6815(x6815, x6814, x6813);
  nand n6816(x6816, x2264, x6812);
  nand n6817(x6817, x6501, x6815);
  nand n6818(x6818, x6817, x6816);
  nand n6819(x6819, x2258, x3291);
  nand n6820(x6820, x6481, x3161);
  nand n6821(x6821, x6820, x6819);
  nand n6822(x6822, x2258, x3031);
  nand n6823(x6823, x6481, x2901);
  nand n6824(x6824, x6823, x6822);
  nand n6825(x6825, x2258, x2771);
  nand n6826(x6826, x6481, x2641);
  nand n6827(x6827, x6826, x6825);
  nand n6828(x6828, x2258, x2511);
  nand n6829(x6829, x6481, x2381);
  nand n6830(x6830, x6829, x6828);
  nand n6831(x6831, x2261, x6821);
  nand n6832(x6832, x6494, x6824);
  nand n6833(x6833, x6832, x6831);
  nand n6834(x6834, x2261, x6827);
  nand n6835(x6835, x6494, x6830);
  nand n6836(x6836, x6835, x6834);
  nand n6837(x6837, x2264, x6833);
  nand n6838(x6838, x6501, x6836);
  nand n6839(x6839, x6838, x6837);
  nand n6840(x6840, x2258, x3295);
  nand n6841(x6841, x6481, x3165);
  nand n6842(x6842, x6841, x6840);
  nand n6843(x6843, x2258, x3035);
  nand n6844(x6844, x6481, x2905);
  nand n6845(x6845, x6844, x6843);
  nand n6846(x6846, x2258, x2775);
  nand n6847(x6847, x6481, x2645);
  nand n6848(x6848, x6847, x6846);
  nand n6849(x6849, x2258, x2515);
  nand n6850(x6850, x6481, x2385);
  nand n6851(x6851, x6850, x6849);
  nand n6852(x6852, x2261, x6842);
  nand n6853(x6853, x6494, x6845);
  nand n6854(x6854, x6853, x6852);
  nand n6855(x6855, x2261, x6848);
  nand n6856(x6856, x6494, x6851);
  nand n6857(x6857, x6856, x6855);
  nand n6858(x6858, x2264, x6854);
  nand n6859(x6859, x6501, x6857);
  nand n6860(x6860, x6859, x6858);
  nand n6861(x6861, x2258, x3299);
  nand n6862(x6862, x6481, x3169);
  nand n6863(x6863, x6862, x6861);
  nand n6864(x6864, x2258, x3039);
  nand n6865(x6865, x6481, x2909);
  nand n6866(x6866, x6865, x6864);
  nand n6867(x6867, x2258, x2779);
  nand n6868(x6868, x6481, x2649);
  nand n6869(x6869, x6868, x6867);
  nand n6870(x6870, x2258, x2519);
  nand n6871(x6871, x6481, x2389);
  nand n6872(x6872, x6871, x6870);
  nand n6873(x6873, x2261, x6863);
  nand n6874(x6874, x6494, x6866);
  nand n6875(x6875, x6874, x6873);
  nand n6876(x6876, x2261, x6869);
  nand n6877(x6877, x6494, x6872);
  nand n6878(x6878, x6877, x6876);
  nand n6879(x6879, x2264, x6875);
  nand n6880(x6880, x6501, x6878);
  nand n6881(x6881, x6880, x6879);
  nand n6882(x6882, x2258, x3303);
  nand n6883(x6883, x6481, x3173);
  nand n6884(x6884, x6883, x6882);
  nand n6885(x6885, x2258, x3043);
  nand n6886(x6886, x6481, x2913);
  nand n6887(x6887, x6886, x6885);
  nand n6888(x6888, x2258, x2783);
  nand n6889(x6889, x6481, x2653);
  nand n6890(x6890, x6889, x6888);
  nand n6891(x6891, x2258, x2523);
  nand n6892(x6892, x6481, x2393);
  nand n6893(x6893, x6892, x6891);
  nand n6894(x6894, x2261, x6884);
  nand n6895(x6895, x6494, x6887);
  nand n6896(x6896, x6895, x6894);
  nand n6897(x6897, x2261, x6890);
  nand n6898(x6898, x6494, x6893);
  nand n6899(x6899, x6898, x6897);
  nand n6900(x6900, x2264, x6896);
  nand n6901(x6901, x6501, x6899);
  nand n6902(x6902, x6901, x6900);
  nand n6903(x6903, x2258, x3307);
  nand n6904(x6904, x6481, x3177);
  nand n6905(x6905, x6904, x6903);
  nand n6906(x6906, x2258, x3047);
  nand n6907(x6907, x6481, x2917);
  nand n6908(x6908, x6907, x6906);
  nand n6909(x6909, x2258, x2787);
  nand n6910(x6910, x6481, x2657);
  nand n6911(x6911, x6910, x6909);
  nand n6912(x6912, x2258, x2527);
  nand n6913(x6913, x6481, x2397);
  nand n6914(x6914, x6913, x6912);
  nand n6915(x6915, x2261, x6905);
  nand n6916(x6916, x6494, x6908);
  nand n6917(x6917, x6916, x6915);
  nand n6918(x6918, x2261, x6911);
  nand n6919(x6919, x6494, x6914);
  nand n6920(x6920, x6919, x6918);
  nand n6921(x6921, x2264, x6917);
  nand n6922(x6922, x6501, x6920);
  nand n6923(x6923, x6922, x6921);
  nand n6924(x6924, x2258, x3311);
  nand n6925(x6925, x6481, x3181);
  nand n6926(x6926, x6925, x6924);
  nand n6927(x6927, x2258, x3051);
  nand n6928(x6928, x6481, x2921);
  nand n6929(x6929, x6928, x6927);
  nand n6930(x6930, x2258, x2791);
  nand n6931(x6931, x6481, x2661);
  nand n6932(x6932, x6931, x6930);
  nand n6933(x6933, x2258, x2531);
  nand n6934(x6934, x6481, x2401);
  nand n6935(x6935, x6934, x6933);
  nand n6936(x6936, x2261, x6926);
  nand n6937(x6937, x6494, x6929);
  nand n6938(x6938, x6937, x6936);
  nand n6939(x6939, x2261, x6932);
  nand n6940(x6940, x6494, x6935);
  nand n6941(x6941, x6940, x6939);
  nand n6942(x6942, x2264, x6938);
  nand n6943(x6943, x6501, x6941);
  nand n6944(x6944, x6943, x6942);
  nand n6945(x6945, x2258, x3315);
  nand n6946(x6946, x6481, x3185);
  nand n6947(x6947, x6946, x6945);
  nand n6948(x6948, x2258, x3055);
  nand n6949(x6949, x6481, x2925);
  nand n6950(x6950, x6949, x6948);
  nand n6951(x6951, x2258, x2795);
  nand n6952(x6952, x6481, x2665);
  nand n6953(x6953, x6952, x6951);
  nand n6954(x6954, x2258, x2535);
  nand n6955(x6955, x6481, x2405);
  nand n6956(x6956, x6955, x6954);
  nand n6957(x6957, x2261, x6947);
  nand n6958(x6958, x6494, x6950);
  nand n6959(x6959, x6958, x6957);
  nand n6960(x6960, x2261, x6953);
  nand n6961(x6961, x6494, x6956);
  nand n6962(x6962, x6961, x6960);
  nand n6963(x6963, x2264, x6959);
  nand n6964(x6964, x6501, x6962);
  nand n6965(x6965, x6964, x6963);
  nand n6966(x6966, x2258, x3319);
  nand n6967(x6967, x6481, x3189);
  nand n6968(x6968, x6967, x6966);
  nand n6969(x6969, x2258, x3059);
  nand n6970(x6970, x6481, x2929);
  nand n6971(x6971, x6970, x6969);
  nand n6972(x6972, x2258, x2799);
  nand n6973(x6973, x6481, x2669);
  nand n6974(x6974, x6973, x6972);
  nand n6975(x6975, x2258, x2539);
  nand n6976(x6976, x6481, x2409);
  nand n6977(x6977, x6976, x6975);
  nand n6978(x6978, x2261, x6968);
  nand n6979(x6979, x6494, x6971);
  nand n6980(x6980, x6979, x6978);
  nand n6981(x6981, x2261, x6974);
  nand n6982(x6982, x6494, x6977);
  nand n6983(x6983, x6982, x6981);
  nand n6984(x6984, x2264, x6980);
  nand n6985(x6985, x6501, x6983);
  nand n6986(x6986, x6985, x6984);
  nand n6987(x6987, x2258, x3323);
  nand n6988(x6988, x6481, x3193);
  nand n6989(x6989, x6988, x6987);
  nand n6990(x6990, x2258, x3063);
  nand n6991(x6991, x6481, x2933);
  nand n6992(x6992, x6991, x6990);
  nand n6993(x6993, x2258, x2803);
  nand n6994(x6994, x6481, x2673);
  nand n6995(x6995, x6994, x6993);
  nand n6996(x6996, x2258, x2543);
  nand n6997(x6997, x6481, x2413);
  nand n6998(x6998, x6997, x6996);
  nand n6999(x6999, x2261, x6989);
  nand n7000(x7000, x6494, x6992);
  nand n7001(x7001, x7000, x6999);
  nand n7002(x7002, x2261, x6995);
  nand n7003(x7003, x6494, x6998);
  nand n7004(x7004, x7003, x7002);
  nand n7005(x7005, x2264, x7001);
  nand n7006(x7006, x6501, x7004);
  nand n7007(x7007, x7006, x7005);
  nand n7008(x7008, x2258, x3327);
  nand n7009(x7009, x6481, x3197);
  nand n7010(x7010, x7009, x7008);
  nand n7011(x7011, x2258, x3067);
  nand n7012(x7012, x6481, x2937);
  nand n7013(x7013, x7012, x7011);
  nand n7014(x7014, x2258, x2807);
  nand n7015(x7015, x6481, x2677);
  nand n7016(x7016, x7015, x7014);
  nand n7017(x7017, x2258, x2547);
  nand n7018(x7018, x6481, x2417);
  nand n7019(x7019, x7018, x7017);
  nand n7020(x7020, x2261, x7010);
  nand n7021(x7021, x6494, x7013);
  nand n7022(x7022, x7021, x7020);
  nand n7023(x7023, x2261, x7016);
  nand n7024(x7024, x6494, x7019);
  nand n7025(x7025, x7024, x7023);
  nand n7026(x7026, x2264, x7022);
  nand n7027(x7027, x6501, x7025);
  nand n7028(x7028, x7027, x7026);
  nand n7029(x7029, x2258, x3331);
  nand n7030(x7030, x6481, x3201);
  nand n7031(x7031, x7030, x7029);
  nand n7032(x7032, x2258, x3071);
  nand n7033(x7033, x6481, x2941);
  nand n7034(x7034, x7033, x7032);
  nand n7035(x7035, x2258, x2811);
  nand n7036(x7036, x6481, x2681);
  nand n7037(x7037, x7036, x7035);
  nand n7038(x7038, x2258, x2551);
  nand n7039(x7039, x6481, x2421);
  nand n7040(x7040, x7039, x7038);
  nand n7041(x7041, x2261, x7031);
  nand n7042(x7042, x6494, x7034);
  nand n7043(x7043, x7042, x7041);
  nand n7044(x7044, x2261, x7037);
  nand n7045(x7045, x6494, x7040);
  nand n7046(x7046, x7045, x7044);
  nand n7047(x7047, x2264, x7043);
  nand n7048(x7048, x6501, x7046);
  nand n7049(x7049, x7048, x7047);
  nand n7050(x7050, x2258, x3335);
  nand n7051(x7051, x6481, x3205);
  nand n7052(x7052, x7051, x7050);
  nand n7053(x7053, x2258, x3075);
  nand n7054(x7054, x6481, x2945);
  nand n7055(x7055, x7054, x7053);
  nand n7056(x7056, x2258, x2815);
  nand n7057(x7057, x6481, x2685);
  nand n7058(x7058, x7057, x7056);
  nand n7059(x7059, x2258, x2555);
  nand n7060(x7060, x6481, x2425);
  nand n7061(x7061, x7060, x7059);
  nand n7062(x7062, x2261, x7052);
  nand n7063(x7063, x6494, x7055);
  nand n7064(x7064, x7063, x7062);
  nand n7065(x7065, x2261, x7058);
  nand n7066(x7066, x6494, x7061);
  nand n7067(x7067, x7066, x7065);
  nand n7068(x7068, x2264, x7064);
  nand n7069(x7069, x6501, x7067);
  nand n7070(x7070, x7069, x7068);
  nand n7071(x7071, x2258, x3339);
  nand n7072(x7072, x6481, x3209);
  nand n7073(x7073, x7072, x7071);
  nand n7074(x7074, x2258, x3079);
  nand n7075(x7075, x6481, x2949);
  nand n7076(x7076, x7075, x7074);
  nand n7077(x7077, x2258, x2819);
  nand n7078(x7078, x6481, x2689);
  nand n7079(x7079, x7078, x7077);
  nand n7080(x7080, x2258, x2559);
  nand n7081(x7081, x6481, x2429);
  nand n7082(x7082, x7081, x7080);
  nand n7083(x7083, x2261, x7073);
  nand n7084(x7084, x6494, x7076);
  nand n7085(x7085, x7084, x7083);
  nand n7086(x7086, x2261, x7079);
  nand n7087(x7087, x6494, x7082);
  nand n7088(x7088, x7087, x7086);
  nand n7089(x7089, x2264, x7085);
  nand n7090(x7090, x6501, x7088);
  nand n7091(x7091, x7090, x7089);
  nand n7092(x7092, x2258, x3343);
  nand n7093(x7093, x6481, x3213);
  nand n7094(x7094, x7093, x7092);
  nand n7095(x7095, x2258, x3083);
  nand n7096(x7096, x6481, x2953);
  nand n7097(x7097, x7096, x7095);
  nand n7098(x7098, x2258, x2823);
  nand n7099(x7099, x6481, x2693);
  nand n7100(x7100, x7099, x7098);
  nand n7101(x7101, x2258, x2563);
  nand n7102(x7102, x6481, x2433);
  nand n7103(x7103, x7102, x7101);
  nand n7104(x7104, x2261, x7094);
  nand n7105(x7105, x6494, x7097);
  nand n7106(x7106, x7105, x7104);
  nand n7107(x7107, x2261, x7100);
  nand n7108(x7108, x6494, x7103);
  nand n7109(x7109, x7108, x7107);
  nand n7110(x7110, x2264, x7106);
  nand n7111(x7111, x6501, x7109);
  nand n7112(x7112, x7111, x7110);
  nand n7113(x7113, x2258, x3347);
  nand n7114(x7114, x6481, x3217);
  nand n7115(x7115, x7114, x7113);
  nand n7116(x7116, x2258, x3087);
  nand n7117(x7117, x6481, x2957);
  nand n7118(x7118, x7117, x7116);
  nand n7119(x7119, x2258, x2827);
  nand n7120(x7120, x6481, x2697);
  nand n7121(x7121, x7120, x7119);
  nand n7122(x7122, x2258, x2567);
  nand n7123(x7123, x6481, x2437);
  nand n7124(x7124, x7123, x7122);
  nand n7125(x7125, x2261, x7115);
  nand n7126(x7126, x6494, x7118);
  nand n7127(x7127, x7126, x7125);
  nand n7128(x7128, x2261, x7121);
  nand n7129(x7129, x6494, x7124);
  nand n7130(x7130, x7129, x7128);
  nand n7131(x7131, x2264, x7127);
  nand n7132(x7132, x6501, x7130);
  nand n7133(x7133, x7132, x7131);
  nand n7134(x7134, x2258, x3351);
  nand n7135(x7135, x6481, x3221);
  nand n7136(x7136, x7135, x7134);
  nand n7137(x7137, x2258, x3091);
  nand n7138(x7138, x6481, x2961);
  nand n7139(x7139, x7138, x7137);
  nand n7140(x7140, x2258, x2831);
  nand n7141(x7141, x6481, x2701);
  nand n7142(x7142, x7141, x7140);
  nand n7143(x7143, x2258, x2571);
  nand n7144(x7144, x6481, x2441);
  nand n7145(x7145, x7144, x7143);
  nand n7146(x7146, x2261, x7136);
  nand n7147(x7147, x6494, x7139);
  nand n7148(x7148, x7147, x7146);
  nand n7149(x7149, x2261, x7142);
  nand n7150(x7150, x6494, x7145);
  nand n7151(x7151, x7150, x7149);
  nand n7152(x7152, x2264, x7148);
  nand n7153(x7153, x6501, x7151);
  nand n7154(x7154, x7153, x7152);
  nand n7155(x7155, x2269, x3227);
  nand n7157(x7157, x7156, x3097);
  nand n7158(x7158, x7157, x7155);
  nand n7159(x7159, x2269, x2967);
  nand n7160(x7160, x7156, x2837);
  nand n7161(x7161, x7160, x7159);
  nand n7162(x7162, x2269, x2707);
  nand n7163(x7163, x7156, x2577);
  nand n7164(x7164, x7163, x7162);
  nand n7165(x7165, x2269, x2447);
  nand n7166(x7166, x7156, x2317);
  nand n7167(x7167, x7166, x7165);
  nand n7168(x7168, x2272, x7158);
  nand n7170(x7170, x7169, x7161);
  nand n7171(x7171, x7170, x7168);
  nand n7172(x7172, x2272, x7164);
  nand n7173(x7173, x7169, x7167);
  nand n7174(x7174, x7173, x7172);
  nand n7175(x7175, x2275, x7171);
  nand n7177(x7177, x7176, x7174);
  nand n7178(x7178, x7177, x7175);
  nand n7179(x7179, x2269, x3231);
  nand n7180(x7180, x7156, x3101);
  nand n7181(x7181, x7180, x7179);
  nand n7182(x7182, x2269, x2971);
  nand n7183(x7183, x7156, x2841);
  nand n7184(x7184, x7183, x7182);
  nand n7185(x7185, x2269, x2711);
  nand n7186(x7186, x7156, x2581);
  nand n7187(x7187, x7186, x7185);
  nand n7188(x7188, x2269, x2451);
  nand n7189(x7189, x7156, x2321);
  nand n7190(x7190, x7189, x7188);
  nand n7191(x7191, x2272, x7181);
  nand n7192(x7192, x7169, x7184);
  nand n7193(x7193, x7192, x7191);
  nand n7194(x7194, x2272, x7187);
  nand n7195(x7195, x7169, x7190);
  nand n7196(x7196, x7195, x7194);
  nand n7197(x7197, x2275, x7193);
  nand n7198(x7198, x7176, x7196);
  nand n7199(x7199, x7198, x7197);
  nand n7200(x7200, x2269, x3235);
  nand n7201(x7201, x7156, x3105);
  nand n7202(x7202, x7201, x7200);
  nand n7203(x7203, x2269, x2975);
  nand n7204(x7204, x7156, x2845);
  nand n7205(x7205, x7204, x7203);
  nand n7206(x7206, x2269, x2715);
  nand n7207(x7207, x7156, x2585);
  nand n7208(x7208, x7207, x7206);
  nand n7209(x7209, x2269, x2455);
  nand n7210(x7210, x7156, x2325);
  nand n7211(x7211, x7210, x7209);
  nand n7212(x7212, x2272, x7202);
  nand n7213(x7213, x7169, x7205);
  nand n7214(x7214, x7213, x7212);
  nand n7215(x7215, x2272, x7208);
  nand n7216(x7216, x7169, x7211);
  nand n7217(x7217, x7216, x7215);
  nand n7218(x7218, x2275, x7214);
  nand n7219(x7219, x7176, x7217);
  nand n7220(x7220, x7219, x7218);
  nand n7221(x7221, x2269, x3239);
  nand n7222(x7222, x7156, x3109);
  nand n7223(x7223, x7222, x7221);
  nand n7224(x7224, x2269, x2979);
  nand n7225(x7225, x7156, x2849);
  nand n7226(x7226, x7225, x7224);
  nand n7227(x7227, x2269, x2719);
  nand n7228(x7228, x7156, x2589);
  nand n7229(x7229, x7228, x7227);
  nand n7230(x7230, x2269, x2459);
  nand n7231(x7231, x7156, x2329);
  nand n7232(x7232, x7231, x7230);
  nand n7233(x7233, x2272, x7223);
  nand n7234(x7234, x7169, x7226);
  nand n7235(x7235, x7234, x7233);
  nand n7236(x7236, x2272, x7229);
  nand n7237(x7237, x7169, x7232);
  nand n7238(x7238, x7237, x7236);
  nand n7239(x7239, x2275, x7235);
  nand n7240(x7240, x7176, x7238);
  nand n7241(x7241, x7240, x7239);
  nand n7242(x7242, x2269, x3243);
  nand n7243(x7243, x7156, x3113);
  nand n7244(x7244, x7243, x7242);
  nand n7245(x7245, x2269, x2983);
  nand n7246(x7246, x7156, x2853);
  nand n7247(x7247, x7246, x7245);
  nand n7248(x7248, x2269, x2723);
  nand n7249(x7249, x7156, x2593);
  nand n7250(x7250, x7249, x7248);
  nand n7251(x7251, x2269, x2463);
  nand n7252(x7252, x7156, x2333);
  nand n7253(x7253, x7252, x7251);
  nand n7254(x7254, x2272, x7244);
  nand n7255(x7255, x7169, x7247);
  nand n7256(x7256, x7255, x7254);
  nand n7257(x7257, x2272, x7250);
  nand n7258(x7258, x7169, x7253);
  nand n7259(x7259, x7258, x7257);
  nand n7260(x7260, x2275, x7256);
  nand n7261(x7261, x7176, x7259);
  nand n7262(x7262, x7261, x7260);
  nand n7263(x7263, x2269, x3247);
  nand n7264(x7264, x7156, x3117);
  nand n7265(x7265, x7264, x7263);
  nand n7266(x7266, x2269, x2987);
  nand n7267(x7267, x7156, x2857);
  nand n7268(x7268, x7267, x7266);
  nand n7269(x7269, x2269, x2727);
  nand n7270(x7270, x7156, x2597);
  nand n7271(x7271, x7270, x7269);
  nand n7272(x7272, x2269, x2467);
  nand n7273(x7273, x7156, x2337);
  nand n7274(x7274, x7273, x7272);
  nand n7275(x7275, x2272, x7265);
  nand n7276(x7276, x7169, x7268);
  nand n7277(x7277, x7276, x7275);
  nand n7278(x7278, x2272, x7271);
  nand n7279(x7279, x7169, x7274);
  nand n7280(x7280, x7279, x7278);
  nand n7281(x7281, x2275, x7277);
  nand n7282(x7282, x7176, x7280);
  nand n7283(x7283, x7282, x7281);
  nand n7284(x7284, x2269, x3251);
  nand n7285(x7285, x7156, x3121);
  nand n7286(x7286, x7285, x7284);
  nand n7287(x7287, x2269, x2991);
  nand n7288(x7288, x7156, x2861);
  nand n7289(x7289, x7288, x7287);
  nand n7290(x7290, x2269, x2731);
  nand n7291(x7291, x7156, x2601);
  nand n7292(x7292, x7291, x7290);
  nand n7293(x7293, x2269, x2471);
  nand n7294(x7294, x7156, x2341);
  nand n7295(x7295, x7294, x7293);
  nand n7296(x7296, x2272, x7286);
  nand n7297(x7297, x7169, x7289);
  nand n7298(x7298, x7297, x7296);
  nand n7299(x7299, x2272, x7292);
  nand n7300(x7300, x7169, x7295);
  nand n7301(x7301, x7300, x7299);
  nand n7302(x7302, x2275, x7298);
  nand n7303(x7303, x7176, x7301);
  nand n7304(x7304, x7303, x7302);
  nand n7305(x7305, x2269, x3255);
  nand n7306(x7306, x7156, x3125);
  nand n7307(x7307, x7306, x7305);
  nand n7308(x7308, x2269, x2995);
  nand n7309(x7309, x7156, x2865);
  nand n7310(x7310, x7309, x7308);
  nand n7311(x7311, x2269, x2735);
  nand n7312(x7312, x7156, x2605);
  nand n7313(x7313, x7312, x7311);
  nand n7314(x7314, x2269, x2475);
  nand n7315(x7315, x7156, x2345);
  nand n7316(x7316, x7315, x7314);
  nand n7317(x7317, x2272, x7307);
  nand n7318(x7318, x7169, x7310);
  nand n7319(x7319, x7318, x7317);
  nand n7320(x7320, x2272, x7313);
  nand n7321(x7321, x7169, x7316);
  nand n7322(x7322, x7321, x7320);
  nand n7323(x7323, x2275, x7319);
  nand n7324(x7324, x7176, x7322);
  nand n7325(x7325, x7324, x7323);
  nand n7326(x7326, x2269, x3259);
  nand n7327(x7327, x7156, x3129);
  nand n7328(x7328, x7327, x7326);
  nand n7329(x7329, x2269, x2999);
  nand n7330(x7330, x7156, x2869);
  nand n7331(x7331, x7330, x7329);
  nand n7332(x7332, x2269, x2739);
  nand n7333(x7333, x7156, x2609);
  nand n7334(x7334, x7333, x7332);
  nand n7335(x7335, x2269, x2479);
  nand n7336(x7336, x7156, x2349);
  nand n7337(x7337, x7336, x7335);
  nand n7338(x7338, x2272, x7328);
  nand n7339(x7339, x7169, x7331);
  nand n7340(x7340, x7339, x7338);
  nand n7341(x7341, x2272, x7334);
  nand n7342(x7342, x7169, x7337);
  nand n7343(x7343, x7342, x7341);
  nand n7344(x7344, x2275, x7340);
  nand n7345(x7345, x7176, x7343);
  nand n7346(x7346, x7345, x7344);
  nand n7347(x7347, x2269, x3263);
  nand n7348(x7348, x7156, x3133);
  nand n7349(x7349, x7348, x7347);
  nand n7350(x7350, x2269, x3003);
  nand n7351(x7351, x7156, x2873);
  nand n7352(x7352, x7351, x7350);
  nand n7353(x7353, x2269, x2743);
  nand n7354(x7354, x7156, x2613);
  nand n7355(x7355, x7354, x7353);
  nand n7356(x7356, x2269, x2483);
  nand n7357(x7357, x7156, x2353);
  nand n7358(x7358, x7357, x7356);
  nand n7359(x7359, x2272, x7349);
  nand n7360(x7360, x7169, x7352);
  nand n7361(x7361, x7360, x7359);
  nand n7362(x7362, x2272, x7355);
  nand n7363(x7363, x7169, x7358);
  nand n7364(x7364, x7363, x7362);
  nand n7365(x7365, x2275, x7361);
  nand n7366(x7366, x7176, x7364);
  nand n7367(x7367, x7366, x7365);
  nand n7368(x7368, x2269, x3267);
  nand n7369(x7369, x7156, x3137);
  nand n7370(x7370, x7369, x7368);
  nand n7371(x7371, x2269, x3007);
  nand n7372(x7372, x7156, x2877);
  nand n7373(x7373, x7372, x7371);
  nand n7374(x7374, x2269, x2747);
  nand n7375(x7375, x7156, x2617);
  nand n7376(x7376, x7375, x7374);
  nand n7377(x7377, x2269, x2487);
  nand n7378(x7378, x7156, x2357);
  nand n7379(x7379, x7378, x7377);
  nand n7380(x7380, x2272, x7370);
  nand n7381(x7381, x7169, x7373);
  nand n7382(x7382, x7381, x7380);
  nand n7383(x7383, x2272, x7376);
  nand n7384(x7384, x7169, x7379);
  nand n7385(x7385, x7384, x7383);
  nand n7386(x7386, x2275, x7382);
  nand n7387(x7387, x7176, x7385);
  nand n7388(x7388, x7387, x7386);
  nand n7389(x7389, x2269, x3271);
  nand n7390(x7390, x7156, x3141);
  nand n7391(x7391, x7390, x7389);
  nand n7392(x7392, x2269, x3011);
  nand n7393(x7393, x7156, x2881);
  nand n7394(x7394, x7393, x7392);
  nand n7395(x7395, x2269, x2751);
  nand n7396(x7396, x7156, x2621);
  nand n7397(x7397, x7396, x7395);
  nand n7398(x7398, x2269, x2491);
  nand n7399(x7399, x7156, x2361);
  nand n7400(x7400, x7399, x7398);
  nand n7401(x7401, x2272, x7391);
  nand n7402(x7402, x7169, x7394);
  nand n7403(x7403, x7402, x7401);
  nand n7404(x7404, x2272, x7397);
  nand n7405(x7405, x7169, x7400);
  nand n7406(x7406, x7405, x7404);
  nand n7407(x7407, x2275, x7403);
  nand n7408(x7408, x7176, x7406);
  nand n7409(x7409, x7408, x7407);
  nand n7410(x7410, x2269, x3275);
  nand n7411(x7411, x7156, x3145);
  nand n7412(x7412, x7411, x7410);
  nand n7413(x7413, x2269, x3015);
  nand n7414(x7414, x7156, x2885);
  nand n7415(x7415, x7414, x7413);
  nand n7416(x7416, x2269, x2755);
  nand n7417(x7417, x7156, x2625);
  nand n7418(x7418, x7417, x7416);
  nand n7419(x7419, x2269, x2495);
  nand n7420(x7420, x7156, x2365);
  nand n7421(x7421, x7420, x7419);
  nand n7422(x7422, x2272, x7412);
  nand n7423(x7423, x7169, x7415);
  nand n7424(x7424, x7423, x7422);
  nand n7425(x7425, x2272, x7418);
  nand n7426(x7426, x7169, x7421);
  nand n7427(x7427, x7426, x7425);
  nand n7428(x7428, x2275, x7424);
  nand n7429(x7429, x7176, x7427);
  nand n7430(x7430, x7429, x7428);
  nand n7431(x7431, x2269, x3279);
  nand n7432(x7432, x7156, x3149);
  nand n7433(x7433, x7432, x7431);
  nand n7434(x7434, x2269, x3019);
  nand n7435(x7435, x7156, x2889);
  nand n7436(x7436, x7435, x7434);
  nand n7437(x7437, x2269, x2759);
  nand n7438(x7438, x7156, x2629);
  nand n7439(x7439, x7438, x7437);
  nand n7440(x7440, x2269, x2499);
  nand n7441(x7441, x7156, x2369);
  nand n7442(x7442, x7441, x7440);
  nand n7443(x7443, x2272, x7433);
  nand n7444(x7444, x7169, x7436);
  nand n7445(x7445, x7444, x7443);
  nand n7446(x7446, x2272, x7439);
  nand n7447(x7447, x7169, x7442);
  nand n7448(x7448, x7447, x7446);
  nand n7449(x7449, x2275, x7445);
  nand n7450(x7450, x7176, x7448);
  nand n7451(x7451, x7450, x7449);
  nand n7452(x7452, x2269, x3283);
  nand n7453(x7453, x7156, x3153);
  nand n7454(x7454, x7453, x7452);
  nand n7455(x7455, x2269, x3023);
  nand n7456(x7456, x7156, x2893);
  nand n7457(x7457, x7456, x7455);
  nand n7458(x7458, x2269, x2763);
  nand n7459(x7459, x7156, x2633);
  nand n7460(x7460, x7459, x7458);
  nand n7461(x7461, x2269, x2503);
  nand n7462(x7462, x7156, x2373);
  nand n7463(x7463, x7462, x7461);
  nand n7464(x7464, x2272, x7454);
  nand n7465(x7465, x7169, x7457);
  nand n7466(x7466, x7465, x7464);
  nand n7467(x7467, x2272, x7460);
  nand n7468(x7468, x7169, x7463);
  nand n7469(x7469, x7468, x7467);
  nand n7470(x7470, x2275, x7466);
  nand n7471(x7471, x7176, x7469);
  nand n7472(x7472, x7471, x7470);
  nand n7473(x7473, x2269, x3287);
  nand n7474(x7474, x7156, x3157);
  nand n7475(x7475, x7474, x7473);
  nand n7476(x7476, x2269, x3027);
  nand n7477(x7477, x7156, x2897);
  nand n7478(x7478, x7477, x7476);
  nand n7479(x7479, x2269, x2767);
  nand n7480(x7480, x7156, x2637);
  nand n7481(x7481, x7480, x7479);
  nand n7482(x7482, x2269, x2507);
  nand n7483(x7483, x7156, x2377);
  nand n7484(x7484, x7483, x7482);
  nand n7485(x7485, x2272, x7475);
  nand n7486(x7486, x7169, x7478);
  nand n7487(x7487, x7486, x7485);
  nand n7488(x7488, x2272, x7481);
  nand n7489(x7489, x7169, x7484);
  nand n7490(x7490, x7489, x7488);
  nand n7491(x7491, x2275, x7487);
  nand n7492(x7492, x7176, x7490);
  nand n7493(x7493, x7492, x7491);
  nand n7494(x7494, x2269, x3291);
  nand n7495(x7495, x7156, x3161);
  nand n7496(x7496, x7495, x7494);
  nand n7497(x7497, x2269, x3031);
  nand n7498(x7498, x7156, x2901);
  nand n7499(x7499, x7498, x7497);
  nand n7500(x7500, x2269, x2771);
  nand n7501(x7501, x7156, x2641);
  nand n7502(x7502, x7501, x7500);
  nand n7503(x7503, x2269, x2511);
  nand n7504(x7504, x7156, x2381);
  nand n7505(x7505, x7504, x7503);
  nand n7506(x7506, x2272, x7496);
  nand n7507(x7507, x7169, x7499);
  nand n7508(x7508, x7507, x7506);
  nand n7509(x7509, x2272, x7502);
  nand n7510(x7510, x7169, x7505);
  nand n7511(x7511, x7510, x7509);
  nand n7512(x7512, x2275, x7508);
  nand n7513(x7513, x7176, x7511);
  nand n7514(x7514, x7513, x7512);
  nand n7515(x7515, x2269, x3295);
  nand n7516(x7516, x7156, x3165);
  nand n7517(x7517, x7516, x7515);
  nand n7518(x7518, x2269, x3035);
  nand n7519(x7519, x7156, x2905);
  nand n7520(x7520, x7519, x7518);
  nand n7521(x7521, x2269, x2775);
  nand n7522(x7522, x7156, x2645);
  nand n7523(x7523, x7522, x7521);
  nand n7524(x7524, x2269, x2515);
  nand n7525(x7525, x7156, x2385);
  nand n7526(x7526, x7525, x7524);
  nand n7527(x7527, x2272, x7517);
  nand n7528(x7528, x7169, x7520);
  nand n7529(x7529, x7528, x7527);
  nand n7530(x7530, x2272, x7523);
  nand n7531(x7531, x7169, x7526);
  nand n7532(x7532, x7531, x7530);
  nand n7533(x7533, x2275, x7529);
  nand n7534(x7534, x7176, x7532);
  nand n7535(x7535, x7534, x7533);
  nand n7536(x7536, x2269, x3299);
  nand n7537(x7537, x7156, x3169);
  nand n7538(x7538, x7537, x7536);
  nand n7539(x7539, x2269, x3039);
  nand n7540(x7540, x7156, x2909);
  nand n7541(x7541, x7540, x7539);
  nand n7542(x7542, x2269, x2779);
  nand n7543(x7543, x7156, x2649);
  nand n7544(x7544, x7543, x7542);
  nand n7545(x7545, x2269, x2519);
  nand n7546(x7546, x7156, x2389);
  nand n7547(x7547, x7546, x7545);
  nand n7548(x7548, x2272, x7538);
  nand n7549(x7549, x7169, x7541);
  nand n7550(x7550, x7549, x7548);
  nand n7551(x7551, x2272, x7544);
  nand n7552(x7552, x7169, x7547);
  nand n7553(x7553, x7552, x7551);
  nand n7554(x7554, x2275, x7550);
  nand n7555(x7555, x7176, x7553);
  nand n7556(x7556, x7555, x7554);
  nand n7557(x7557, x2269, x3303);
  nand n7558(x7558, x7156, x3173);
  nand n7559(x7559, x7558, x7557);
  nand n7560(x7560, x2269, x3043);
  nand n7561(x7561, x7156, x2913);
  nand n7562(x7562, x7561, x7560);
  nand n7563(x7563, x2269, x2783);
  nand n7564(x7564, x7156, x2653);
  nand n7565(x7565, x7564, x7563);
  nand n7566(x7566, x2269, x2523);
  nand n7567(x7567, x7156, x2393);
  nand n7568(x7568, x7567, x7566);
  nand n7569(x7569, x2272, x7559);
  nand n7570(x7570, x7169, x7562);
  nand n7571(x7571, x7570, x7569);
  nand n7572(x7572, x2272, x7565);
  nand n7573(x7573, x7169, x7568);
  nand n7574(x7574, x7573, x7572);
  nand n7575(x7575, x2275, x7571);
  nand n7576(x7576, x7176, x7574);
  nand n7577(x7577, x7576, x7575);
  nand n7578(x7578, x2269, x3307);
  nand n7579(x7579, x7156, x3177);
  nand n7580(x7580, x7579, x7578);
  nand n7581(x7581, x2269, x3047);
  nand n7582(x7582, x7156, x2917);
  nand n7583(x7583, x7582, x7581);
  nand n7584(x7584, x2269, x2787);
  nand n7585(x7585, x7156, x2657);
  nand n7586(x7586, x7585, x7584);
  nand n7587(x7587, x2269, x2527);
  nand n7588(x7588, x7156, x2397);
  nand n7589(x7589, x7588, x7587);
  nand n7590(x7590, x2272, x7580);
  nand n7591(x7591, x7169, x7583);
  nand n7592(x7592, x7591, x7590);
  nand n7593(x7593, x2272, x7586);
  nand n7594(x7594, x7169, x7589);
  nand n7595(x7595, x7594, x7593);
  nand n7596(x7596, x2275, x7592);
  nand n7597(x7597, x7176, x7595);
  nand n7598(x7598, x7597, x7596);
  nand n7599(x7599, x2269, x3311);
  nand n7600(x7600, x7156, x3181);
  nand n7601(x7601, x7600, x7599);
  nand n7602(x7602, x2269, x3051);
  nand n7603(x7603, x7156, x2921);
  nand n7604(x7604, x7603, x7602);
  nand n7605(x7605, x2269, x2791);
  nand n7606(x7606, x7156, x2661);
  nand n7607(x7607, x7606, x7605);
  nand n7608(x7608, x2269, x2531);
  nand n7609(x7609, x7156, x2401);
  nand n7610(x7610, x7609, x7608);
  nand n7611(x7611, x2272, x7601);
  nand n7612(x7612, x7169, x7604);
  nand n7613(x7613, x7612, x7611);
  nand n7614(x7614, x2272, x7607);
  nand n7615(x7615, x7169, x7610);
  nand n7616(x7616, x7615, x7614);
  nand n7617(x7617, x2275, x7613);
  nand n7618(x7618, x7176, x7616);
  nand n7619(x7619, x7618, x7617);
  nand n7620(x7620, x2269, x3315);
  nand n7621(x7621, x7156, x3185);
  nand n7622(x7622, x7621, x7620);
  nand n7623(x7623, x2269, x3055);
  nand n7624(x7624, x7156, x2925);
  nand n7625(x7625, x7624, x7623);
  nand n7626(x7626, x2269, x2795);
  nand n7627(x7627, x7156, x2665);
  nand n7628(x7628, x7627, x7626);
  nand n7629(x7629, x2269, x2535);
  nand n7630(x7630, x7156, x2405);
  nand n7631(x7631, x7630, x7629);
  nand n7632(x7632, x2272, x7622);
  nand n7633(x7633, x7169, x7625);
  nand n7634(x7634, x7633, x7632);
  nand n7635(x7635, x2272, x7628);
  nand n7636(x7636, x7169, x7631);
  nand n7637(x7637, x7636, x7635);
  nand n7638(x7638, x2275, x7634);
  nand n7639(x7639, x7176, x7637);
  nand n7640(x7640, x7639, x7638);
  nand n7641(x7641, x2269, x3319);
  nand n7642(x7642, x7156, x3189);
  nand n7643(x7643, x7642, x7641);
  nand n7644(x7644, x2269, x3059);
  nand n7645(x7645, x7156, x2929);
  nand n7646(x7646, x7645, x7644);
  nand n7647(x7647, x2269, x2799);
  nand n7648(x7648, x7156, x2669);
  nand n7649(x7649, x7648, x7647);
  nand n7650(x7650, x2269, x2539);
  nand n7651(x7651, x7156, x2409);
  nand n7652(x7652, x7651, x7650);
  nand n7653(x7653, x2272, x7643);
  nand n7654(x7654, x7169, x7646);
  nand n7655(x7655, x7654, x7653);
  nand n7656(x7656, x2272, x7649);
  nand n7657(x7657, x7169, x7652);
  nand n7658(x7658, x7657, x7656);
  nand n7659(x7659, x2275, x7655);
  nand n7660(x7660, x7176, x7658);
  nand n7661(x7661, x7660, x7659);
  nand n7662(x7662, x2269, x3323);
  nand n7663(x7663, x7156, x3193);
  nand n7664(x7664, x7663, x7662);
  nand n7665(x7665, x2269, x3063);
  nand n7666(x7666, x7156, x2933);
  nand n7667(x7667, x7666, x7665);
  nand n7668(x7668, x2269, x2803);
  nand n7669(x7669, x7156, x2673);
  nand n7670(x7670, x7669, x7668);
  nand n7671(x7671, x2269, x2543);
  nand n7672(x7672, x7156, x2413);
  nand n7673(x7673, x7672, x7671);
  nand n7674(x7674, x2272, x7664);
  nand n7675(x7675, x7169, x7667);
  nand n7676(x7676, x7675, x7674);
  nand n7677(x7677, x2272, x7670);
  nand n7678(x7678, x7169, x7673);
  nand n7679(x7679, x7678, x7677);
  nand n7680(x7680, x2275, x7676);
  nand n7681(x7681, x7176, x7679);
  nand n7682(x7682, x7681, x7680);
  nand n7683(x7683, x2269, x3327);
  nand n7684(x7684, x7156, x3197);
  nand n7685(x7685, x7684, x7683);
  nand n7686(x7686, x2269, x3067);
  nand n7687(x7687, x7156, x2937);
  nand n7688(x7688, x7687, x7686);
  nand n7689(x7689, x2269, x2807);
  nand n7690(x7690, x7156, x2677);
  nand n7691(x7691, x7690, x7689);
  nand n7692(x7692, x2269, x2547);
  nand n7693(x7693, x7156, x2417);
  nand n7694(x7694, x7693, x7692);
  nand n7695(x7695, x2272, x7685);
  nand n7696(x7696, x7169, x7688);
  nand n7697(x7697, x7696, x7695);
  nand n7698(x7698, x2272, x7691);
  nand n7699(x7699, x7169, x7694);
  nand n7700(x7700, x7699, x7698);
  nand n7701(x7701, x2275, x7697);
  nand n7702(x7702, x7176, x7700);
  nand n7703(x7703, x7702, x7701);
  nand n7704(x7704, x2269, x3331);
  nand n7705(x7705, x7156, x3201);
  nand n7706(x7706, x7705, x7704);
  nand n7707(x7707, x2269, x3071);
  nand n7708(x7708, x7156, x2941);
  nand n7709(x7709, x7708, x7707);
  nand n7710(x7710, x2269, x2811);
  nand n7711(x7711, x7156, x2681);
  nand n7712(x7712, x7711, x7710);
  nand n7713(x7713, x2269, x2551);
  nand n7714(x7714, x7156, x2421);
  nand n7715(x7715, x7714, x7713);
  nand n7716(x7716, x2272, x7706);
  nand n7717(x7717, x7169, x7709);
  nand n7718(x7718, x7717, x7716);
  nand n7719(x7719, x2272, x7712);
  nand n7720(x7720, x7169, x7715);
  nand n7721(x7721, x7720, x7719);
  nand n7722(x7722, x2275, x7718);
  nand n7723(x7723, x7176, x7721);
  nand n7724(x7724, x7723, x7722);
  nand n7725(x7725, x2269, x3335);
  nand n7726(x7726, x7156, x3205);
  nand n7727(x7727, x7726, x7725);
  nand n7728(x7728, x2269, x3075);
  nand n7729(x7729, x7156, x2945);
  nand n7730(x7730, x7729, x7728);
  nand n7731(x7731, x2269, x2815);
  nand n7732(x7732, x7156, x2685);
  nand n7733(x7733, x7732, x7731);
  nand n7734(x7734, x2269, x2555);
  nand n7735(x7735, x7156, x2425);
  nand n7736(x7736, x7735, x7734);
  nand n7737(x7737, x2272, x7727);
  nand n7738(x7738, x7169, x7730);
  nand n7739(x7739, x7738, x7737);
  nand n7740(x7740, x2272, x7733);
  nand n7741(x7741, x7169, x7736);
  nand n7742(x7742, x7741, x7740);
  nand n7743(x7743, x2275, x7739);
  nand n7744(x7744, x7176, x7742);
  nand n7745(x7745, x7744, x7743);
  nand n7746(x7746, x2269, x3339);
  nand n7747(x7747, x7156, x3209);
  nand n7748(x7748, x7747, x7746);
  nand n7749(x7749, x2269, x3079);
  nand n7750(x7750, x7156, x2949);
  nand n7751(x7751, x7750, x7749);
  nand n7752(x7752, x2269, x2819);
  nand n7753(x7753, x7156, x2689);
  nand n7754(x7754, x7753, x7752);
  nand n7755(x7755, x2269, x2559);
  nand n7756(x7756, x7156, x2429);
  nand n7757(x7757, x7756, x7755);
  nand n7758(x7758, x2272, x7748);
  nand n7759(x7759, x7169, x7751);
  nand n7760(x7760, x7759, x7758);
  nand n7761(x7761, x2272, x7754);
  nand n7762(x7762, x7169, x7757);
  nand n7763(x7763, x7762, x7761);
  nand n7764(x7764, x2275, x7760);
  nand n7765(x7765, x7176, x7763);
  nand n7766(x7766, x7765, x7764);
  nand n7767(x7767, x2269, x3343);
  nand n7768(x7768, x7156, x3213);
  nand n7769(x7769, x7768, x7767);
  nand n7770(x7770, x2269, x3083);
  nand n7771(x7771, x7156, x2953);
  nand n7772(x7772, x7771, x7770);
  nand n7773(x7773, x2269, x2823);
  nand n7774(x7774, x7156, x2693);
  nand n7775(x7775, x7774, x7773);
  nand n7776(x7776, x2269, x2563);
  nand n7777(x7777, x7156, x2433);
  nand n7778(x7778, x7777, x7776);
  nand n7779(x7779, x2272, x7769);
  nand n7780(x7780, x7169, x7772);
  nand n7781(x7781, x7780, x7779);
  nand n7782(x7782, x2272, x7775);
  nand n7783(x7783, x7169, x7778);
  nand n7784(x7784, x7783, x7782);
  nand n7785(x7785, x2275, x7781);
  nand n7786(x7786, x7176, x7784);
  nand n7787(x7787, x7786, x7785);
  nand n7788(x7788, x2269, x3347);
  nand n7789(x7789, x7156, x3217);
  nand n7790(x7790, x7789, x7788);
  nand n7791(x7791, x2269, x3087);
  nand n7792(x7792, x7156, x2957);
  nand n7793(x7793, x7792, x7791);
  nand n7794(x7794, x2269, x2827);
  nand n7795(x7795, x7156, x2697);
  nand n7796(x7796, x7795, x7794);
  nand n7797(x7797, x2269, x2567);
  nand n7798(x7798, x7156, x2437);
  nand n7799(x7799, x7798, x7797);
  nand n7800(x7800, x2272, x7790);
  nand n7801(x7801, x7169, x7793);
  nand n7802(x7802, x7801, x7800);
  nand n7803(x7803, x2272, x7796);
  nand n7804(x7804, x7169, x7799);
  nand n7805(x7805, x7804, x7803);
  nand n7806(x7806, x2275, x7802);
  nand n7807(x7807, x7176, x7805);
  nand n7808(x7808, x7807, x7806);
  nand n7809(x7809, x2269, x3351);
  nand n7810(x7810, x7156, x3221);
  nand n7811(x7811, x7810, x7809);
  nand n7812(x7812, x2269, x3091);
  nand n7813(x7813, x7156, x2961);
  nand n7814(x7814, x7813, x7812);
  nand n7815(x7815, x2269, x2831);
  nand n7816(x7816, x7156, x2701);
  nand n7817(x7817, x7816, x7815);
  nand n7818(x7818, x2269, x2571);
  nand n7819(x7819, x7156, x2441);
  nand n7820(x7820, x7819, x7818);
  nand n7821(x7821, x2272, x7811);
  nand n7822(x7822, x7169, x7814);
  nand n7823(x7823, x7822, x7821);
  nand n7824(x7824, x2272, x7817);
  nand n7825(x7825, x7169, x7820);
  nand n7826(x7826, x7825, x7824);
  nand n7827(x7827, x2275, x7823);
  nand n7828(x7828, x7176, x7826);
  nand n7829(x7829, x7828, x7827);
  nand n7830(x7830, x71202, x3227);
  nand n7831(x7831, x1448, x3097);
  nand n7832(x7832, x7831, x7830);
  nand n7833(x7833, x71202, x2967);
  nand n7834(x7834, x1448, x2837);
  nand n7835(x7835, x7834, x7833);
  nand n7836(x7836, x71202, x2707);
  nand n7837(x7837, x1448, x2577);
  nand n7838(x7838, x7837, x7836);
  nand n7839(x7839, x71202, x2447);
  nand n7840(x7840, x1448, x2317);
  nand n7841(x7841, x7840, x7839);
  nand n7842(x7842, x71205, x7832);
  nand n7843(x7843, x1461, x7835);
  nand n7844(x7844, x7843, x7842);
  nand n7845(x7845, x71205, x7838);
  nand n7846(x7846, x1461, x7841);
  nand n7847(x7847, x7846, x7845);
  nand n7848(x7848, x71210, x7844);
  nand n7849(x7849, x1468, x7847);
  nand n7850(x7850, x7849, x7848);
  nand n7851(x7851, x71202, x3231);
  nand n7852(x7852, x1448, x3101);
  nand n7853(x7853, x7852, x7851);
  nand n7854(x7854, x71202, x2971);
  nand n7855(x7855, x1448, x2841);
  nand n7856(x7856, x7855, x7854);
  nand n7857(x7857, x71202, x2711);
  nand n7858(x7858, x1448, x2581);
  nand n7859(x7859, x7858, x7857);
  nand n7860(x7860, x71202, x2451);
  nand n7861(x7861, x1448, x2321);
  nand n7862(x7862, x7861, x7860);
  nand n7863(x7863, x71205, x7853);
  nand n7864(x7864, x1461, x7856);
  nand n7865(x7865, x7864, x7863);
  nand n7866(x7866, x71205, x7859);
  nand n7867(x7867, x1461, x7862);
  nand n7868(x7868, x7867, x7866);
  nand n7869(x7869, x71210, x7865);
  nand n7870(x7870, x1468, x7868);
  nand n7871(x7871, x7870, x7869);
  nand n7872(x7872, x71202, x3235);
  nand n7873(x7873, x1448, x3105);
  nand n7874(x7874, x7873, x7872);
  nand n7875(x7875, x71202, x2975);
  nand n7876(x7876, x1448, x2845);
  nand n7877(x7877, x7876, x7875);
  nand n7878(x7878, x71202, x2715);
  nand n7879(x7879, x1448, x2585);
  nand n7880(x7880, x7879, x7878);
  nand n7881(x7881, x71202, x2455);
  nand n7882(x7882, x1448, x2325);
  nand n7883(x7883, x7882, x7881);
  nand n7884(x7884, x71205, x7874);
  nand n7885(x7885, x1461, x7877);
  nand n7886(x7886, x7885, x7884);
  nand n7887(x7887, x71205, x7880);
  nand n7888(x7888, x1461, x7883);
  nand n7889(x7889, x7888, x7887);
  nand n7890(x7890, x71210, x7886);
  nand n7891(x7891, x1468, x7889);
  nand n7892(x7892, x7891, x7890);
  nand n7893(x7893, x71202, x3239);
  nand n7894(x7894, x1448, x3109);
  nand n7895(x7895, x7894, x7893);
  nand n7896(x7896, x71202, x2979);
  nand n7897(x7897, x1448, x2849);
  nand n7898(x7898, x7897, x7896);
  nand n7899(x7899, x71202, x2719);
  nand n7900(x7900, x1448, x2589);
  nand n7901(x7901, x7900, x7899);
  nand n7902(x7902, x71202, x2459);
  nand n7903(x7903, x1448, x2329);
  nand n7904(x7904, x7903, x7902);
  nand n7905(x7905, x71205, x7895);
  nand n7906(x7906, x1461, x7898);
  nand n7907(x7907, x7906, x7905);
  nand n7908(x7908, x71205, x7901);
  nand n7909(x7909, x1461, x7904);
  nand n7910(x7910, x7909, x7908);
  nand n7911(x7911, x71210, x7907);
  nand n7912(x7912, x1468, x7910);
  nand n7913(x7913, x7912, x7911);
  nand n7914(x7914, x71202, x3243);
  nand n7915(x7915, x1448, x3113);
  nand n7916(x7916, x7915, x7914);
  nand n7917(x7917, x71202, x2983);
  nand n7918(x7918, x1448, x2853);
  nand n7919(x7919, x7918, x7917);
  nand n7920(x7920, x71202, x2723);
  nand n7921(x7921, x1448, x2593);
  nand n7922(x7922, x7921, x7920);
  nand n7923(x7923, x71202, x2463);
  nand n7924(x7924, x1448, x2333);
  nand n7925(x7925, x7924, x7923);
  nand n7926(x7926, x71205, x7916);
  nand n7927(x7927, x1461, x7919);
  nand n7928(x7928, x7927, x7926);
  nand n7929(x7929, x71205, x7922);
  nand n7930(x7930, x1461, x7925);
  nand n7931(x7931, x7930, x7929);
  nand n7932(x7932, x71210, x7928);
  nand n7933(x7933, x1468, x7931);
  nand n7934(x7934, x7933, x7932);
  nand n7935(x7935, x71202, x3247);
  nand n7936(x7936, x1448, x3117);
  nand n7937(x7937, x7936, x7935);
  nand n7938(x7938, x71202, x2987);
  nand n7939(x7939, x1448, x2857);
  nand n7940(x7940, x7939, x7938);
  nand n7941(x7941, x71202, x2727);
  nand n7942(x7942, x1448, x2597);
  nand n7943(x7943, x7942, x7941);
  nand n7944(x7944, x71202, x2467);
  nand n7945(x7945, x1448, x2337);
  nand n7946(x7946, x7945, x7944);
  nand n7947(x7947, x71205, x7937);
  nand n7948(x7948, x1461, x7940);
  nand n7949(x7949, x7948, x7947);
  nand n7950(x7950, x71205, x7943);
  nand n7951(x7951, x1461, x7946);
  nand n7952(x7952, x7951, x7950);
  nand n7953(x7953, x71210, x7949);
  nand n7954(x7954, x1468, x7952);
  nand n7955(x7955, x7954, x7953);
  nand n7956(x7956, x71202, x3251);
  nand n7957(x7957, x1448, x3121);
  nand n7958(x7958, x7957, x7956);
  nand n7959(x7959, x71202, x2991);
  nand n7960(x7960, x1448, x2861);
  nand n7961(x7961, x7960, x7959);
  nand n7962(x7962, x71202, x2731);
  nand n7963(x7963, x1448, x2601);
  nand n7964(x7964, x7963, x7962);
  nand n7965(x7965, x71202, x2471);
  nand n7966(x7966, x1448, x2341);
  nand n7967(x7967, x7966, x7965);
  nand n7968(x7968, x71205, x7958);
  nand n7969(x7969, x1461, x7961);
  nand n7970(x7970, x7969, x7968);
  nand n7971(x7971, x71205, x7964);
  nand n7972(x7972, x1461, x7967);
  nand n7973(x7973, x7972, x7971);
  nand n7974(x7974, x71210, x7970);
  nand n7975(x7975, x1468, x7973);
  nand n7976(x7976, x7975, x7974);
  nand n7977(x7977, x71202, x3255);
  nand n7978(x7978, x1448, x3125);
  nand n7979(x7979, x7978, x7977);
  nand n7980(x7980, x71202, x2995);
  nand n7981(x7981, x1448, x2865);
  nand n7982(x7982, x7981, x7980);
  nand n7983(x7983, x71202, x2735);
  nand n7984(x7984, x1448, x2605);
  nand n7985(x7985, x7984, x7983);
  nand n7986(x7986, x71202, x2475);
  nand n7987(x7987, x1448, x2345);
  nand n7988(x7988, x7987, x7986);
  nand n7989(x7989, x71205, x7979);
  nand n7990(x7990, x1461, x7982);
  nand n7991(x7991, x7990, x7989);
  nand n7992(x7992, x71205, x7985);
  nand n7993(x7993, x1461, x7988);
  nand n7994(x7994, x7993, x7992);
  nand n7995(x7995, x71210, x7991);
  nand n7996(x7996, x1468, x7994);
  nand n7997(x7997, x7996, x7995);
  nand n7998(x7998, x71202, x3259);
  nand n7999(x7999, x1448, x3129);
  nand n8000(x8000, x7999, x7998);
  nand n8001(x8001, x71202, x2999);
  nand n8002(x8002, x1448, x2869);
  nand n8003(x8003, x8002, x8001);
  nand n8004(x8004, x71202, x2739);
  nand n8005(x8005, x1448, x2609);
  nand n8006(x8006, x8005, x8004);
  nand n8007(x8007, x71202, x2479);
  nand n8008(x8008, x1448, x2349);
  nand n8009(x8009, x8008, x8007);
  nand n8010(x8010, x71205, x8000);
  nand n8011(x8011, x1461, x8003);
  nand n8012(x8012, x8011, x8010);
  nand n8013(x8013, x71205, x8006);
  nand n8014(x8014, x1461, x8009);
  nand n8015(x8015, x8014, x8013);
  nand n8016(x8016, x71210, x8012);
  nand n8017(x8017, x1468, x8015);
  nand n8018(x8018, x8017, x8016);
  nand n8019(x8019, x71202, x3263);
  nand n8020(x8020, x1448, x3133);
  nand n8021(x8021, x8020, x8019);
  nand n8022(x8022, x71202, x3003);
  nand n8023(x8023, x1448, x2873);
  nand n8024(x8024, x8023, x8022);
  nand n8025(x8025, x71202, x2743);
  nand n8026(x8026, x1448, x2613);
  nand n8027(x8027, x8026, x8025);
  nand n8028(x8028, x71202, x2483);
  nand n8029(x8029, x1448, x2353);
  nand n8030(x8030, x8029, x8028);
  nand n8031(x8031, x71205, x8021);
  nand n8032(x8032, x1461, x8024);
  nand n8033(x8033, x8032, x8031);
  nand n8034(x8034, x71205, x8027);
  nand n8035(x8035, x1461, x8030);
  nand n8036(x8036, x8035, x8034);
  nand n8037(x8037, x71210, x8033);
  nand n8038(x8038, x1468, x8036);
  nand n8039(x8039, x8038, x8037);
  nand n8040(x8040, x71202, x3267);
  nand n8041(x8041, x1448, x3137);
  nand n8042(x8042, x8041, x8040);
  nand n8043(x8043, x71202, x3007);
  nand n8044(x8044, x1448, x2877);
  nand n8045(x8045, x8044, x8043);
  nand n8046(x8046, x71202, x2747);
  nand n8047(x8047, x1448, x2617);
  nand n8048(x8048, x8047, x8046);
  nand n8049(x8049, x71202, x2487);
  nand n8050(x8050, x1448, x2357);
  nand n8051(x8051, x8050, x8049);
  nand n8052(x8052, x71205, x8042);
  nand n8053(x8053, x1461, x8045);
  nand n8054(x8054, x8053, x8052);
  nand n8055(x8055, x71205, x8048);
  nand n8056(x8056, x1461, x8051);
  nand n8057(x8057, x8056, x8055);
  nand n8058(x8058, x71210, x8054);
  nand n8059(x8059, x1468, x8057);
  nand n8060(x8060, x8059, x8058);
  nand n8061(x8061, x71202, x3271);
  nand n8062(x8062, x1448, x3141);
  nand n8063(x8063, x8062, x8061);
  nand n8064(x8064, x71202, x3011);
  nand n8065(x8065, x1448, x2881);
  nand n8066(x8066, x8065, x8064);
  nand n8067(x8067, x71202, x2751);
  nand n8068(x8068, x1448, x2621);
  nand n8069(x8069, x8068, x8067);
  nand n8070(x8070, x71202, x2491);
  nand n8071(x8071, x1448, x2361);
  nand n8072(x8072, x8071, x8070);
  nand n8073(x8073, x71205, x8063);
  nand n8074(x8074, x1461, x8066);
  nand n8075(x8075, x8074, x8073);
  nand n8076(x8076, x71205, x8069);
  nand n8077(x8077, x1461, x8072);
  nand n8078(x8078, x8077, x8076);
  nand n8079(x8079, x71210, x8075);
  nand n8080(x8080, x1468, x8078);
  nand n8081(x8081, x8080, x8079);
  nand n8082(x8082, x71202, x3275);
  nand n8083(x8083, x1448, x3145);
  nand n8084(x8084, x8083, x8082);
  nand n8085(x8085, x71202, x3015);
  nand n8086(x8086, x1448, x2885);
  nand n8087(x8087, x8086, x8085);
  nand n8088(x8088, x71202, x2755);
  nand n8089(x8089, x1448, x2625);
  nand n8090(x8090, x8089, x8088);
  nand n8091(x8091, x71202, x2495);
  nand n8092(x8092, x1448, x2365);
  nand n8093(x8093, x8092, x8091);
  nand n8094(x8094, x71205, x8084);
  nand n8095(x8095, x1461, x8087);
  nand n8096(x8096, x8095, x8094);
  nand n8097(x8097, x71205, x8090);
  nand n8098(x8098, x1461, x8093);
  nand n8099(x8099, x8098, x8097);
  nand n8100(x8100, x71210, x8096);
  nand n8101(x8101, x1468, x8099);
  nand n8102(x8102, x8101, x8100);
  nand n8103(x8103, x71202, x3279);
  nand n8104(x8104, x1448, x3149);
  nand n8105(x8105, x8104, x8103);
  nand n8106(x8106, x71202, x3019);
  nand n8107(x8107, x1448, x2889);
  nand n8108(x8108, x8107, x8106);
  nand n8109(x8109, x71202, x2759);
  nand n8110(x8110, x1448, x2629);
  nand n8111(x8111, x8110, x8109);
  nand n8112(x8112, x71202, x2499);
  nand n8113(x8113, x1448, x2369);
  nand n8114(x8114, x8113, x8112);
  nand n8115(x8115, x71205, x8105);
  nand n8116(x8116, x1461, x8108);
  nand n8117(x8117, x8116, x8115);
  nand n8118(x8118, x71205, x8111);
  nand n8119(x8119, x1461, x8114);
  nand n8120(x8120, x8119, x8118);
  nand n8121(x8121, x71210, x8117);
  nand n8122(x8122, x1468, x8120);
  nand n8123(x8123, x8122, x8121);
  nand n8124(x8124, x71202, x3283);
  nand n8125(x8125, x1448, x3153);
  nand n8126(x8126, x8125, x8124);
  nand n8127(x8127, x71202, x3023);
  nand n8128(x8128, x1448, x2893);
  nand n8129(x8129, x8128, x8127);
  nand n8130(x8130, x71202, x2763);
  nand n8131(x8131, x1448, x2633);
  nand n8132(x8132, x8131, x8130);
  nand n8133(x8133, x71202, x2503);
  nand n8134(x8134, x1448, x2373);
  nand n8135(x8135, x8134, x8133);
  nand n8136(x8136, x71205, x8126);
  nand n8137(x8137, x1461, x8129);
  nand n8138(x8138, x8137, x8136);
  nand n8139(x8139, x71205, x8132);
  nand n8140(x8140, x1461, x8135);
  nand n8141(x8141, x8140, x8139);
  nand n8142(x8142, x71210, x8138);
  nand n8143(x8143, x1468, x8141);
  nand n8144(x8144, x8143, x8142);
  nand n8145(x8145, x71202, x3287);
  nand n8146(x8146, x1448, x3157);
  nand n8147(x8147, x8146, x8145);
  nand n8148(x8148, x71202, x3027);
  nand n8149(x8149, x1448, x2897);
  nand n8150(x8150, x8149, x8148);
  nand n8151(x8151, x71202, x2767);
  nand n8152(x8152, x1448, x2637);
  nand n8153(x8153, x8152, x8151);
  nand n8154(x8154, x71202, x2507);
  nand n8155(x8155, x1448, x2377);
  nand n8156(x8156, x8155, x8154);
  nand n8157(x8157, x71205, x8147);
  nand n8158(x8158, x1461, x8150);
  nand n8159(x8159, x8158, x8157);
  nand n8160(x8160, x71205, x8153);
  nand n8161(x8161, x1461, x8156);
  nand n8162(x8162, x8161, x8160);
  nand n8163(x8163, x71210, x8159);
  nand n8164(x8164, x1468, x8162);
  nand n8165(x8165, x8164, x8163);
  nand n8166(x8166, x71202, x3291);
  nand n8167(x8167, x1448, x3161);
  nand n8168(x8168, x8167, x8166);
  nand n8169(x8169, x71202, x3031);
  nand n8170(x8170, x1448, x2901);
  nand n8171(x8171, x8170, x8169);
  nand n8172(x8172, x71202, x2771);
  nand n8173(x8173, x1448, x2641);
  nand n8174(x8174, x8173, x8172);
  nand n8175(x8175, x71202, x2511);
  nand n8176(x8176, x1448, x2381);
  nand n8177(x8177, x8176, x8175);
  nand n8178(x8178, x71205, x8168);
  nand n8179(x8179, x1461, x8171);
  nand n8180(x8180, x8179, x8178);
  nand n8181(x8181, x71205, x8174);
  nand n8182(x8182, x1461, x8177);
  nand n8183(x8183, x8182, x8181);
  nand n8184(x8184, x71210, x8180);
  nand n8185(x8185, x1468, x8183);
  nand n8186(x8186, x8185, x8184);
  nand n8187(x8187, x71202, x3295);
  nand n8188(x8188, x1448, x3165);
  nand n8189(x8189, x8188, x8187);
  nand n8190(x8190, x71202, x3035);
  nand n8191(x8191, x1448, x2905);
  nand n8192(x8192, x8191, x8190);
  nand n8193(x8193, x71202, x2775);
  nand n8194(x8194, x1448, x2645);
  nand n8195(x8195, x8194, x8193);
  nand n8196(x8196, x71202, x2515);
  nand n8197(x8197, x1448, x2385);
  nand n8198(x8198, x8197, x8196);
  nand n8199(x8199, x71205, x8189);
  nand n8200(x8200, x1461, x8192);
  nand n8201(x8201, x8200, x8199);
  nand n8202(x8202, x71205, x8195);
  nand n8203(x8203, x1461, x8198);
  nand n8204(x8204, x8203, x8202);
  nand n8205(x8205, x71210, x8201);
  nand n8206(x8206, x1468, x8204);
  nand n8207(x8207, x8206, x8205);
  nand n8208(x8208, x71202, x3299);
  nand n8209(x8209, x1448, x3169);
  nand n8210(x8210, x8209, x8208);
  nand n8211(x8211, x71202, x3039);
  nand n8212(x8212, x1448, x2909);
  nand n8213(x8213, x8212, x8211);
  nand n8214(x8214, x71202, x2779);
  nand n8215(x8215, x1448, x2649);
  nand n8216(x8216, x8215, x8214);
  nand n8217(x8217, x71202, x2519);
  nand n8218(x8218, x1448, x2389);
  nand n8219(x8219, x8218, x8217);
  nand n8220(x8220, x71205, x8210);
  nand n8221(x8221, x1461, x8213);
  nand n8222(x8222, x8221, x8220);
  nand n8223(x8223, x71205, x8216);
  nand n8224(x8224, x1461, x8219);
  nand n8225(x8225, x8224, x8223);
  nand n8226(x8226, x71210, x8222);
  nand n8227(x8227, x1468, x8225);
  nand n8228(x8228, x8227, x8226);
  nand n8229(x8229, x71202, x3303);
  nand n8230(x8230, x1448, x3173);
  nand n8231(x8231, x8230, x8229);
  nand n8232(x8232, x71202, x3043);
  nand n8233(x8233, x1448, x2913);
  nand n8234(x8234, x8233, x8232);
  nand n8235(x8235, x71202, x2783);
  nand n8236(x8236, x1448, x2653);
  nand n8237(x8237, x8236, x8235);
  nand n8238(x8238, x71202, x2523);
  nand n8239(x8239, x1448, x2393);
  nand n8240(x8240, x8239, x8238);
  nand n8241(x8241, x71205, x8231);
  nand n8242(x8242, x1461, x8234);
  nand n8243(x8243, x8242, x8241);
  nand n8244(x8244, x71205, x8237);
  nand n8245(x8245, x1461, x8240);
  nand n8246(x8246, x8245, x8244);
  nand n8247(x8247, x71210, x8243);
  nand n8248(x8248, x1468, x8246);
  nand n8249(x8249, x8248, x8247);
  nand n8250(x8250, x71202, x3307);
  nand n8251(x8251, x1448, x3177);
  nand n8252(x8252, x8251, x8250);
  nand n8253(x8253, x71202, x3047);
  nand n8254(x8254, x1448, x2917);
  nand n8255(x8255, x8254, x8253);
  nand n8256(x8256, x71202, x2787);
  nand n8257(x8257, x1448, x2657);
  nand n8258(x8258, x8257, x8256);
  nand n8259(x8259, x71202, x2527);
  nand n8260(x8260, x1448, x2397);
  nand n8261(x8261, x8260, x8259);
  nand n8262(x8262, x71205, x8252);
  nand n8263(x8263, x1461, x8255);
  nand n8264(x8264, x8263, x8262);
  nand n8265(x8265, x71205, x8258);
  nand n8266(x8266, x1461, x8261);
  nand n8267(x8267, x8266, x8265);
  nand n8268(x8268, x71210, x8264);
  nand n8269(x8269, x1468, x8267);
  nand n8270(x8270, x8269, x8268);
  nand n8271(x8271, x71202, x3311);
  nand n8272(x8272, x1448, x3181);
  nand n8273(x8273, x8272, x8271);
  nand n8274(x8274, x71202, x3051);
  nand n8275(x8275, x1448, x2921);
  nand n8276(x8276, x8275, x8274);
  nand n8277(x8277, x71202, x2791);
  nand n8278(x8278, x1448, x2661);
  nand n8279(x8279, x8278, x8277);
  nand n8280(x8280, x71202, x2531);
  nand n8281(x8281, x1448, x2401);
  nand n8282(x8282, x8281, x8280);
  nand n8283(x8283, x71205, x8273);
  nand n8284(x8284, x1461, x8276);
  nand n8285(x8285, x8284, x8283);
  nand n8286(x8286, x71205, x8279);
  nand n8287(x8287, x1461, x8282);
  nand n8288(x8288, x8287, x8286);
  nand n8289(x8289, x71210, x8285);
  nand n8290(x8290, x1468, x8288);
  nand n8291(x8291, x8290, x8289);
  nand n8292(x8292, x71202, x3315);
  nand n8293(x8293, x1448, x3185);
  nand n8294(x8294, x8293, x8292);
  nand n8295(x8295, x71202, x3055);
  nand n8296(x8296, x1448, x2925);
  nand n8297(x8297, x8296, x8295);
  nand n8298(x8298, x71202, x2795);
  nand n8299(x8299, x1448, x2665);
  nand n8300(x8300, x8299, x8298);
  nand n8301(x8301, x71202, x2535);
  nand n8302(x8302, x1448, x2405);
  nand n8303(x8303, x8302, x8301);
  nand n8304(x8304, x71205, x8294);
  nand n8305(x8305, x1461, x8297);
  nand n8306(x8306, x8305, x8304);
  nand n8307(x8307, x71205, x8300);
  nand n8308(x8308, x1461, x8303);
  nand n8309(x8309, x8308, x8307);
  nand n8310(x8310, x71210, x8306);
  nand n8311(x8311, x1468, x8309);
  nand n8312(x8312, x8311, x8310);
  nand n8313(x8313, x71202, x3319);
  nand n8314(x8314, x1448, x3189);
  nand n8315(x8315, x8314, x8313);
  nand n8316(x8316, x71202, x3059);
  nand n8317(x8317, x1448, x2929);
  nand n8318(x8318, x8317, x8316);
  nand n8319(x8319, x71202, x2799);
  nand n8320(x8320, x1448, x2669);
  nand n8321(x8321, x8320, x8319);
  nand n8322(x8322, x71202, x2539);
  nand n8323(x8323, x1448, x2409);
  nand n8324(x8324, x8323, x8322);
  nand n8325(x8325, x71205, x8315);
  nand n8326(x8326, x1461, x8318);
  nand n8327(x8327, x8326, x8325);
  nand n8328(x8328, x71205, x8321);
  nand n8329(x8329, x1461, x8324);
  nand n8330(x8330, x8329, x8328);
  nand n8331(x8331, x71210, x8327);
  nand n8332(x8332, x1468, x8330);
  nand n8333(x8333, x8332, x8331);
  nand n8334(x8334, x71202, x3323);
  nand n8335(x8335, x1448, x3193);
  nand n8336(x8336, x8335, x8334);
  nand n8337(x8337, x71202, x3063);
  nand n8338(x8338, x1448, x2933);
  nand n8339(x8339, x8338, x8337);
  nand n8340(x8340, x71202, x2803);
  nand n8341(x8341, x1448, x2673);
  nand n8342(x8342, x8341, x8340);
  nand n8343(x8343, x71202, x2543);
  nand n8344(x8344, x1448, x2413);
  nand n8345(x8345, x8344, x8343);
  nand n8346(x8346, x71205, x8336);
  nand n8347(x8347, x1461, x8339);
  nand n8348(x8348, x8347, x8346);
  nand n8349(x8349, x71205, x8342);
  nand n8350(x8350, x1461, x8345);
  nand n8351(x8351, x8350, x8349);
  nand n8352(x8352, x71210, x8348);
  nand n8353(x8353, x1468, x8351);
  nand n8354(x8354, x8353, x8352);
  nand n8355(x8355, x71202, x3327);
  nand n8356(x8356, x1448, x3197);
  nand n8357(x8357, x8356, x8355);
  nand n8358(x8358, x71202, x3067);
  nand n8359(x8359, x1448, x2937);
  nand n8360(x8360, x8359, x8358);
  nand n8361(x8361, x71202, x2807);
  nand n8362(x8362, x1448, x2677);
  nand n8363(x8363, x8362, x8361);
  nand n8364(x8364, x71202, x2547);
  nand n8365(x8365, x1448, x2417);
  nand n8366(x8366, x8365, x8364);
  nand n8367(x8367, x71205, x8357);
  nand n8368(x8368, x1461, x8360);
  nand n8369(x8369, x8368, x8367);
  nand n8370(x8370, x71205, x8363);
  nand n8371(x8371, x1461, x8366);
  nand n8372(x8372, x8371, x8370);
  nand n8373(x8373, x71210, x8369);
  nand n8374(x8374, x1468, x8372);
  nand n8375(x8375, x8374, x8373);
  nand n8376(x8376, x71202, x3331);
  nand n8377(x8377, x1448, x3201);
  nand n8378(x8378, x8377, x8376);
  nand n8379(x8379, x71202, x3071);
  nand n8380(x8380, x1448, x2941);
  nand n8381(x8381, x8380, x8379);
  nand n8382(x8382, x71202, x2811);
  nand n8383(x8383, x1448, x2681);
  nand n8384(x8384, x8383, x8382);
  nand n8385(x8385, x71202, x2551);
  nand n8386(x8386, x1448, x2421);
  nand n8387(x8387, x8386, x8385);
  nand n8388(x8388, x71205, x8378);
  nand n8389(x8389, x1461, x8381);
  nand n8390(x8390, x8389, x8388);
  nand n8391(x8391, x71205, x8384);
  nand n8392(x8392, x1461, x8387);
  nand n8393(x8393, x8392, x8391);
  nand n8394(x8394, x71210, x8390);
  nand n8395(x8395, x1468, x8393);
  nand n8396(x8396, x8395, x8394);
  nand n8397(x8397, x71202, x3335);
  nand n8398(x8398, x1448, x3205);
  nand n8399(x8399, x8398, x8397);
  nand n8400(x8400, x71202, x3075);
  nand n8401(x8401, x1448, x2945);
  nand n8402(x8402, x8401, x8400);
  nand n8403(x8403, x71202, x2815);
  nand n8404(x8404, x1448, x2685);
  nand n8405(x8405, x8404, x8403);
  nand n8406(x8406, x71202, x2555);
  nand n8407(x8407, x1448, x2425);
  nand n8408(x8408, x8407, x8406);
  nand n8409(x8409, x71205, x8399);
  nand n8410(x8410, x1461, x8402);
  nand n8411(x8411, x8410, x8409);
  nand n8412(x8412, x71205, x8405);
  nand n8413(x8413, x1461, x8408);
  nand n8414(x8414, x8413, x8412);
  nand n8415(x8415, x71210, x8411);
  nand n8416(x8416, x1468, x8414);
  nand n8417(x8417, x8416, x8415);
  nand n8418(x8418, x71202, x3339);
  nand n8419(x8419, x1448, x3209);
  nand n8420(x8420, x8419, x8418);
  nand n8421(x8421, x71202, x3079);
  nand n8422(x8422, x1448, x2949);
  nand n8423(x8423, x8422, x8421);
  nand n8424(x8424, x71202, x2819);
  nand n8425(x8425, x1448, x2689);
  nand n8426(x8426, x8425, x8424);
  nand n8427(x8427, x71202, x2559);
  nand n8428(x8428, x1448, x2429);
  nand n8429(x8429, x8428, x8427);
  nand n8430(x8430, x71205, x8420);
  nand n8431(x8431, x1461, x8423);
  nand n8432(x8432, x8431, x8430);
  nand n8433(x8433, x71205, x8426);
  nand n8434(x8434, x1461, x8429);
  nand n8435(x8435, x8434, x8433);
  nand n8436(x8436, x71210, x8432);
  nand n8437(x8437, x1468, x8435);
  nand n8438(x8438, x8437, x8436);
  nand n8439(x8439, x71202, x3343);
  nand n8440(x8440, x1448, x3213);
  nand n8441(x8441, x8440, x8439);
  nand n8442(x8442, x71202, x3083);
  nand n8443(x8443, x1448, x2953);
  nand n8444(x8444, x8443, x8442);
  nand n8445(x8445, x71202, x2823);
  nand n8446(x8446, x1448, x2693);
  nand n8447(x8447, x8446, x8445);
  nand n8448(x8448, x71202, x2563);
  nand n8449(x8449, x1448, x2433);
  nand n8450(x8450, x8449, x8448);
  nand n8451(x8451, x71205, x8441);
  nand n8452(x8452, x1461, x8444);
  nand n8453(x8453, x8452, x8451);
  nand n8454(x8454, x71205, x8447);
  nand n8455(x8455, x1461, x8450);
  nand n8456(x8456, x8455, x8454);
  nand n8457(x8457, x71210, x8453);
  nand n8458(x8458, x1468, x8456);
  nand n8459(x8459, x8458, x8457);
  nand n8460(x8460, x71202, x3347);
  nand n8461(x8461, x1448, x3217);
  nand n8462(x8462, x8461, x8460);
  nand n8463(x8463, x71202, x3087);
  nand n8464(x8464, x1448, x2957);
  nand n8465(x8465, x8464, x8463);
  nand n8466(x8466, x71202, x2827);
  nand n8467(x8467, x1448, x2697);
  nand n8468(x8468, x8467, x8466);
  nand n8469(x8469, x71202, x2567);
  nand n8470(x8470, x1448, x2437);
  nand n8471(x8471, x8470, x8469);
  nand n8472(x8472, x71205, x8462);
  nand n8473(x8473, x1461, x8465);
  nand n8474(x8474, x8473, x8472);
  nand n8475(x8475, x71205, x8468);
  nand n8476(x8476, x1461, x8471);
  nand n8477(x8477, x8476, x8475);
  nand n8478(x8478, x71210, x8474);
  nand n8479(x8479, x1468, x8477);
  nand n8480(x8480, x8479, x8478);
  nand n8481(x8481, x71202, x3351);
  nand n8482(x8482, x1448, x3221);
  nand n8483(x8483, x8482, x8481);
  nand n8484(x8484, x71202, x3091);
  nand n8485(x8485, x1448, x2961);
  nand n8486(x8486, x8485, x8484);
  nand n8487(x8487, x71202, x2831);
  nand n8488(x8488, x1448, x2701);
  nand n8489(x8489, x8488, x8487);
  nand n8490(x8490, x71202, x2571);
  nand n8491(x8491, x1448, x2441);
  nand n8492(x8492, x8491, x8490);
  nand n8493(x8493, x71205, x8483);
  nand n8494(x8494, x1461, x8486);
  nand n8495(x8495, x8494, x8493);
  nand n8496(x8496, x71205, x8489);
  nand n8497(x8497, x1461, x8492);
  nand n8498(x8498, x8497, x8496);
  nand n8499(x8499, x71210, x8495);
  nand n8500(x8500, x1468, x8498);
  nand n8501(x8501, x8500, x8499);
  nand n8502(x8502, x2258, x4269);
  nand n8503(x8503, x6481, x4139);
  nand n8504(x8504, x8503, x8502);
  nand n8505(x8505, x2258, x4009);
  nand n8506(x8506, x6481, x3879);
  nand n8507(x8507, x8506, x8505);
  nand n8508(x8508, x2258, x3749);
  nand n8509(x8509, x6481, x3619);
  nand n8510(x8510, x8509, x8508);
  nand n8511(x8511, x2258, x3489);
  nand n8512(x8512, x6481, x3359);
  nand n8513(x8513, x8512, x8511);
  nand n8514(x8514, x2261, x8504);
  nand n8515(x8515, x6494, x8507);
  nand n8516(x8516, x8515, x8514);
  nand n8517(x8517, x2261, x8510);
  nand n8518(x8518, x6494, x8513);
  nand n8519(x8519, x8518, x8517);
  nand n8520(x8520, x2264, x8516);
  nand n8521(x8521, x6501, x8519);
  nand n8522(x8522, x8521, x8520);
  nand n8523(x8523, x2258, x4273);
  nand n8524(x8524, x6481, x4143);
  nand n8525(x8525, x8524, x8523);
  nand n8526(x8526, x2258, x4013);
  nand n8527(x8527, x6481, x3883);
  nand n8528(x8528, x8527, x8526);
  nand n8529(x8529, x2258, x3753);
  nand n8530(x8530, x6481, x3623);
  nand n8531(x8531, x8530, x8529);
  nand n8532(x8532, x2258, x3493);
  nand n8533(x8533, x6481, x3363);
  nand n8534(x8534, x8533, x8532);
  nand n8535(x8535, x2261, x8525);
  nand n8536(x8536, x6494, x8528);
  nand n8537(x8537, x8536, x8535);
  nand n8538(x8538, x2261, x8531);
  nand n8539(x8539, x6494, x8534);
  nand n8540(x8540, x8539, x8538);
  nand n8541(x8541, x2264, x8537);
  nand n8542(x8542, x6501, x8540);
  nand n8543(x8543, x8542, x8541);
  nand n8544(x8544, x2258, x4277);
  nand n8545(x8545, x6481, x4147);
  nand n8546(x8546, x8545, x8544);
  nand n8547(x8547, x2258, x4017);
  nand n8548(x8548, x6481, x3887);
  nand n8549(x8549, x8548, x8547);
  nand n8550(x8550, x2258, x3757);
  nand n8551(x8551, x6481, x3627);
  nand n8552(x8552, x8551, x8550);
  nand n8553(x8553, x2258, x3497);
  nand n8554(x8554, x6481, x3367);
  nand n8555(x8555, x8554, x8553);
  nand n8556(x8556, x2261, x8546);
  nand n8557(x8557, x6494, x8549);
  nand n8558(x8558, x8557, x8556);
  nand n8559(x8559, x2261, x8552);
  nand n8560(x8560, x6494, x8555);
  nand n8561(x8561, x8560, x8559);
  nand n8562(x8562, x2264, x8558);
  nand n8563(x8563, x6501, x8561);
  nand n8564(x8564, x8563, x8562);
  nand n8565(x8565, x2258, x4281);
  nand n8566(x8566, x6481, x4151);
  nand n8567(x8567, x8566, x8565);
  nand n8568(x8568, x2258, x4021);
  nand n8569(x8569, x6481, x3891);
  nand n8570(x8570, x8569, x8568);
  nand n8571(x8571, x2258, x3761);
  nand n8572(x8572, x6481, x3631);
  nand n8573(x8573, x8572, x8571);
  nand n8574(x8574, x2258, x3501);
  nand n8575(x8575, x6481, x3371);
  nand n8576(x8576, x8575, x8574);
  nand n8577(x8577, x2261, x8567);
  nand n8578(x8578, x6494, x8570);
  nand n8579(x8579, x8578, x8577);
  nand n8580(x8580, x2261, x8573);
  nand n8581(x8581, x6494, x8576);
  nand n8582(x8582, x8581, x8580);
  nand n8583(x8583, x2264, x8579);
  nand n8584(x8584, x6501, x8582);
  nand n8585(x8585, x8584, x8583);
  nand n8586(x8586, x2258, x4285);
  nand n8587(x8587, x6481, x4155);
  nand n8588(x8588, x8587, x8586);
  nand n8589(x8589, x2258, x4025);
  nand n8590(x8590, x6481, x3895);
  nand n8591(x8591, x8590, x8589);
  nand n8592(x8592, x2258, x3765);
  nand n8593(x8593, x6481, x3635);
  nand n8594(x8594, x8593, x8592);
  nand n8595(x8595, x2258, x3505);
  nand n8596(x8596, x6481, x3375);
  nand n8597(x8597, x8596, x8595);
  nand n8598(x8598, x2261, x8588);
  nand n8599(x8599, x6494, x8591);
  nand n8600(x8600, x8599, x8598);
  nand n8601(x8601, x2261, x8594);
  nand n8602(x8602, x6494, x8597);
  nand n8603(x8603, x8602, x8601);
  nand n8604(x8604, x2264, x8600);
  nand n8605(x8605, x6501, x8603);
  nand n8606(x8606, x8605, x8604);
  nand n8607(x8607, x2258, x4289);
  nand n8608(x8608, x6481, x4159);
  nand n8609(x8609, x8608, x8607);
  nand n8610(x8610, x2258, x4029);
  nand n8611(x8611, x6481, x3899);
  nand n8612(x8612, x8611, x8610);
  nand n8613(x8613, x2258, x3769);
  nand n8614(x8614, x6481, x3639);
  nand n8615(x8615, x8614, x8613);
  nand n8616(x8616, x2258, x3509);
  nand n8617(x8617, x6481, x3379);
  nand n8618(x8618, x8617, x8616);
  nand n8619(x8619, x2261, x8609);
  nand n8620(x8620, x6494, x8612);
  nand n8621(x8621, x8620, x8619);
  nand n8622(x8622, x2261, x8615);
  nand n8623(x8623, x6494, x8618);
  nand n8624(x8624, x8623, x8622);
  nand n8625(x8625, x2264, x8621);
  nand n8626(x8626, x6501, x8624);
  nand n8627(x8627, x8626, x8625);
  nand n8628(x8628, x2258, x4293);
  nand n8629(x8629, x6481, x4163);
  nand n8630(x8630, x8629, x8628);
  nand n8631(x8631, x2258, x4033);
  nand n8632(x8632, x6481, x3903);
  nand n8633(x8633, x8632, x8631);
  nand n8634(x8634, x2258, x3773);
  nand n8635(x8635, x6481, x3643);
  nand n8636(x8636, x8635, x8634);
  nand n8637(x8637, x2258, x3513);
  nand n8638(x8638, x6481, x3383);
  nand n8639(x8639, x8638, x8637);
  nand n8640(x8640, x2261, x8630);
  nand n8641(x8641, x6494, x8633);
  nand n8642(x8642, x8641, x8640);
  nand n8643(x8643, x2261, x8636);
  nand n8644(x8644, x6494, x8639);
  nand n8645(x8645, x8644, x8643);
  nand n8646(x8646, x2264, x8642);
  nand n8647(x8647, x6501, x8645);
  nand n8648(x8648, x8647, x8646);
  nand n8649(x8649, x2258, x4297);
  nand n8650(x8650, x6481, x4167);
  nand n8651(x8651, x8650, x8649);
  nand n8652(x8652, x2258, x4037);
  nand n8653(x8653, x6481, x3907);
  nand n8654(x8654, x8653, x8652);
  nand n8655(x8655, x2258, x3777);
  nand n8656(x8656, x6481, x3647);
  nand n8657(x8657, x8656, x8655);
  nand n8658(x8658, x2258, x3517);
  nand n8659(x8659, x6481, x3387);
  nand n8660(x8660, x8659, x8658);
  nand n8661(x8661, x2261, x8651);
  nand n8662(x8662, x6494, x8654);
  nand n8663(x8663, x8662, x8661);
  nand n8664(x8664, x2261, x8657);
  nand n8665(x8665, x6494, x8660);
  nand n8666(x8666, x8665, x8664);
  nand n8667(x8667, x2264, x8663);
  nand n8668(x8668, x6501, x8666);
  nand n8669(x8669, x8668, x8667);
  nand n8670(x8670, x2258, x4301);
  nand n8671(x8671, x6481, x4171);
  nand n8672(x8672, x8671, x8670);
  nand n8673(x8673, x2258, x4041);
  nand n8674(x8674, x6481, x3911);
  nand n8675(x8675, x8674, x8673);
  nand n8676(x8676, x2258, x3781);
  nand n8677(x8677, x6481, x3651);
  nand n8678(x8678, x8677, x8676);
  nand n8679(x8679, x2258, x3521);
  nand n8680(x8680, x6481, x3391);
  nand n8681(x8681, x8680, x8679);
  nand n8682(x8682, x2261, x8672);
  nand n8683(x8683, x6494, x8675);
  nand n8684(x8684, x8683, x8682);
  nand n8685(x8685, x2261, x8678);
  nand n8686(x8686, x6494, x8681);
  nand n8687(x8687, x8686, x8685);
  nand n8688(x8688, x2264, x8684);
  nand n8689(x8689, x6501, x8687);
  nand n8690(x8690, x8689, x8688);
  nand n8691(x8691, x2258, x4305);
  nand n8692(x8692, x6481, x4175);
  nand n8693(x8693, x8692, x8691);
  nand n8694(x8694, x2258, x4045);
  nand n8695(x8695, x6481, x3915);
  nand n8696(x8696, x8695, x8694);
  nand n8697(x8697, x2258, x3785);
  nand n8698(x8698, x6481, x3655);
  nand n8699(x8699, x8698, x8697);
  nand n8700(x8700, x2258, x3525);
  nand n8701(x8701, x6481, x3395);
  nand n8702(x8702, x8701, x8700);
  nand n8703(x8703, x2261, x8693);
  nand n8704(x8704, x6494, x8696);
  nand n8705(x8705, x8704, x8703);
  nand n8706(x8706, x2261, x8699);
  nand n8707(x8707, x6494, x8702);
  nand n8708(x8708, x8707, x8706);
  nand n8709(x8709, x2264, x8705);
  nand n8710(x8710, x6501, x8708);
  nand n8711(x8711, x8710, x8709);
  nand n8712(x8712, x2258, x4309);
  nand n8713(x8713, x6481, x4179);
  nand n8714(x8714, x8713, x8712);
  nand n8715(x8715, x2258, x4049);
  nand n8716(x8716, x6481, x3919);
  nand n8717(x8717, x8716, x8715);
  nand n8718(x8718, x2258, x3789);
  nand n8719(x8719, x6481, x3659);
  nand n8720(x8720, x8719, x8718);
  nand n8721(x8721, x2258, x3529);
  nand n8722(x8722, x6481, x3399);
  nand n8723(x8723, x8722, x8721);
  nand n8724(x8724, x2261, x8714);
  nand n8725(x8725, x6494, x8717);
  nand n8726(x8726, x8725, x8724);
  nand n8727(x8727, x2261, x8720);
  nand n8728(x8728, x6494, x8723);
  nand n8729(x8729, x8728, x8727);
  nand n8730(x8730, x2264, x8726);
  nand n8731(x8731, x6501, x8729);
  nand n8732(x8732, x8731, x8730);
  nand n8733(x8733, x2258, x4313);
  nand n8734(x8734, x6481, x4183);
  nand n8735(x8735, x8734, x8733);
  nand n8736(x8736, x2258, x4053);
  nand n8737(x8737, x6481, x3923);
  nand n8738(x8738, x8737, x8736);
  nand n8739(x8739, x2258, x3793);
  nand n8740(x8740, x6481, x3663);
  nand n8741(x8741, x8740, x8739);
  nand n8742(x8742, x2258, x3533);
  nand n8743(x8743, x6481, x3403);
  nand n8744(x8744, x8743, x8742);
  nand n8745(x8745, x2261, x8735);
  nand n8746(x8746, x6494, x8738);
  nand n8747(x8747, x8746, x8745);
  nand n8748(x8748, x2261, x8741);
  nand n8749(x8749, x6494, x8744);
  nand n8750(x8750, x8749, x8748);
  nand n8751(x8751, x2264, x8747);
  nand n8752(x8752, x6501, x8750);
  nand n8753(x8753, x8752, x8751);
  nand n8754(x8754, x2258, x4317);
  nand n8755(x8755, x6481, x4187);
  nand n8756(x8756, x8755, x8754);
  nand n8757(x8757, x2258, x4057);
  nand n8758(x8758, x6481, x3927);
  nand n8759(x8759, x8758, x8757);
  nand n8760(x8760, x2258, x3797);
  nand n8761(x8761, x6481, x3667);
  nand n8762(x8762, x8761, x8760);
  nand n8763(x8763, x2258, x3537);
  nand n8764(x8764, x6481, x3407);
  nand n8765(x8765, x8764, x8763);
  nand n8766(x8766, x2261, x8756);
  nand n8767(x8767, x6494, x8759);
  nand n8768(x8768, x8767, x8766);
  nand n8769(x8769, x2261, x8762);
  nand n8770(x8770, x6494, x8765);
  nand n8771(x8771, x8770, x8769);
  nand n8772(x8772, x2264, x8768);
  nand n8773(x8773, x6501, x8771);
  nand n8774(x8774, x8773, x8772);
  nand n8775(x8775, x2258, x4321);
  nand n8776(x8776, x6481, x4191);
  nand n8777(x8777, x8776, x8775);
  nand n8778(x8778, x2258, x4061);
  nand n8779(x8779, x6481, x3931);
  nand n8780(x8780, x8779, x8778);
  nand n8781(x8781, x2258, x3801);
  nand n8782(x8782, x6481, x3671);
  nand n8783(x8783, x8782, x8781);
  nand n8784(x8784, x2258, x3541);
  nand n8785(x8785, x6481, x3411);
  nand n8786(x8786, x8785, x8784);
  nand n8787(x8787, x2261, x8777);
  nand n8788(x8788, x6494, x8780);
  nand n8789(x8789, x8788, x8787);
  nand n8790(x8790, x2261, x8783);
  nand n8791(x8791, x6494, x8786);
  nand n8792(x8792, x8791, x8790);
  nand n8793(x8793, x2264, x8789);
  nand n8794(x8794, x6501, x8792);
  nand n8795(x8795, x8794, x8793);
  nand n8796(x8796, x2258, x4325);
  nand n8797(x8797, x6481, x4195);
  nand n8798(x8798, x8797, x8796);
  nand n8799(x8799, x2258, x4065);
  nand n8800(x8800, x6481, x3935);
  nand n8801(x8801, x8800, x8799);
  nand n8802(x8802, x2258, x3805);
  nand n8803(x8803, x6481, x3675);
  nand n8804(x8804, x8803, x8802);
  nand n8805(x8805, x2258, x3545);
  nand n8806(x8806, x6481, x3415);
  nand n8807(x8807, x8806, x8805);
  nand n8808(x8808, x2261, x8798);
  nand n8809(x8809, x6494, x8801);
  nand n8810(x8810, x8809, x8808);
  nand n8811(x8811, x2261, x8804);
  nand n8812(x8812, x6494, x8807);
  nand n8813(x8813, x8812, x8811);
  nand n8814(x8814, x2264, x8810);
  nand n8815(x8815, x6501, x8813);
  nand n8816(x8816, x8815, x8814);
  nand n8817(x8817, x2258, x4329);
  nand n8818(x8818, x6481, x4199);
  nand n8819(x8819, x8818, x8817);
  nand n8820(x8820, x2258, x4069);
  nand n8821(x8821, x6481, x3939);
  nand n8822(x8822, x8821, x8820);
  nand n8823(x8823, x2258, x3809);
  nand n8824(x8824, x6481, x3679);
  nand n8825(x8825, x8824, x8823);
  nand n8826(x8826, x2258, x3549);
  nand n8827(x8827, x6481, x3419);
  nand n8828(x8828, x8827, x8826);
  nand n8829(x8829, x2261, x8819);
  nand n8830(x8830, x6494, x8822);
  nand n8831(x8831, x8830, x8829);
  nand n8832(x8832, x2261, x8825);
  nand n8833(x8833, x6494, x8828);
  nand n8834(x8834, x8833, x8832);
  nand n8835(x8835, x2264, x8831);
  nand n8836(x8836, x6501, x8834);
  nand n8837(x8837, x8836, x8835);
  nand n8838(x8838, x2258, x4333);
  nand n8839(x8839, x6481, x4203);
  nand n8840(x8840, x8839, x8838);
  nand n8841(x8841, x2258, x4073);
  nand n8842(x8842, x6481, x3943);
  nand n8843(x8843, x8842, x8841);
  nand n8844(x8844, x2258, x3813);
  nand n8845(x8845, x6481, x3683);
  nand n8846(x8846, x8845, x8844);
  nand n8847(x8847, x2258, x3553);
  nand n8848(x8848, x6481, x3423);
  nand n8849(x8849, x8848, x8847);
  nand n8850(x8850, x2261, x8840);
  nand n8851(x8851, x6494, x8843);
  nand n8852(x8852, x8851, x8850);
  nand n8853(x8853, x2261, x8846);
  nand n8854(x8854, x6494, x8849);
  nand n8855(x8855, x8854, x8853);
  nand n8856(x8856, x2264, x8852);
  nand n8857(x8857, x6501, x8855);
  nand n8858(x8858, x8857, x8856);
  nand n8859(x8859, x2258, x4337);
  nand n8860(x8860, x6481, x4207);
  nand n8861(x8861, x8860, x8859);
  nand n8862(x8862, x2258, x4077);
  nand n8863(x8863, x6481, x3947);
  nand n8864(x8864, x8863, x8862);
  nand n8865(x8865, x2258, x3817);
  nand n8866(x8866, x6481, x3687);
  nand n8867(x8867, x8866, x8865);
  nand n8868(x8868, x2258, x3557);
  nand n8869(x8869, x6481, x3427);
  nand n8870(x8870, x8869, x8868);
  nand n8871(x8871, x2261, x8861);
  nand n8872(x8872, x6494, x8864);
  nand n8873(x8873, x8872, x8871);
  nand n8874(x8874, x2261, x8867);
  nand n8875(x8875, x6494, x8870);
  nand n8876(x8876, x8875, x8874);
  nand n8877(x8877, x2264, x8873);
  nand n8878(x8878, x6501, x8876);
  nand n8879(x8879, x8878, x8877);
  nand n8880(x8880, x2258, x4341);
  nand n8881(x8881, x6481, x4211);
  nand n8882(x8882, x8881, x8880);
  nand n8883(x8883, x2258, x4081);
  nand n8884(x8884, x6481, x3951);
  nand n8885(x8885, x8884, x8883);
  nand n8886(x8886, x2258, x3821);
  nand n8887(x8887, x6481, x3691);
  nand n8888(x8888, x8887, x8886);
  nand n8889(x8889, x2258, x3561);
  nand n8890(x8890, x6481, x3431);
  nand n8891(x8891, x8890, x8889);
  nand n8892(x8892, x2261, x8882);
  nand n8893(x8893, x6494, x8885);
  nand n8894(x8894, x8893, x8892);
  nand n8895(x8895, x2261, x8888);
  nand n8896(x8896, x6494, x8891);
  nand n8897(x8897, x8896, x8895);
  nand n8898(x8898, x2264, x8894);
  nand n8899(x8899, x6501, x8897);
  nand n8900(x8900, x8899, x8898);
  nand n8901(x8901, x2258, x4345);
  nand n8902(x8902, x6481, x4215);
  nand n8903(x8903, x8902, x8901);
  nand n8904(x8904, x2258, x4085);
  nand n8905(x8905, x6481, x3955);
  nand n8906(x8906, x8905, x8904);
  nand n8907(x8907, x2258, x3825);
  nand n8908(x8908, x6481, x3695);
  nand n8909(x8909, x8908, x8907);
  nand n8910(x8910, x2258, x3565);
  nand n8911(x8911, x6481, x3435);
  nand n8912(x8912, x8911, x8910);
  nand n8913(x8913, x2261, x8903);
  nand n8914(x8914, x6494, x8906);
  nand n8915(x8915, x8914, x8913);
  nand n8916(x8916, x2261, x8909);
  nand n8917(x8917, x6494, x8912);
  nand n8918(x8918, x8917, x8916);
  nand n8919(x8919, x2264, x8915);
  nand n8920(x8920, x6501, x8918);
  nand n8921(x8921, x8920, x8919);
  nand n8922(x8922, x2258, x4349);
  nand n8923(x8923, x6481, x4219);
  nand n8924(x8924, x8923, x8922);
  nand n8925(x8925, x2258, x4089);
  nand n8926(x8926, x6481, x3959);
  nand n8927(x8927, x8926, x8925);
  nand n8928(x8928, x2258, x3829);
  nand n8929(x8929, x6481, x3699);
  nand n8930(x8930, x8929, x8928);
  nand n8931(x8931, x2258, x3569);
  nand n8932(x8932, x6481, x3439);
  nand n8933(x8933, x8932, x8931);
  nand n8934(x8934, x2261, x8924);
  nand n8935(x8935, x6494, x8927);
  nand n8936(x8936, x8935, x8934);
  nand n8937(x8937, x2261, x8930);
  nand n8938(x8938, x6494, x8933);
  nand n8939(x8939, x8938, x8937);
  nand n8940(x8940, x2264, x8936);
  nand n8941(x8941, x6501, x8939);
  nand n8942(x8942, x8941, x8940);
  nand n8943(x8943, x2258, x4353);
  nand n8944(x8944, x6481, x4223);
  nand n8945(x8945, x8944, x8943);
  nand n8946(x8946, x2258, x4093);
  nand n8947(x8947, x6481, x3963);
  nand n8948(x8948, x8947, x8946);
  nand n8949(x8949, x2258, x3833);
  nand n8950(x8950, x6481, x3703);
  nand n8951(x8951, x8950, x8949);
  nand n8952(x8952, x2258, x3573);
  nand n8953(x8953, x6481, x3443);
  nand n8954(x8954, x8953, x8952);
  nand n8955(x8955, x2261, x8945);
  nand n8956(x8956, x6494, x8948);
  nand n8957(x8957, x8956, x8955);
  nand n8958(x8958, x2261, x8951);
  nand n8959(x8959, x6494, x8954);
  nand n8960(x8960, x8959, x8958);
  nand n8961(x8961, x2264, x8957);
  nand n8962(x8962, x6501, x8960);
  nand n8963(x8963, x8962, x8961);
  nand n8964(x8964, x2258, x4357);
  nand n8965(x8965, x6481, x4227);
  nand n8966(x8966, x8965, x8964);
  nand n8967(x8967, x2258, x4097);
  nand n8968(x8968, x6481, x3967);
  nand n8969(x8969, x8968, x8967);
  nand n8970(x8970, x2258, x3837);
  nand n8971(x8971, x6481, x3707);
  nand n8972(x8972, x8971, x8970);
  nand n8973(x8973, x2258, x3577);
  nand n8974(x8974, x6481, x3447);
  nand n8975(x8975, x8974, x8973);
  nand n8976(x8976, x2261, x8966);
  nand n8977(x8977, x6494, x8969);
  nand n8978(x8978, x8977, x8976);
  nand n8979(x8979, x2261, x8972);
  nand n8980(x8980, x6494, x8975);
  nand n8981(x8981, x8980, x8979);
  nand n8982(x8982, x2264, x8978);
  nand n8983(x8983, x6501, x8981);
  nand n8984(x8984, x8983, x8982);
  nand n8985(x8985, x2258, x4361);
  nand n8986(x8986, x6481, x4231);
  nand n8987(x8987, x8986, x8985);
  nand n8988(x8988, x2258, x4101);
  nand n8989(x8989, x6481, x3971);
  nand n8990(x8990, x8989, x8988);
  nand n8991(x8991, x2258, x3841);
  nand n8992(x8992, x6481, x3711);
  nand n8993(x8993, x8992, x8991);
  nand n8994(x8994, x2258, x3581);
  nand n8995(x8995, x6481, x3451);
  nand n8996(x8996, x8995, x8994);
  nand n8997(x8997, x2261, x8987);
  nand n8998(x8998, x6494, x8990);
  nand n8999(x8999, x8998, x8997);
  nand n9000(x9000, x2261, x8993);
  nand n9001(x9001, x6494, x8996);
  nand n9002(x9002, x9001, x9000);
  nand n9003(x9003, x2264, x8999);
  nand n9004(x9004, x6501, x9002);
  nand n9005(x9005, x9004, x9003);
  nand n9006(x9006, x2258, x4365);
  nand n9007(x9007, x6481, x4235);
  nand n9008(x9008, x9007, x9006);
  nand n9009(x9009, x2258, x4105);
  nand n9010(x9010, x6481, x3975);
  nand n9011(x9011, x9010, x9009);
  nand n9012(x9012, x2258, x3845);
  nand n9013(x9013, x6481, x3715);
  nand n9014(x9014, x9013, x9012);
  nand n9015(x9015, x2258, x3585);
  nand n9016(x9016, x6481, x3455);
  nand n9017(x9017, x9016, x9015);
  nand n9018(x9018, x2261, x9008);
  nand n9019(x9019, x6494, x9011);
  nand n9020(x9020, x9019, x9018);
  nand n9021(x9021, x2261, x9014);
  nand n9022(x9022, x6494, x9017);
  nand n9023(x9023, x9022, x9021);
  nand n9024(x9024, x2264, x9020);
  nand n9025(x9025, x6501, x9023);
  nand n9026(x9026, x9025, x9024);
  nand n9027(x9027, x2258, x4369);
  nand n9028(x9028, x6481, x4239);
  nand n9029(x9029, x9028, x9027);
  nand n9030(x9030, x2258, x4109);
  nand n9031(x9031, x6481, x3979);
  nand n9032(x9032, x9031, x9030);
  nand n9033(x9033, x2258, x3849);
  nand n9034(x9034, x6481, x3719);
  nand n9035(x9035, x9034, x9033);
  nand n9036(x9036, x2258, x3589);
  nand n9037(x9037, x6481, x3459);
  nand n9038(x9038, x9037, x9036);
  nand n9039(x9039, x2261, x9029);
  nand n9040(x9040, x6494, x9032);
  nand n9041(x9041, x9040, x9039);
  nand n9042(x9042, x2261, x9035);
  nand n9043(x9043, x6494, x9038);
  nand n9044(x9044, x9043, x9042);
  nand n9045(x9045, x2264, x9041);
  nand n9046(x9046, x6501, x9044);
  nand n9047(x9047, x9046, x9045);
  nand n9048(x9048, x2258, x4373);
  nand n9049(x9049, x6481, x4243);
  nand n9050(x9050, x9049, x9048);
  nand n9051(x9051, x2258, x4113);
  nand n9052(x9052, x6481, x3983);
  nand n9053(x9053, x9052, x9051);
  nand n9054(x9054, x2258, x3853);
  nand n9055(x9055, x6481, x3723);
  nand n9056(x9056, x9055, x9054);
  nand n9057(x9057, x2258, x3593);
  nand n9058(x9058, x6481, x3463);
  nand n9059(x9059, x9058, x9057);
  nand n9060(x9060, x2261, x9050);
  nand n9061(x9061, x6494, x9053);
  nand n9062(x9062, x9061, x9060);
  nand n9063(x9063, x2261, x9056);
  nand n9064(x9064, x6494, x9059);
  nand n9065(x9065, x9064, x9063);
  nand n9066(x9066, x2264, x9062);
  nand n9067(x9067, x6501, x9065);
  nand n9068(x9068, x9067, x9066);
  nand n9069(x9069, x2258, x4377);
  nand n9070(x9070, x6481, x4247);
  nand n9071(x9071, x9070, x9069);
  nand n9072(x9072, x2258, x4117);
  nand n9073(x9073, x6481, x3987);
  nand n9074(x9074, x9073, x9072);
  nand n9075(x9075, x2258, x3857);
  nand n9076(x9076, x6481, x3727);
  nand n9077(x9077, x9076, x9075);
  nand n9078(x9078, x2258, x3597);
  nand n9079(x9079, x6481, x3467);
  nand n9080(x9080, x9079, x9078);
  nand n9081(x9081, x2261, x9071);
  nand n9082(x9082, x6494, x9074);
  nand n9083(x9083, x9082, x9081);
  nand n9084(x9084, x2261, x9077);
  nand n9085(x9085, x6494, x9080);
  nand n9086(x9086, x9085, x9084);
  nand n9087(x9087, x2264, x9083);
  nand n9088(x9088, x6501, x9086);
  nand n9089(x9089, x9088, x9087);
  nand n9090(x9090, x2258, x4381);
  nand n9091(x9091, x6481, x4251);
  nand n9092(x9092, x9091, x9090);
  nand n9093(x9093, x2258, x4121);
  nand n9094(x9094, x6481, x3991);
  nand n9095(x9095, x9094, x9093);
  nand n9096(x9096, x2258, x3861);
  nand n9097(x9097, x6481, x3731);
  nand n9098(x9098, x9097, x9096);
  nand n9099(x9099, x2258, x3601);
  nand n9100(x9100, x6481, x3471);
  nand n9101(x9101, x9100, x9099);
  nand n9102(x9102, x2261, x9092);
  nand n9103(x9103, x6494, x9095);
  nand n9104(x9104, x9103, x9102);
  nand n9105(x9105, x2261, x9098);
  nand n9106(x9106, x6494, x9101);
  nand n9107(x9107, x9106, x9105);
  nand n9108(x9108, x2264, x9104);
  nand n9109(x9109, x6501, x9107);
  nand n9110(x9110, x9109, x9108);
  nand n9111(x9111, x2258, x4385);
  nand n9112(x9112, x6481, x4255);
  nand n9113(x9113, x9112, x9111);
  nand n9114(x9114, x2258, x4125);
  nand n9115(x9115, x6481, x3995);
  nand n9116(x9116, x9115, x9114);
  nand n9117(x9117, x2258, x3865);
  nand n9118(x9118, x6481, x3735);
  nand n9119(x9119, x9118, x9117);
  nand n9120(x9120, x2258, x3605);
  nand n9121(x9121, x6481, x3475);
  nand n9122(x9122, x9121, x9120);
  nand n9123(x9123, x2261, x9113);
  nand n9124(x9124, x6494, x9116);
  nand n9125(x9125, x9124, x9123);
  nand n9126(x9126, x2261, x9119);
  nand n9127(x9127, x6494, x9122);
  nand n9128(x9128, x9127, x9126);
  nand n9129(x9129, x2264, x9125);
  nand n9130(x9130, x6501, x9128);
  nand n9131(x9131, x9130, x9129);
  nand n9132(x9132, x2258, x4389);
  nand n9133(x9133, x6481, x4259);
  nand n9134(x9134, x9133, x9132);
  nand n9135(x9135, x2258, x4129);
  nand n9136(x9136, x6481, x3999);
  nand n9137(x9137, x9136, x9135);
  nand n9138(x9138, x2258, x3869);
  nand n9139(x9139, x6481, x3739);
  nand n9140(x9140, x9139, x9138);
  nand n9141(x9141, x2258, x3609);
  nand n9142(x9142, x6481, x3479);
  nand n9143(x9143, x9142, x9141);
  nand n9144(x9144, x2261, x9134);
  nand n9145(x9145, x6494, x9137);
  nand n9146(x9146, x9145, x9144);
  nand n9147(x9147, x2261, x9140);
  nand n9148(x9148, x6494, x9143);
  nand n9149(x9149, x9148, x9147);
  nand n9150(x9150, x2264, x9146);
  nand n9151(x9151, x6501, x9149);
  nand n9152(x9152, x9151, x9150);
  nand n9153(x9153, x2258, x4393);
  nand n9154(x9154, x6481, x4263);
  nand n9155(x9155, x9154, x9153);
  nand n9156(x9156, x2258, x4133);
  nand n9157(x9157, x6481, x4003);
  nand n9158(x9158, x9157, x9156);
  nand n9159(x9159, x2258, x3873);
  nand n9160(x9160, x6481, x3743);
  nand n9161(x9161, x9160, x9159);
  nand n9162(x9162, x2258, x3613);
  nand n9163(x9163, x6481, x3483);
  nand n9164(x9164, x9163, x9162);
  nand n9165(x9165, x2261, x9155);
  nand n9166(x9166, x6494, x9158);
  nand n9167(x9167, x9166, x9165);
  nand n9168(x9168, x2261, x9161);
  nand n9169(x9169, x6494, x9164);
  nand n9170(x9170, x9169, x9168);
  nand n9171(x9171, x2264, x9167);
  nand n9172(x9172, x6501, x9170);
  nand n9173(x9173, x9172, x9171);
  nand n9174(x9174, x2269, x4269);
  nand n9175(x9175, x7156, x4139);
  nand n9176(x9176, x9175, x9174);
  nand n9177(x9177, x2269, x4009);
  nand n9178(x9178, x7156, x3879);
  nand n9179(x9179, x9178, x9177);
  nand n9180(x9180, x2269, x3749);
  nand n9181(x9181, x7156, x3619);
  nand n9182(x9182, x9181, x9180);
  nand n9183(x9183, x2269, x3489);
  nand n9184(x9184, x7156, x3359);
  nand n9185(x9185, x9184, x9183);
  nand n9186(x9186, x2272, x9176);
  nand n9187(x9187, x7169, x9179);
  nand n9188(x9188, x9187, x9186);
  nand n9189(x9189, x2272, x9182);
  nand n9190(x9190, x7169, x9185);
  nand n9191(x9191, x9190, x9189);
  nand n9192(x9192, x2275, x9188);
  nand n9193(x9193, x7176, x9191);
  nand n9194(x9194, x9193, x9192);
  nand n9195(x9195, x2269, x4273);
  nand n9196(x9196, x7156, x4143);
  nand n9197(x9197, x9196, x9195);
  nand n9198(x9198, x2269, x4013);
  nand n9199(x9199, x7156, x3883);
  nand n9200(x9200, x9199, x9198);
  nand n9201(x9201, x2269, x3753);
  nand n9202(x9202, x7156, x3623);
  nand n9203(x9203, x9202, x9201);
  nand n9204(x9204, x2269, x3493);
  nand n9205(x9205, x7156, x3363);
  nand n9206(x9206, x9205, x9204);
  nand n9207(x9207, x2272, x9197);
  nand n9208(x9208, x7169, x9200);
  nand n9209(x9209, x9208, x9207);
  nand n9210(x9210, x2272, x9203);
  nand n9211(x9211, x7169, x9206);
  nand n9212(x9212, x9211, x9210);
  nand n9213(x9213, x2275, x9209);
  nand n9214(x9214, x7176, x9212);
  nand n9215(x9215, x9214, x9213);
  nand n9216(x9216, x2269, x4277);
  nand n9217(x9217, x7156, x4147);
  nand n9218(x9218, x9217, x9216);
  nand n9219(x9219, x2269, x4017);
  nand n9220(x9220, x7156, x3887);
  nand n9221(x9221, x9220, x9219);
  nand n9222(x9222, x2269, x3757);
  nand n9223(x9223, x7156, x3627);
  nand n9224(x9224, x9223, x9222);
  nand n9225(x9225, x2269, x3497);
  nand n9226(x9226, x7156, x3367);
  nand n9227(x9227, x9226, x9225);
  nand n9228(x9228, x2272, x9218);
  nand n9229(x9229, x7169, x9221);
  nand n9230(x9230, x9229, x9228);
  nand n9231(x9231, x2272, x9224);
  nand n9232(x9232, x7169, x9227);
  nand n9233(x9233, x9232, x9231);
  nand n9234(x9234, x2275, x9230);
  nand n9235(x9235, x7176, x9233);
  nand n9236(x9236, x9235, x9234);
  nand n9237(x9237, x2269, x4281);
  nand n9238(x9238, x7156, x4151);
  nand n9239(x9239, x9238, x9237);
  nand n9240(x9240, x2269, x4021);
  nand n9241(x9241, x7156, x3891);
  nand n9242(x9242, x9241, x9240);
  nand n9243(x9243, x2269, x3761);
  nand n9244(x9244, x7156, x3631);
  nand n9245(x9245, x9244, x9243);
  nand n9246(x9246, x2269, x3501);
  nand n9247(x9247, x7156, x3371);
  nand n9248(x9248, x9247, x9246);
  nand n9249(x9249, x2272, x9239);
  nand n9250(x9250, x7169, x9242);
  nand n9251(x9251, x9250, x9249);
  nand n9252(x9252, x2272, x9245);
  nand n9253(x9253, x7169, x9248);
  nand n9254(x9254, x9253, x9252);
  nand n9255(x9255, x2275, x9251);
  nand n9256(x9256, x7176, x9254);
  nand n9257(x9257, x9256, x9255);
  nand n9258(x9258, x2269, x4285);
  nand n9259(x9259, x7156, x4155);
  nand n9260(x9260, x9259, x9258);
  nand n9261(x9261, x2269, x4025);
  nand n9262(x9262, x7156, x3895);
  nand n9263(x9263, x9262, x9261);
  nand n9264(x9264, x2269, x3765);
  nand n9265(x9265, x7156, x3635);
  nand n9266(x9266, x9265, x9264);
  nand n9267(x9267, x2269, x3505);
  nand n9268(x9268, x7156, x3375);
  nand n9269(x9269, x9268, x9267);
  nand n9270(x9270, x2272, x9260);
  nand n9271(x9271, x7169, x9263);
  nand n9272(x9272, x9271, x9270);
  nand n9273(x9273, x2272, x9266);
  nand n9274(x9274, x7169, x9269);
  nand n9275(x9275, x9274, x9273);
  nand n9276(x9276, x2275, x9272);
  nand n9277(x9277, x7176, x9275);
  nand n9278(x9278, x9277, x9276);
  nand n9279(x9279, x2269, x4289);
  nand n9280(x9280, x7156, x4159);
  nand n9281(x9281, x9280, x9279);
  nand n9282(x9282, x2269, x4029);
  nand n9283(x9283, x7156, x3899);
  nand n9284(x9284, x9283, x9282);
  nand n9285(x9285, x2269, x3769);
  nand n9286(x9286, x7156, x3639);
  nand n9287(x9287, x9286, x9285);
  nand n9288(x9288, x2269, x3509);
  nand n9289(x9289, x7156, x3379);
  nand n9290(x9290, x9289, x9288);
  nand n9291(x9291, x2272, x9281);
  nand n9292(x9292, x7169, x9284);
  nand n9293(x9293, x9292, x9291);
  nand n9294(x9294, x2272, x9287);
  nand n9295(x9295, x7169, x9290);
  nand n9296(x9296, x9295, x9294);
  nand n9297(x9297, x2275, x9293);
  nand n9298(x9298, x7176, x9296);
  nand n9299(x9299, x9298, x9297);
  nand n9300(x9300, x2269, x4293);
  nand n9301(x9301, x7156, x4163);
  nand n9302(x9302, x9301, x9300);
  nand n9303(x9303, x2269, x4033);
  nand n9304(x9304, x7156, x3903);
  nand n9305(x9305, x9304, x9303);
  nand n9306(x9306, x2269, x3773);
  nand n9307(x9307, x7156, x3643);
  nand n9308(x9308, x9307, x9306);
  nand n9309(x9309, x2269, x3513);
  nand n9310(x9310, x7156, x3383);
  nand n9311(x9311, x9310, x9309);
  nand n9312(x9312, x2272, x9302);
  nand n9313(x9313, x7169, x9305);
  nand n9314(x9314, x9313, x9312);
  nand n9315(x9315, x2272, x9308);
  nand n9316(x9316, x7169, x9311);
  nand n9317(x9317, x9316, x9315);
  nand n9318(x9318, x2275, x9314);
  nand n9319(x9319, x7176, x9317);
  nand n9320(x9320, x9319, x9318);
  nand n9321(x9321, x2269, x4297);
  nand n9322(x9322, x7156, x4167);
  nand n9323(x9323, x9322, x9321);
  nand n9324(x9324, x2269, x4037);
  nand n9325(x9325, x7156, x3907);
  nand n9326(x9326, x9325, x9324);
  nand n9327(x9327, x2269, x3777);
  nand n9328(x9328, x7156, x3647);
  nand n9329(x9329, x9328, x9327);
  nand n9330(x9330, x2269, x3517);
  nand n9331(x9331, x7156, x3387);
  nand n9332(x9332, x9331, x9330);
  nand n9333(x9333, x2272, x9323);
  nand n9334(x9334, x7169, x9326);
  nand n9335(x9335, x9334, x9333);
  nand n9336(x9336, x2272, x9329);
  nand n9337(x9337, x7169, x9332);
  nand n9338(x9338, x9337, x9336);
  nand n9339(x9339, x2275, x9335);
  nand n9340(x9340, x7176, x9338);
  nand n9341(x9341, x9340, x9339);
  nand n9342(x9342, x2269, x4301);
  nand n9343(x9343, x7156, x4171);
  nand n9344(x9344, x9343, x9342);
  nand n9345(x9345, x2269, x4041);
  nand n9346(x9346, x7156, x3911);
  nand n9347(x9347, x9346, x9345);
  nand n9348(x9348, x2269, x3781);
  nand n9349(x9349, x7156, x3651);
  nand n9350(x9350, x9349, x9348);
  nand n9351(x9351, x2269, x3521);
  nand n9352(x9352, x7156, x3391);
  nand n9353(x9353, x9352, x9351);
  nand n9354(x9354, x2272, x9344);
  nand n9355(x9355, x7169, x9347);
  nand n9356(x9356, x9355, x9354);
  nand n9357(x9357, x2272, x9350);
  nand n9358(x9358, x7169, x9353);
  nand n9359(x9359, x9358, x9357);
  nand n9360(x9360, x2275, x9356);
  nand n9361(x9361, x7176, x9359);
  nand n9362(x9362, x9361, x9360);
  nand n9363(x9363, x2269, x4305);
  nand n9364(x9364, x7156, x4175);
  nand n9365(x9365, x9364, x9363);
  nand n9366(x9366, x2269, x4045);
  nand n9367(x9367, x7156, x3915);
  nand n9368(x9368, x9367, x9366);
  nand n9369(x9369, x2269, x3785);
  nand n9370(x9370, x7156, x3655);
  nand n9371(x9371, x9370, x9369);
  nand n9372(x9372, x2269, x3525);
  nand n9373(x9373, x7156, x3395);
  nand n9374(x9374, x9373, x9372);
  nand n9375(x9375, x2272, x9365);
  nand n9376(x9376, x7169, x9368);
  nand n9377(x9377, x9376, x9375);
  nand n9378(x9378, x2272, x9371);
  nand n9379(x9379, x7169, x9374);
  nand n9380(x9380, x9379, x9378);
  nand n9381(x9381, x2275, x9377);
  nand n9382(x9382, x7176, x9380);
  nand n9383(x9383, x9382, x9381);
  nand n9384(x9384, x2269, x4309);
  nand n9385(x9385, x7156, x4179);
  nand n9386(x9386, x9385, x9384);
  nand n9387(x9387, x2269, x4049);
  nand n9388(x9388, x7156, x3919);
  nand n9389(x9389, x9388, x9387);
  nand n9390(x9390, x2269, x3789);
  nand n9391(x9391, x7156, x3659);
  nand n9392(x9392, x9391, x9390);
  nand n9393(x9393, x2269, x3529);
  nand n9394(x9394, x7156, x3399);
  nand n9395(x9395, x9394, x9393);
  nand n9396(x9396, x2272, x9386);
  nand n9397(x9397, x7169, x9389);
  nand n9398(x9398, x9397, x9396);
  nand n9399(x9399, x2272, x9392);
  nand n9400(x9400, x7169, x9395);
  nand n9401(x9401, x9400, x9399);
  nand n9402(x9402, x2275, x9398);
  nand n9403(x9403, x7176, x9401);
  nand n9404(x9404, x9403, x9402);
  nand n9405(x9405, x2269, x4313);
  nand n9406(x9406, x7156, x4183);
  nand n9407(x9407, x9406, x9405);
  nand n9408(x9408, x2269, x4053);
  nand n9409(x9409, x7156, x3923);
  nand n9410(x9410, x9409, x9408);
  nand n9411(x9411, x2269, x3793);
  nand n9412(x9412, x7156, x3663);
  nand n9413(x9413, x9412, x9411);
  nand n9414(x9414, x2269, x3533);
  nand n9415(x9415, x7156, x3403);
  nand n9416(x9416, x9415, x9414);
  nand n9417(x9417, x2272, x9407);
  nand n9418(x9418, x7169, x9410);
  nand n9419(x9419, x9418, x9417);
  nand n9420(x9420, x2272, x9413);
  nand n9421(x9421, x7169, x9416);
  nand n9422(x9422, x9421, x9420);
  nand n9423(x9423, x2275, x9419);
  nand n9424(x9424, x7176, x9422);
  nand n9425(x9425, x9424, x9423);
  nand n9426(x9426, x2269, x4317);
  nand n9427(x9427, x7156, x4187);
  nand n9428(x9428, x9427, x9426);
  nand n9429(x9429, x2269, x4057);
  nand n9430(x9430, x7156, x3927);
  nand n9431(x9431, x9430, x9429);
  nand n9432(x9432, x2269, x3797);
  nand n9433(x9433, x7156, x3667);
  nand n9434(x9434, x9433, x9432);
  nand n9435(x9435, x2269, x3537);
  nand n9436(x9436, x7156, x3407);
  nand n9437(x9437, x9436, x9435);
  nand n9438(x9438, x2272, x9428);
  nand n9439(x9439, x7169, x9431);
  nand n9440(x9440, x9439, x9438);
  nand n9441(x9441, x2272, x9434);
  nand n9442(x9442, x7169, x9437);
  nand n9443(x9443, x9442, x9441);
  nand n9444(x9444, x2275, x9440);
  nand n9445(x9445, x7176, x9443);
  nand n9446(x9446, x9445, x9444);
  nand n9447(x9447, x2269, x4321);
  nand n9448(x9448, x7156, x4191);
  nand n9449(x9449, x9448, x9447);
  nand n9450(x9450, x2269, x4061);
  nand n9451(x9451, x7156, x3931);
  nand n9452(x9452, x9451, x9450);
  nand n9453(x9453, x2269, x3801);
  nand n9454(x9454, x7156, x3671);
  nand n9455(x9455, x9454, x9453);
  nand n9456(x9456, x2269, x3541);
  nand n9457(x9457, x7156, x3411);
  nand n9458(x9458, x9457, x9456);
  nand n9459(x9459, x2272, x9449);
  nand n9460(x9460, x7169, x9452);
  nand n9461(x9461, x9460, x9459);
  nand n9462(x9462, x2272, x9455);
  nand n9463(x9463, x7169, x9458);
  nand n9464(x9464, x9463, x9462);
  nand n9465(x9465, x2275, x9461);
  nand n9466(x9466, x7176, x9464);
  nand n9467(x9467, x9466, x9465);
  nand n9468(x9468, x2269, x4325);
  nand n9469(x9469, x7156, x4195);
  nand n9470(x9470, x9469, x9468);
  nand n9471(x9471, x2269, x4065);
  nand n9472(x9472, x7156, x3935);
  nand n9473(x9473, x9472, x9471);
  nand n9474(x9474, x2269, x3805);
  nand n9475(x9475, x7156, x3675);
  nand n9476(x9476, x9475, x9474);
  nand n9477(x9477, x2269, x3545);
  nand n9478(x9478, x7156, x3415);
  nand n9479(x9479, x9478, x9477);
  nand n9480(x9480, x2272, x9470);
  nand n9481(x9481, x7169, x9473);
  nand n9482(x9482, x9481, x9480);
  nand n9483(x9483, x2272, x9476);
  nand n9484(x9484, x7169, x9479);
  nand n9485(x9485, x9484, x9483);
  nand n9486(x9486, x2275, x9482);
  nand n9487(x9487, x7176, x9485);
  nand n9488(x9488, x9487, x9486);
  nand n9489(x9489, x2269, x4329);
  nand n9490(x9490, x7156, x4199);
  nand n9491(x9491, x9490, x9489);
  nand n9492(x9492, x2269, x4069);
  nand n9493(x9493, x7156, x3939);
  nand n9494(x9494, x9493, x9492);
  nand n9495(x9495, x2269, x3809);
  nand n9496(x9496, x7156, x3679);
  nand n9497(x9497, x9496, x9495);
  nand n9498(x9498, x2269, x3549);
  nand n9499(x9499, x7156, x3419);
  nand n9500(x9500, x9499, x9498);
  nand n9501(x9501, x2272, x9491);
  nand n9502(x9502, x7169, x9494);
  nand n9503(x9503, x9502, x9501);
  nand n9504(x9504, x2272, x9497);
  nand n9505(x9505, x7169, x9500);
  nand n9506(x9506, x9505, x9504);
  nand n9507(x9507, x2275, x9503);
  nand n9508(x9508, x7176, x9506);
  nand n9509(x9509, x9508, x9507);
  nand n9510(x9510, x2269, x4333);
  nand n9511(x9511, x7156, x4203);
  nand n9512(x9512, x9511, x9510);
  nand n9513(x9513, x2269, x4073);
  nand n9514(x9514, x7156, x3943);
  nand n9515(x9515, x9514, x9513);
  nand n9516(x9516, x2269, x3813);
  nand n9517(x9517, x7156, x3683);
  nand n9518(x9518, x9517, x9516);
  nand n9519(x9519, x2269, x3553);
  nand n9520(x9520, x7156, x3423);
  nand n9521(x9521, x9520, x9519);
  nand n9522(x9522, x2272, x9512);
  nand n9523(x9523, x7169, x9515);
  nand n9524(x9524, x9523, x9522);
  nand n9525(x9525, x2272, x9518);
  nand n9526(x9526, x7169, x9521);
  nand n9527(x9527, x9526, x9525);
  nand n9528(x9528, x2275, x9524);
  nand n9529(x9529, x7176, x9527);
  nand n9530(x9530, x9529, x9528);
  nand n9531(x9531, x2269, x4337);
  nand n9532(x9532, x7156, x4207);
  nand n9533(x9533, x9532, x9531);
  nand n9534(x9534, x2269, x4077);
  nand n9535(x9535, x7156, x3947);
  nand n9536(x9536, x9535, x9534);
  nand n9537(x9537, x2269, x3817);
  nand n9538(x9538, x7156, x3687);
  nand n9539(x9539, x9538, x9537);
  nand n9540(x9540, x2269, x3557);
  nand n9541(x9541, x7156, x3427);
  nand n9542(x9542, x9541, x9540);
  nand n9543(x9543, x2272, x9533);
  nand n9544(x9544, x7169, x9536);
  nand n9545(x9545, x9544, x9543);
  nand n9546(x9546, x2272, x9539);
  nand n9547(x9547, x7169, x9542);
  nand n9548(x9548, x9547, x9546);
  nand n9549(x9549, x2275, x9545);
  nand n9550(x9550, x7176, x9548);
  nand n9551(x9551, x9550, x9549);
  nand n9552(x9552, x2269, x4341);
  nand n9553(x9553, x7156, x4211);
  nand n9554(x9554, x9553, x9552);
  nand n9555(x9555, x2269, x4081);
  nand n9556(x9556, x7156, x3951);
  nand n9557(x9557, x9556, x9555);
  nand n9558(x9558, x2269, x3821);
  nand n9559(x9559, x7156, x3691);
  nand n9560(x9560, x9559, x9558);
  nand n9561(x9561, x2269, x3561);
  nand n9562(x9562, x7156, x3431);
  nand n9563(x9563, x9562, x9561);
  nand n9564(x9564, x2272, x9554);
  nand n9565(x9565, x7169, x9557);
  nand n9566(x9566, x9565, x9564);
  nand n9567(x9567, x2272, x9560);
  nand n9568(x9568, x7169, x9563);
  nand n9569(x9569, x9568, x9567);
  nand n9570(x9570, x2275, x9566);
  nand n9571(x9571, x7176, x9569);
  nand n9572(x9572, x9571, x9570);
  nand n9573(x9573, x2269, x4345);
  nand n9574(x9574, x7156, x4215);
  nand n9575(x9575, x9574, x9573);
  nand n9576(x9576, x2269, x4085);
  nand n9577(x9577, x7156, x3955);
  nand n9578(x9578, x9577, x9576);
  nand n9579(x9579, x2269, x3825);
  nand n9580(x9580, x7156, x3695);
  nand n9581(x9581, x9580, x9579);
  nand n9582(x9582, x2269, x3565);
  nand n9583(x9583, x7156, x3435);
  nand n9584(x9584, x9583, x9582);
  nand n9585(x9585, x2272, x9575);
  nand n9586(x9586, x7169, x9578);
  nand n9587(x9587, x9586, x9585);
  nand n9588(x9588, x2272, x9581);
  nand n9589(x9589, x7169, x9584);
  nand n9590(x9590, x9589, x9588);
  nand n9591(x9591, x2275, x9587);
  nand n9592(x9592, x7176, x9590);
  nand n9593(x9593, x9592, x9591);
  nand n9594(x9594, x2269, x4349);
  nand n9595(x9595, x7156, x4219);
  nand n9596(x9596, x9595, x9594);
  nand n9597(x9597, x2269, x4089);
  nand n9598(x9598, x7156, x3959);
  nand n9599(x9599, x9598, x9597);
  nand n9600(x9600, x2269, x3829);
  nand n9601(x9601, x7156, x3699);
  nand n9602(x9602, x9601, x9600);
  nand n9603(x9603, x2269, x3569);
  nand n9604(x9604, x7156, x3439);
  nand n9605(x9605, x9604, x9603);
  nand n9606(x9606, x2272, x9596);
  nand n9607(x9607, x7169, x9599);
  nand n9608(x9608, x9607, x9606);
  nand n9609(x9609, x2272, x9602);
  nand n9610(x9610, x7169, x9605);
  nand n9611(x9611, x9610, x9609);
  nand n9612(x9612, x2275, x9608);
  nand n9613(x9613, x7176, x9611);
  nand n9614(x9614, x9613, x9612);
  nand n9615(x9615, x2269, x4353);
  nand n9616(x9616, x7156, x4223);
  nand n9617(x9617, x9616, x9615);
  nand n9618(x9618, x2269, x4093);
  nand n9619(x9619, x7156, x3963);
  nand n9620(x9620, x9619, x9618);
  nand n9621(x9621, x2269, x3833);
  nand n9622(x9622, x7156, x3703);
  nand n9623(x9623, x9622, x9621);
  nand n9624(x9624, x2269, x3573);
  nand n9625(x9625, x7156, x3443);
  nand n9626(x9626, x9625, x9624);
  nand n9627(x9627, x2272, x9617);
  nand n9628(x9628, x7169, x9620);
  nand n9629(x9629, x9628, x9627);
  nand n9630(x9630, x2272, x9623);
  nand n9631(x9631, x7169, x9626);
  nand n9632(x9632, x9631, x9630);
  nand n9633(x9633, x2275, x9629);
  nand n9634(x9634, x7176, x9632);
  nand n9635(x9635, x9634, x9633);
  nand n9636(x9636, x2269, x4357);
  nand n9637(x9637, x7156, x4227);
  nand n9638(x9638, x9637, x9636);
  nand n9639(x9639, x2269, x4097);
  nand n9640(x9640, x7156, x3967);
  nand n9641(x9641, x9640, x9639);
  nand n9642(x9642, x2269, x3837);
  nand n9643(x9643, x7156, x3707);
  nand n9644(x9644, x9643, x9642);
  nand n9645(x9645, x2269, x3577);
  nand n9646(x9646, x7156, x3447);
  nand n9647(x9647, x9646, x9645);
  nand n9648(x9648, x2272, x9638);
  nand n9649(x9649, x7169, x9641);
  nand n9650(x9650, x9649, x9648);
  nand n9651(x9651, x2272, x9644);
  nand n9652(x9652, x7169, x9647);
  nand n9653(x9653, x9652, x9651);
  nand n9654(x9654, x2275, x9650);
  nand n9655(x9655, x7176, x9653);
  nand n9656(x9656, x9655, x9654);
  nand n9657(x9657, x2269, x4361);
  nand n9658(x9658, x7156, x4231);
  nand n9659(x9659, x9658, x9657);
  nand n9660(x9660, x2269, x4101);
  nand n9661(x9661, x7156, x3971);
  nand n9662(x9662, x9661, x9660);
  nand n9663(x9663, x2269, x3841);
  nand n9664(x9664, x7156, x3711);
  nand n9665(x9665, x9664, x9663);
  nand n9666(x9666, x2269, x3581);
  nand n9667(x9667, x7156, x3451);
  nand n9668(x9668, x9667, x9666);
  nand n9669(x9669, x2272, x9659);
  nand n9670(x9670, x7169, x9662);
  nand n9671(x9671, x9670, x9669);
  nand n9672(x9672, x2272, x9665);
  nand n9673(x9673, x7169, x9668);
  nand n9674(x9674, x9673, x9672);
  nand n9675(x9675, x2275, x9671);
  nand n9676(x9676, x7176, x9674);
  nand n9677(x9677, x9676, x9675);
  nand n9678(x9678, x2269, x4365);
  nand n9679(x9679, x7156, x4235);
  nand n9680(x9680, x9679, x9678);
  nand n9681(x9681, x2269, x4105);
  nand n9682(x9682, x7156, x3975);
  nand n9683(x9683, x9682, x9681);
  nand n9684(x9684, x2269, x3845);
  nand n9685(x9685, x7156, x3715);
  nand n9686(x9686, x9685, x9684);
  nand n9687(x9687, x2269, x3585);
  nand n9688(x9688, x7156, x3455);
  nand n9689(x9689, x9688, x9687);
  nand n9690(x9690, x2272, x9680);
  nand n9691(x9691, x7169, x9683);
  nand n9692(x9692, x9691, x9690);
  nand n9693(x9693, x2272, x9686);
  nand n9694(x9694, x7169, x9689);
  nand n9695(x9695, x9694, x9693);
  nand n9696(x9696, x2275, x9692);
  nand n9697(x9697, x7176, x9695);
  nand n9698(x9698, x9697, x9696);
  nand n9699(x9699, x2269, x4369);
  nand n9700(x9700, x7156, x4239);
  nand n9701(x9701, x9700, x9699);
  nand n9702(x9702, x2269, x4109);
  nand n9703(x9703, x7156, x3979);
  nand n9704(x9704, x9703, x9702);
  nand n9705(x9705, x2269, x3849);
  nand n9706(x9706, x7156, x3719);
  nand n9707(x9707, x9706, x9705);
  nand n9708(x9708, x2269, x3589);
  nand n9709(x9709, x7156, x3459);
  nand n9710(x9710, x9709, x9708);
  nand n9711(x9711, x2272, x9701);
  nand n9712(x9712, x7169, x9704);
  nand n9713(x9713, x9712, x9711);
  nand n9714(x9714, x2272, x9707);
  nand n9715(x9715, x7169, x9710);
  nand n9716(x9716, x9715, x9714);
  nand n9717(x9717, x2275, x9713);
  nand n9718(x9718, x7176, x9716);
  nand n9719(x9719, x9718, x9717);
  nand n9720(x9720, x2269, x4373);
  nand n9721(x9721, x7156, x4243);
  nand n9722(x9722, x9721, x9720);
  nand n9723(x9723, x2269, x4113);
  nand n9724(x9724, x7156, x3983);
  nand n9725(x9725, x9724, x9723);
  nand n9726(x9726, x2269, x3853);
  nand n9727(x9727, x7156, x3723);
  nand n9728(x9728, x9727, x9726);
  nand n9729(x9729, x2269, x3593);
  nand n9730(x9730, x7156, x3463);
  nand n9731(x9731, x9730, x9729);
  nand n9732(x9732, x2272, x9722);
  nand n9733(x9733, x7169, x9725);
  nand n9734(x9734, x9733, x9732);
  nand n9735(x9735, x2272, x9728);
  nand n9736(x9736, x7169, x9731);
  nand n9737(x9737, x9736, x9735);
  nand n9738(x9738, x2275, x9734);
  nand n9739(x9739, x7176, x9737);
  nand n9740(x9740, x9739, x9738);
  nand n9741(x9741, x2269, x4377);
  nand n9742(x9742, x7156, x4247);
  nand n9743(x9743, x9742, x9741);
  nand n9744(x9744, x2269, x4117);
  nand n9745(x9745, x7156, x3987);
  nand n9746(x9746, x9745, x9744);
  nand n9747(x9747, x2269, x3857);
  nand n9748(x9748, x7156, x3727);
  nand n9749(x9749, x9748, x9747);
  nand n9750(x9750, x2269, x3597);
  nand n9751(x9751, x7156, x3467);
  nand n9752(x9752, x9751, x9750);
  nand n9753(x9753, x2272, x9743);
  nand n9754(x9754, x7169, x9746);
  nand n9755(x9755, x9754, x9753);
  nand n9756(x9756, x2272, x9749);
  nand n9757(x9757, x7169, x9752);
  nand n9758(x9758, x9757, x9756);
  nand n9759(x9759, x2275, x9755);
  nand n9760(x9760, x7176, x9758);
  nand n9761(x9761, x9760, x9759);
  nand n9762(x9762, x2269, x4381);
  nand n9763(x9763, x7156, x4251);
  nand n9764(x9764, x9763, x9762);
  nand n9765(x9765, x2269, x4121);
  nand n9766(x9766, x7156, x3991);
  nand n9767(x9767, x9766, x9765);
  nand n9768(x9768, x2269, x3861);
  nand n9769(x9769, x7156, x3731);
  nand n9770(x9770, x9769, x9768);
  nand n9771(x9771, x2269, x3601);
  nand n9772(x9772, x7156, x3471);
  nand n9773(x9773, x9772, x9771);
  nand n9774(x9774, x2272, x9764);
  nand n9775(x9775, x7169, x9767);
  nand n9776(x9776, x9775, x9774);
  nand n9777(x9777, x2272, x9770);
  nand n9778(x9778, x7169, x9773);
  nand n9779(x9779, x9778, x9777);
  nand n9780(x9780, x2275, x9776);
  nand n9781(x9781, x7176, x9779);
  nand n9782(x9782, x9781, x9780);
  nand n9783(x9783, x2269, x4385);
  nand n9784(x9784, x7156, x4255);
  nand n9785(x9785, x9784, x9783);
  nand n9786(x9786, x2269, x4125);
  nand n9787(x9787, x7156, x3995);
  nand n9788(x9788, x9787, x9786);
  nand n9789(x9789, x2269, x3865);
  nand n9790(x9790, x7156, x3735);
  nand n9791(x9791, x9790, x9789);
  nand n9792(x9792, x2269, x3605);
  nand n9793(x9793, x7156, x3475);
  nand n9794(x9794, x9793, x9792);
  nand n9795(x9795, x2272, x9785);
  nand n9796(x9796, x7169, x9788);
  nand n9797(x9797, x9796, x9795);
  nand n9798(x9798, x2272, x9791);
  nand n9799(x9799, x7169, x9794);
  nand n9800(x9800, x9799, x9798);
  nand n9801(x9801, x2275, x9797);
  nand n9802(x9802, x7176, x9800);
  nand n9803(x9803, x9802, x9801);
  nand n9804(x9804, x2269, x4389);
  nand n9805(x9805, x7156, x4259);
  nand n9806(x9806, x9805, x9804);
  nand n9807(x9807, x2269, x4129);
  nand n9808(x9808, x7156, x3999);
  nand n9809(x9809, x9808, x9807);
  nand n9810(x9810, x2269, x3869);
  nand n9811(x9811, x7156, x3739);
  nand n9812(x9812, x9811, x9810);
  nand n9813(x9813, x2269, x3609);
  nand n9814(x9814, x7156, x3479);
  nand n9815(x9815, x9814, x9813);
  nand n9816(x9816, x2272, x9806);
  nand n9817(x9817, x7169, x9809);
  nand n9818(x9818, x9817, x9816);
  nand n9819(x9819, x2272, x9812);
  nand n9820(x9820, x7169, x9815);
  nand n9821(x9821, x9820, x9819);
  nand n9822(x9822, x2275, x9818);
  nand n9823(x9823, x7176, x9821);
  nand n9824(x9824, x9823, x9822);
  nand n9825(x9825, x2269, x4393);
  nand n9826(x9826, x7156, x4263);
  nand n9827(x9827, x9826, x9825);
  nand n9828(x9828, x2269, x4133);
  nand n9829(x9829, x7156, x4003);
  nand n9830(x9830, x9829, x9828);
  nand n9831(x9831, x2269, x3873);
  nand n9832(x9832, x7156, x3743);
  nand n9833(x9833, x9832, x9831);
  nand n9834(x9834, x2269, x3613);
  nand n9835(x9835, x7156, x3483);
  nand n9836(x9836, x9835, x9834);
  nand n9837(x9837, x2272, x9827);
  nand n9838(x9838, x7169, x9830);
  nand n9839(x9839, x9838, x9837);
  nand n9840(x9840, x2272, x9833);
  nand n9841(x9841, x7169, x9836);
  nand n9842(x9842, x9841, x9840);
  nand n9843(x9843, x2275, x9839);
  nand n9844(x9844, x7176, x9842);
  nand n9845(x9845, x9844, x9843);
  nand n9846(x9846, x71202, x4269);
  nand n9847(x9847, x1448, x4139);
  nand n9848(x9848, x9847, x9846);
  nand n9849(x9849, x71202, x4009);
  nand n9850(x9850, x1448, x3879);
  nand n9851(x9851, x9850, x9849);
  nand n9852(x9852, x71202, x3749);
  nand n9853(x9853, x1448, x3619);
  nand n9854(x9854, x9853, x9852);
  nand n9855(x9855, x71202, x3489);
  nand n9856(x9856, x1448, x3359);
  nand n9857(x9857, x9856, x9855);
  nand n9858(x9858, x71205, x9848);
  nand n9859(x9859, x1461, x9851);
  nand n9860(x9860, x9859, x9858);
  nand n9861(x9861, x71205, x9854);
  nand n9862(x9862, x1461, x9857);
  nand n9863(x9863, x9862, x9861);
  nand n9864(x9864, x71210, x9860);
  nand n9865(x9865, x1468, x9863);
  nand n9866(x9866, x9865, x9864);
  nand n9867(x9867, x71202, x4273);
  nand n9868(x9868, x1448, x4143);
  nand n9869(x9869, x9868, x9867);
  nand n9870(x9870, x71202, x4013);
  nand n9871(x9871, x1448, x3883);
  nand n9872(x9872, x9871, x9870);
  nand n9873(x9873, x71202, x3753);
  nand n9874(x9874, x1448, x3623);
  nand n9875(x9875, x9874, x9873);
  nand n9876(x9876, x71202, x3493);
  nand n9877(x9877, x1448, x3363);
  nand n9878(x9878, x9877, x9876);
  nand n9879(x9879, x71205, x9869);
  nand n9880(x9880, x1461, x9872);
  nand n9881(x9881, x9880, x9879);
  nand n9882(x9882, x71205, x9875);
  nand n9883(x9883, x1461, x9878);
  nand n9884(x9884, x9883, x9882);
  nand n9885(x9885, x71210, x9881);
  nand n9886(x9886, x1468, x9884);
  nand n9887(x9887, x9886, x9885);
  nand n9888(x9888, x71202, x4277);
  nand n9889(x9889, x1448, x4147);
  nand n9890(x9890, x9889, x9888);
  nand n9891(x9891, x71202, x4017);
  nand n9892(x9892, x1448, x3887);
  nand n9893(x9893, x9892, x9891);
  nand n9894(x9894, x71202, x3757);
  nand n9895(x9895, x1448, x3627);
  nand n9896(x9896, x9895, x9894);
  nand n9897(x9897, x71202, x3497);
  nand n9898(x9898, x1448, x3367);
  nand n9899(x9899, x9898, x9897);
  nand n9900(x9900, x71205, x9890);
  nand n9901(x9901, x1461, x9893);
  nand n9902(x9902, x9901, x9900);
  nand n9903(x9903, x71205, x9896);
  nand n9904(x9904, x1461, x9899);
  nand n9905(x9905, x9904, x9903);
  nand n9906(x9906, x71210, x9902);
  nand n9907(x9907, x1468, x9905);
  nand n9908(x9908, x9907, x9906);
  nand n9909(x9909, x71202, x4281);
  nand n9910(x9910, x1448, x4151);
  nand n9911(x9911, x9910, x9909);
  nand n9912(x9912, x71202, x4021);
  nand n9913(x9913, x1448, x3891);
  nand n9914(x9914, x9913, x9912);
  nand n9915(x9915, x71202, x3761);
  nand n9916(x9916, x1448, x3631);
  nand n9917(x9917, x9916, x9915);
  nand n9918(x9918, x71202, x3501);
  nand n9919(x9919, x1448, x3371);
  nand n9920(x9920, x9919, x9918);
  nand n9921(x9921, x71205, x9911);
  nand n9922(x9922, x1461, x9914);
  nand n9923(x9923, x9922, x9921);
  nand n9924(x9924, x71205, x9917);
  nand n9925(x9925, x1461, x9920);
  nand n9926(x9926, x9925, x9924);
  nand n9927(x9927, x71210, x9923);
  nand n9928(x9928, x1468, x9926);
  nand n9929(x9929, x9928, x9927);
  nand n9930(x9930, x71202, x4285);
  nand n9931(x9931, x1448, x4155);
  nand n9932(x9932, x9931, x9930);
  nand n9933(x9933, x71202, x4025);
  nand n9934(x9934, x1448, x3895);
  nand n9935(x9935, x9934, x9933);
  nand n9936(x9936, x71202, x3765);
  nand n9937(x9937, x1448, x3635);
  nand n9938(x9938, x9937, x9936);
  nand n9939(x9939, x71202, x3505);
  nand n9940(x9940, x1448, x3375);
  nand n9941(x9941, x9940, x9939);
  nand n9942(x9942, x71205, x9932);
  nand n9943(x9943, x1461, x9935);
  nand n9944(x9944, x9943, x9942);
  nand n9945(x9945, x71205, x9938);
  nand n9946(x9946, x1461, x9941);
  nand n9947(x9947, x9946, x9945);
  nand n9948(x9948, x71210, x9944);
  nand n9949(x9949, x1468, x9947);
  nand n9950(x9950, x9949, x9948);
  nand n9951(x9951, x71202, x4289);
  nand n9952(x9952, x1448, x4159);
  nand n9953(x9953, x9952, x9951);
  nand n9954(x9954, x71202, x4029);
  nand n9955(x9955, x1448, x3899);
  nand n9956(x9956, x9955, x9954);
  nand n9957(x9957, x71202, x3769);
  nand n9958(x9958, x1448, x3639);
  nand n9959(x9959, x9958, x9957);
  nand n9960(x9960, x71202, x3509);
  nand n9961(x9961, x1448, x3379);
  nand n9962(x9962, x9961, x9960);
  nand n9963(x9963, x71205, x9953);
  nand n9964(x9964, x1461, x9956);
  nand n9965(x9965, x9964, x9963);
  nand n9966(x9966, x71205, x9959);
  nand n9967(x9967, x1461, x9962);
  nand n9968(x9968, x9967, x9966);
  nand n9969(x9969, x71210, x9965);
  nand n9970(x9970, x1468, x9968);
  nand n9971(x9971, x9970, x9969);
  nand n9972(x9972, x71202, x4293);
  nand n9973(x9973, x1448, x4163);
  nand n9974(x9974, x9973, x9972);
  nand n9975(x9975, x71202, x4033);
  nand n9976(x9976, x1448, x3903);
  nand n9977(x9977, x9976, x9975);
  nand n9978(x9978, x71202, x3773);
  nand n9979(x9979, x1448, x3643);
  nand n9980(x9980, x9979, x9978);
  nand n9981(x9981, x71202, x3513);
  nand n9982(x9982, x1448, x3383);
  nand n9983(x9983, x9982, x9981);
  nand n9984(x9984, x71205, x9974);
  nand n9985(x9985, x1461, x9977);
  nand n9986(x9986, x9985, x9984);
  nand n9987(x9987, x71205, x9980);
  nand n9988(x9988, x1461, x9983);
  nand n9989(x9989, x9988, x9987);
  nand n9990(x9990, x71210, x9986);
  nand n9991(x9991, x1468, x9989);
  nand n9992(x9992, x9991, x9990);
  nand n9993(x9993, x71202, x4297);
  nand n9994(x9994, x1448, x4167);
  nand n9995(x9995, x9994, x9993);
  nand n9996(x9996, x71202, x4037);
  nand n9997(x9997, x1448, x3907);
  nand n9998(x9998, x9997, x9996);
  nand n9999(x9999, x71202, x3777);
  nand n10000(x10000, x1448, x3647);
  nand n10001(x10001, x10000, x9999);
  nand n10002(x10002, x71202, x3517);
  nand n10003(x10003, x1448, x3387);
  nand n10004(x10004, x10003, x10002);
  nand n10005(x10005, x71205, x9995);
  nand n10006(x10006, x1461, x9998);
  nand n10007(x10007, x10006, x10005);
  nand n10008(x10008, x71205, x10001);
  nand n10009(x10009, x1461, x10004);
  nand n10010(x10010, x10009, x10008);
  nand n10011(x10011, x71210, x10007);
  nand n10012(x10012, x1468, x10010);
  nand n10013(x10013, x10012, x10011);
  nand n10014(x10014, x71202, x4301);
  nand n10015(x10015, x1448, x4171);
  nand n10016(x10016, x10015, x10014);
  nand n10017(x10017, x71202, x4041);
  nand n10018(x10018, x1448, x3911);
  nand n10019(x10019, x10018, x10017);
  nand n10020(x10020, x71202, x3781);
  nand n10021(x10021, x1448, x3651);
  nand n10022(x10022, x10021, x10020);
  nand n10023(x10023, x71202, x3521);
  nand n10024(x10024, x1448, x3391);
  nand n10025(x10025, x10024, x10023);
  nand n10026(x10026, x71205, x10016);
  nand n10027(x10027, x1461, x10019);
  nand n10028(x10028, x10027, x10026);
  nand n10029(x10029, x71205, x10022);
  nand n10030(x10030, x1461, x10025);
  nand n10031(x10031, x10030, x10029);
  nand n10032(x10032, x71210, x10028);
  nand n10033(x10033, x1468, x10031);
  nand n10034(x10034, x10033, x10032);
  nand n10035(x10035, x71202, x4305);
  nand n10036(x10036, x1448, x4175);
  nand n10037(x10037, x10036, x10035);
  nand n10038(x10038, x71202, x4045);
  nand n10039(x10039, x1448, x3915);
  nand n10040(x10040, x10039, x10038);
  nand n10041(x10041, x71202, x3785);
  nand n10042(x10042, x1448, x3655);
  nand n10043(x10043, x10042, x10041);
  nand n10044(x10044, x71202, x3525);
  nand n10045(x10045, x1448, x3395);
  nand n10046(x10046, x10045, x10044);
  nand n10047(x10047, x71205, x10037);
  nand n10048(x10048, x1461, x10040);
  nand n10049(x10049, x10048, x10047);
  nand n10050(x10050, x71205, x10043);
  nand n10051(x10051, x1461, x10046);
  nand n10052(x10052, x10051, x10050);
  nand n10053(x10053, x71210, x10049);
  nand n10054(x10054, x1468, x10052);
  nand n10055(x10055, x10054, x10053);
  nand n10056(x10056, x71202, x4309);
  nand n10057(x10057, x1448, x4179);
  nand n10058(x10058, x10057, x10056);
  nand n10059(x10059, x71202, x4049);
  nand n10060(x10060, x1448, x3919);
  nand n10061(x10061, x10060, x10059);
  nand n10062(x10062, x71202, x3789);
  nand n10063(x10063, x1448, x3659);
  nand n10064(x10064, x10063, x10062);
  nand n10065(x10065, x71202, x3529);
  nand n10066(x10066, x1448, x3399);
  nand n10067(x10067, x10066, x10065);
  nand n10068(x10068, x71205, x10058);
  nand n10069(x10069, x1461, x10061);
  nand n10070(x10070, x10069, x10068);
  nand n10071(x10071, x71205, x10064);
  nand n10072(x10072, x1461, x10067);
  nand n10073(x10073, x10072, x10071);
  nand n10074(x10074, x71210, x10070);
  nand n10075(x10075, x1468, x10073);
  nand n10076(x10076, x10075, x10074);
  nand n10077(x10077, x71202, x4313);
  nand n10078(x10078, x1448, x4183);
  nand n10079(x10079, x10078, x10077);
  nand n10080(x10080, x71202, x4053);
  nand n10081(x10081, x1448, x3923);
  nand n10082(x10082, x10081, x10080);
  nand n10083(x10083, x71202, x3793);
  nand n10084(x10084, x1448, x3663);
  nand n10085(x10085, x10084, x10083);
  nand n10086(x10086, x71202, x3533);
  nand n10087(x10087, x1448, x3403);
  nand n10088(x10088, x10087, x10086);
  nand n10089(x10089, x71205, x10079);
  nand n10090(x10090, x1461, x10082);
  nand n10091(x10091, x10090, x10089);
  nand n10092(x10092, x71205, x10085);
  nand n10093(x10093, x1461, x10088);
  nand n10094(x10094, x10093, x10092);
  nand n10095(x10095, x71210, x10091);
  nand n10096(x10096, x1468, x10094);
  nand n10097(x10097, x10096, x10095);
  nand n10098(x10098, x71202, x4317);
  nand n10099(x10099, x1448, x4187);
  nand n10100(x10100, x10099, x10098);
  nand n10101(x10101, x71202, x4057);
  nand n10102(x10102, x1448, x3927);
  nand n10103(x10103, x10102, x10101);
  nand n10104(x10104, x71202, x3797);
  nand n10105(x10105, x1448, x3667);
  nand n10106(x10106, x10105, x10104);
  nand n10107(x10107, x71202, x3537);
  nand n10108(x10108, x1448, x3407);
  nand n10109(x10109, x10108, x10107);
  nand n10110(x10110, x71205, x10100);
  nand n10111(x10111, x1461, x10103);
  nand n10112(x10112, x10111, x10110);
  nand n10113(x10113, x71205, x10106);
  nand n10114(x10114, x1461, x10109);
  nand n10115(x10115, x10114, x10113);
  nand n10116(x10116, x71210, x10112);
  nand n10117(x10117, x1468, x10115);
  nand n10118(x10118, x10117, x10116);
  nand n10119(x10119, x71202, x4321);
  nand n10120(x10120, x1448, x4191);
  nand n10121(x10121, x10120, x10119);
  nand n10122(x10122, x71202, x4061);
  nand n10123(x10123, x1448, x3931);
  nand n10124(x10124, x10123, x10122);
  nand n10125(x10125, x71202, x3801);
  nand n10126(x10126, x1448, x3671);
  nand n10127(x10127, x10126, x10125);
  nand n10128(x10128, x71202, x3541);
  nand n10129(x10129, x1448, x3411);
  nand n10130(x10130, x10129, x10128);
  nand n10131(x10131, x71205, x10121);
  nand n10132(x10132, x1461, x10124);
  nand n10133(x10133, x10132, x10131);
  nand n10134(x10134, x71205, x10127);
  nand n10135(x10135, x1461, x10130);
  nand n10136(x10136, x10135, x10134);
  nand n10137(x10137, x71210, x10133);
  nand n10138(x10138, x1468, x10136);
  nand n10139(x10139, x10138, x10137);
  nand n10140(x10140, x71202, x4325);
  nand n10141(x10141, x1448, x4195);
  nand n10142(x10142, x10141, x10140);
  nand n10143(x10143, x71202, x4065);
  nand n10144(x10144, x1448, x3935);
  nand n10145(x10145, x10144, x10143);
  nand n10146(x10146, x71202, x3805);
  nand n10147(x10147, x1448, x3675);
  nand n10148(x10148, x10147, x10146);
  nand n10149(x10149, x71202, x3545);
  nand n10150(x10150, x1448, x3415);
  nand n10151(x10151, x10150, x10149);
  nand n10152(x10152, x71205, x10142);
  nand n10153(x10153, x1461, x10145);
  nand n10154(x10154, x10153, x10152);
  nand n10155(x10155, x71205, x10148);
  nand n10156(x10156, x1461, x10151);
  nand n10157(x10157, x10156, x10155);
  nand n10158(x10158, x71210, x10154);
  nand n10159(x10159, x1468, x10157);
  nand n10160(x10160, x10159, x10158);
  nand n10161(x10161, x71202, x4329);
  nand n10162(x10162, x1448, x4199);
  nand n10163(x10163, x10162, x10161);
  nand n10164(x10164, x71202, x4069);
  nand n10165(x10165, x1448, x3939);
  nand n10166(x10166, x10165, x10164);
  nand n10167(x10167, x71202, x3809);
  nand n10168(x10168, x1448, x3679);
  nand n10169(x10169, x10168, x10167);
  nand n10170(x10170, x71202, x3549);
  nand n10171(x10171, x1448, x3419);
  nand n10172(x10172, x10171, x10170);
  nand n10173(x10173, x71205, x10163);
  nand n10174(x10174, x1461, x10166);
  nand n10175(x10175, x10174, x10173);
  nand n10176(x10176, x71205, x10169);
  nand n10177(x10177, x1461, x10172);
  nand n10178(x10178, x10177, x10176);
  nand n10179(x10179, x71210, x10175);
  nand n10180(x10180, x1468, x10178);
  nand n10181(x10181, x10180, x10179);
  nand n10182(x10182, x71202, x4333);
  nand n10183(x10183, x1448, x4203);
  nand n10184(x10184, x10183, x10182);
  nand n10185(x10185, x71202, x4073);
  nand n10186(x10186, x1448, x3943);
  nand n10187(x10187, x10186, x10185);
  nand n10188(x10188, x71202, x3813);
  nand n10189(x10189, x1448, x3683);
  nand n10190(x10190, x10189, x10188);
  nand n10191(x10191, x71202, x3553);
  nand n10192(x10192, x1448, x3423);
  nand n10193(x10193, x10192, x10191);
  nand n10194(x10194, x71205, x10184);
  nand n10195(x10195, x1461, x10187);
  nand n10196(x10196, x10195, x10194);
  nand n10197(x10197, x71205, x10190);
  nand n10198(x10198, x1461, x10193);
  nand n10199(x10199, x10198, x10197);
  nand n10200(x10200, x71210, x10196);
  nand n10201(x10201, x1468, x10199);
  nand n10202(x10202, x10201, x10200);
  nand n10203(x10203, x71202, x4337);
  nand n10204(x10204, x1448, x4207);
  nand n10205(x10205, x10204, x10203);
  nand n10206(x10206, x71202, x4077);
  nand n10207(x10207, x1448, x3947);
  nand n10208(x10208, x10207, x10206);
  nand n10209(x10209, x71202, x3817);
  nand n10210(x10210, x1448, x3687);
  nand n10211(x10211, x10210, x10209);
  nand n10212(x10212, x71202, x3557);
  nand n10213(x10213, x1448, x3427);
  nand n10214(x10214, x10213, x10212);
  nand n10215(x10215, x71205, x10205);
  nand n10216(x10216, x1461, x10208);
  nand n10217(x10217, x10216, x10215);
  nand n10218(x10218, x71205, x10211);
  nand n10219(x10219, x1461, x10214);
  nand n10220(x10220, x10219, x10218);
  nand n10221(x10221, x71210, x10217);
  nand n10222(x10222, x1468, x10220);
  nand n10223(x10223, x10222, x10221);
  nand n10224(x10224, x71202, x4341);
  nand n10225(x10225, x1448, x4211);
  nand n10226(x10226, x10225, x10224);
  nand n10227(x10227, x71202, x4081);
  nand n10228(x10228, x1448, x3951);
  nand n10229(x10229, x10228, x10227);
  nand n10230(x10230, x71202, x3821);
  nand n10231(x10231, x1448, x3691);
  nand n10232(x10232, x10231, x10230);
  nand n10233(x10233, x71202, x3561);
  nand n10234(x10234, x1448, x3431);
  nand n10235(x10235, x10234, x10233);
  nand n10236(x10236, x71205, x10226);
  nand n10237(x10237, x1461, x10229);
  nand n10238(x10238, x10237, x10236);
  nand n10239(x10239, x71205, x10232);
  nand n10240(x10240, x1461, x10235);
  nand n10241(x10241, x10240, x10239);
  nand n10242(x10242, x71210, x10238);
  nand n10243(x10243, x1468, x10241);
  nand n10244(x10244, x10243, x10242);
  nand n10245(x10245, x71202, x4345);
  nand n10246(x10246, x1448, x4215);
  nand n10247(x10247, x10246, x10245);
  nand n10248(x10248, x71202, x4085);
  nand n10249(x10249, x1448, x3955);
  nand n10250(x10250, x10249, x10248);
  nand n10251(x10251, x71202, x3825);
  nand n10252(x10252, x1448, x3695);
  nand n10253(x10253, x10252, x10251);
  nand n10254(x10254, x71202, x3565);
  nand n10255(x10255, x1448, x3435);
  nand n10256(x10256, x10255, x10254);
  nand n10257(x10257, x71205, x10247);
  nand n10258(x10258, x1461, x10250);
  nand n10259(x10259, x10258, x10257);
  nand n10260(x10260, x71205, x10253);
  nand n10261(x10261, x1461, x10256);
  nand n10262(x10262, x10261, x10260);
  nand n10263(x10263, x71210, x10259);
  nand n10264(x10264, x1468, x10262);
  nand n10265(x10265, x10264, x10263);
  nand n10266(x10266, x71202, x4349);
  nand n10267(x10267, x1448, x4219);
  nand n10268(x10268, x10267, x10266);
  nand n10269(x10269, x71202, x4089);
  nand n10270(x10270, x1448, x3959);
  nand n10271(x10271, x10270, x10269);
  nand n10272(x10272, x71202, x3829);
  nand n10273(x10273, x1448, x3699);
  nand n10274(x10274, x10273, x10272);
  nand n10275(x10275, x71202, x3569);
  nand n10276(x10276, x1448, x3439);
  nand n10277(x10277, x10276, x10275);
  nand n10278(x10278, x71205, x10268);
  nand n10279(x10279, x1461, x10271);
  nand n10280(x10280, x10279, x10278);
  nand n10281(x10281, x71205, x10274);
  nand n10282(x10282, x1461, x10277);
  nand n10283(x10283, x10282, x10281);
  nand n10284(x10284, x71210, x10280);
  nand n10285(x10285, x1468, x10283);
  nand n10286(x10286, x10285, x10284);
  nand n10287(x10287, x71202, x4353);
  nand n10288(x10288, x1448, x4223);
  nand n10289(x10289, x10288, x10287);
  nand n10290(x10290, x71202, x4093);
  nand n10291(x10291, x1448, x3963);
  nand n10292(x10292, x10291, x10290);
  nand n10293(x10293, x71202, x3833);
  nand n10294(x10294, x1448, x3703);
  nand n10295(x10295, x10294, x10293);
  nand n10296(x10296, x71202, x3573);
  nand n10297(x10297, x1448, x3443);
  nand n10298(x10298, x10297, x10296);
  nand n10299(x10299, x71205, x10289);
  nand n10300(x10300, x1461, x10292);
  nand n10301(x10301, x10300, x10299);
  nand n10302(x10302, x71205, x10295);
  nand n10303(x10303, x1461, x10298);
  nand n10304(x10304, x10303, x10302);
  nand n10305(x10305, x71210, x10301);
  nand n10306(x10306, x1468, x10304);
  nand n10307(x10307, x10306, x10305);
  nand n10308(x10308, x71202, x4357);
  nand n10309(x10309, x1448, x4227);
  nand n10310(x10310, x10309, x10308);
  nand n10311(x10311, x71202, x4097);
  nand n10312(x10312, x1448, x3967);
  nand n10313(x10313, x10312, x10311);
  nand n10314(x10314, x71202, x3837);
  nand n10315(x10315, x1448, x3707);
  nand n10316(x10316, x10315, x10314);
  nand n10317(x10317, x71202, x3577);
  nand n10318(x10318, x1448, x3447);
  nand n10319(x10319, x10318, x10317);
  nand n10320(x10320, x71205, x10310);
  nand n10321(x10321, x1461, x10313);
  nand n10322(x10322, x10321, x10320);
  nand n10323(x10323, x71205, x10316);
  nand n10324(x10324, x1461, x10319);
  nand n10325(x10325, x10324, x10323);
  nand n10326(x10326, x71210, x10322);
  nand n10327(x10327, x1468, x10325);
  nand n10328(x10328, x10327, x10326);
  nand n10329(x10329, x71202, x4361);
  nand n10330(x10330, x1448, x4231);
  nand n10331(x10331, x10330, x10329);
  nand n10332(x10332, x71202, x4101);
  nand n10333(x10333, x1448, x3971);
  nand n10334(x10334, x10333, x10332);
  nand n10335(x10335, x71202, x3841);
  nand n10336(x10336, x1448, x3711);
  nand n10337(x10337, x10336, x10335);
  nand n10338(x10338, x71202, x3581);
  nand n10339(x10339, x1448, x3451);
  nand n10340(x10340, x10339, x10338);
  nand n10341(x10341, x71205, x10331);
  nand n10342(x10342, x1461, x10334);
  nand n10343(x10343, x10342, x10341);
  nand n10344(x10344, x71205, x10337);
  nand n10345(x10345, x1461, x10340);
  nand n10346(x10346, x10345, x10344);
  nand n10347(x10347, x71210, x10343);
  nand n10348(x10348, x1468, x10346);
  nand n10349(x10349, x10348, x10347);
  nand n10350(x10350, x71202, x4365);
  nand n10351(x10351, x1448, x4235);
  nand n10352(x10352, x10351, x10350);
  nand n10353(x10353, x71202, x4105);
  nand n10354(x10354, x1448, x3975);
  nand n10355(x10355, x10354, x10353);
  nand n10356(x10356, x71202, x3845);
  nand n10357(x10357, x1448, x3715);
  nand n10358(x10358, x10357, x10356);
  nand n10359(x10359, x71202, x3585);
  nand n10360(x10360, x1448, x3455);
  nand n10361(x10361, x10360, x10359);
  nand n10362(x10362, x71205, x10352);
  nand n10363(x10363, x1461, x10355);
  nand n10364(x10364, x10363, x10362);
  nand n10365(x10365, x71205, x10358);
  nand n10366(x10366, x1461, x10361);
  nand n10367(x10367, x10366, x10365);
  nand n10368(x10368, x71210, x10364);
  nand n10369(x10369, x1468, x10367);
  nand n10370(x10370, x10369, x10368);
  nand n10371(x10371, x71202, x4369);
  nand n10372(x10372, x1448, x4239);
  nand n10373(x10373, x10372, x10371);
  nand n10374(x10374, x71202, x4109);
  nand n10375(x10375, x1448, x3979);
  nand n10376(x10376, x10375, x10374);
  nand n10377(x10377, x71202, x3849);
  nand n10378(x10378, x1448, x3719);
  nand n10379(x10379, x10378, x10377);
  nand n10380(x10380, x71202, x3589);
  nand n10381(x10381, x1448, x3459);
  nand n10382(x10382, x10381, x10380);
  nand n10383(x10383, x71205, x10373);
  nand n10384(x10384, x1461, x10376);
  nand n10385(x10385, x10384, x10383);
  nand n10386(x10386, x71205, x10379);
  nand n10387(x10387, x1461, x10382);
  nand n10388(x10388, x10387, x10386);
  nand n10389(x10389, x71210, x10385);
  nand n10390(x10390, x1468, x10388);
  nand n10391(x10391, x10390, x10389);
  nand n10392(x10392, x71202, x4373);
  nand n10393(x10393, x1448, x4243);
  nand n10394(x10394, x10393, x10392);
  nand n10395(x10395, x71202, x4113);
  nand n10396(x10396, x1448, x3983);
  nand n10397(x10397, x10396, x10395);
  nand n10398(x10398, x71202, x3853);
  nand n10399(x10399, x1448, x3723);
  nand n10400(x10400, x10399, x10398);
  nand n10401(x10401, x71202, x3593);
  nand n10402(x10402, x1448, x3463);
  nand n10403(x10403, x10402, x10401);
  nand n10404(x10404, x71205, x10394);
  nand n10405(x10405, x1461, x10397);
  nand n10406(x10406, x10405, x10404);
  nand n10407(x10407, x71205, x10400);
  nand n10408(x10408, x1461, x10403);
  nand n10409(x10409, x10408, x10407);
  nand n10410(x10410, x71210, x10406);
  nand n10411(x10411, x1468, x10409);
  nand n10412(x10412, x10411, x10410);
  nand n10413(x10413, x71202, x4377);
  nand n10414(x10414, x1448, x4247);
  nand n10415(x10415, x10414, x10413);
  nand n10416(x10416, x71202, x4117);
  nand n10417(x10417, x1448, x3987);
  nand n10418(x10418, x10417, x10416);
  nand n10419(x10419, x71202, x3857);
  nand n10420(x10420, x1448, x3727);
  nand n10421(x10421, x10420, x10419);
  nand n10422(x10422, x71202, x3597);
  nand n10423(x10423, x1448, x3467);
  nand n10424(x10424, x10423, x10422);
  nand n10425(x10425, x71205, x10415);
  nand n10426(x10426, x1461, x10418);
  nand n10427(x10427, x10426, x10425);
  nand n10428(x10428, x71205, x10421);
  nand n10429(x10429, x1461, x10424);
  nand n10430(x10430, x10429, x10428);
  nand n10431(x10431, x71210, x10427);
  nand n10432(x10432, x1468, x10430);
  nand n10433(x10433, x10432, x10431);
  nand n10434(x10434, x71202, x4381);
  nand n10435(x10435, x1448, x4251);
  nand n10436(x10436, x10435, x10434);
  nand n10437(x10437, x71202, x4121);
  nand n10438(x10438, x1448, x3991);
  nand n10439(x10439, x10438, x10437);
  nand n10440(x10440, x71202, x3861);
  nand n10441(x10441, x1448, x3731);
  nand n10442(x10442, x10441, x10440);
  nand n10443(x10443, x71202, x3601);
  nand n10444(x10444, x1448, x3471);
  nand n10445(x10445, x10444, x10443);
  nand n10446(x10446, x71205, x10436);
  nand n10447(x10447, x1461, x10439);
  nand n10448(x10448, x10447, x10446);
  nand n10449(x10449, x71205, x10442);
  nand n10450(x10450, x1461, x10445);
  nand n10451(x10451, x10450, x10449);
  nand n10452(x10452, x71210, x10448);
  nand n10453(x10453, x1468, x10451);
  nand n10454(x10454, x10453, x10452);
  nand n10455(x10455, x71202, x4385);
  nand n10456(x10456, x1448, x4255);
  nand n10457(x10457, x10456, x10455);
  nand n10458(x10458, x71202, x4125);
  nand n10459(x10459, x1448, x3995);
  nand n10460(x10460, x10459, x10458);
  nand n10461(x10461, x71202, x3865);
  nand n10462(x10462, x1448, x3735);
  nand n10463(x10463, x10462, x10461);
  nand n10464(x10464, x71202, x3605);
  nand n10465(x10465, x1448, x3475);
  nand n10466(x10466, x10465, x10464);
  nand n10467(x10467, x71205, x10457);
  nand n10468(x10468, x1461, x10460);
  nand n10469(x10469, x10468, x10467);
  nand n10470(x10470, x71205, x10463);
  nand n10471(x10471, x1461, x10466);
  nand n10472(x10472, x10471, x10470);
  nand n10473(x10473, x71210, x10469);
  nand n10474(x10474, x1468, x10472);
  nand n10475(x10475, x10474, x10473);
  nand n10476(x10476, x71202, x4389);
  nand n10477(x10477, x1448, x4259);
  nand n10478(x10478, x10477, x10476);
  nand n10479(x10479, x71202, x4129);
  nand n10480(x10480, x1448, x3999);
  nand n10481(x10481, x10480, x10479);
  nand n10482(x10482, x71202, x3869);
  nand n10483(x10483, x1448, x3739);
  nand n10484(x10484, x10483, x10482);
  nand n10485(x10485, x71202, x3609);
  nand n10486(x10486, x1448, x3479);
  nand n10487(x10487, x10486, x10485);
  nand n10488(x10488, x71205, x10478);
  nand n10489(x10489, x1461, x10481);
  nand n10490(x10490, x10489, x10488);
  nand n10491(x10491, x71205, x10484);
  nand n10492(x10492, x1461, x10487);
  nand n10493(x10493, x10492, x10491);
  nand n10494(x10494, x71210, x10490);
  nand n10495(x10495, x1468, x10493);
  nand n10496(x10496, x10495, x10494);
  nand n10497(x10497, x71202, x4393);
  nand n10498(x10498, x1448, x4263);
  nand n10499(x10499, x10498, x10497);
  nand n10500(x10500, x71202, x4133);
  nand n10501(x10501, x1448, x4003);
  nand n10502(x10502, x10501, x10500);
  nand n10503(x10503, x71202, x3873);
  nand n10504(x10504, x1448, x3743);
  nand n10505(x10505, x10504, x10503);
  nand n10506(x10506, x71202, x3613);
  nand n10507(x10507, x1448, x3483);
  nand n10508(x10508, x10507, x10506);
  nand n10509(x10509, x71205, x10499);
  nand n10510(x10510, x1461, x10502);
  nand n10511(x10511, x10510, x10509);
  nand n10512(x10512, x71205, x10505);
  nand n10513(x10513, x1461, x10508);
  nand n10514(x10514, x10513, x10512);
  nand n10515(x10515, x71210, x10511);
  nand n10516(x10516, x1468, x10514);
  nand n10517(x10517, x10516, x10515);
  nand n10518(x10518, x2258, x5311);
  nand n10519(x10519, x6481, x5181);
  nand n10520(x10520, x10519, x10518);
  nand n10521(x10521, x2258, x5051);
  nand n10522(x10522, x6481, x4921);
  nand n10523(x10523, x10522, x10521);
  nand n10524(x10524, x2258, x4791);
  nand n10525(x10525, x6481, x4661);
  nand n10526(x10526, x10525, x10524);
  nand n10527(x10527, x2258, x4531);
  nand n10528(x10528, x6481, x4399);
  nand n10529(x10529, x10528, x10527);
  nand n10530(x10530, x2261, x10520);
  nand n10531(x10531, x6494, x10523);
  nand n10532(x10532, x10531, x10530);
  nand n10533(x10533, x2261, x10526);
  nand n10534(x10534, x6494, x10529);
  nand n10535(x10535, x10534, x10533);
  nand n10536(x10536, x2264, x10532);
  nand n10537(x10537, x6501, x10535);
  nand n10538(x10538, x10537, x10536);
  nand n10539(x10539, x2258, x5315);
  nand n10540(x10540, x6481, x5185);
  nand n10541(x10541, x10540, x10539);
  nand n10542(x10542, x2258, x5055);
  nand n10543(x10543, x6481, x4925);
  nand n10544(x10544, x10543, x10542);
  nand n10545(x10545, x2258, x4795);
  nand n10546(x10546, x6481, x4665);
  nand n10547(x10547, x10546, x10545);
  nand n10548(x10548, x2258, x4535);
  nand n10549(x10549, x6481, x4405);
  nand n10550(x10550, x10549, x10548);
  nand n10551(x10551, x2261, x10541);
  nand n10552(x10552, x6494, x10544);
  nand n10553(x10553, x10552, x10551);
  nand n10554(x10554, x2261, x10547);
  nand n10555(x10555, x6494, x10550);
  nand n10556(x10556, x10555, x10554);
  nand n10557(x10557, x2264, x10553);
  nand n10558(x10558, x6501, x10556);
  nand n10559(x10559, x10558, x10557);
  nand n10560(x10560, x2258, x5319);
  nand n10561(x10561, x6481, x5189);
  nand n10562(x10562, x10561, x10560);
  nand n10563(x10563, x2258, x5059);
  nand n10564(x10564, x6481, x4929);
  nand n10565(x10565, x10564, x10563);
  nand n10566(x10566, x2258, x4799);
  nand n10567(x10567, x6481, x4669);
  nand n10568(x10568, x10567, x10566);
  nand n10569(x10569, x2258, x4539);
  nand n10570(x10570, x6481, x4409);
  nand n10571(x10571, x10570, x10569);
  nand n10572(x10572, x2261, x10562);
  nand n10573(x10573, x6494, x10565);
  nand n10574(x10574, x10573, x10572);
  nand n10575(x10575, x2261, x10568);
  nand n10576(x10576, x6494, x10571);
  nand n10577(x10577, x10576, x10575);
  nand n10578(x10578, x2264, x10574);
  nand n10579(x10579, x6501, x10577);
  nand n10580(x10580, x10579, x10578);
  nand n10581(x10581, x2258, x5323);
  nand n10582(x10582, x6481, x5193);
  nand n10583(x10583, x10582, x10581);
  nand n10584(x10584, x2258, x5063);
  nand n10585(x10585, x6481, x4933);
  nand n10586(x10586, x10585, x10584);
  nand n10587(x10587, x2258, x4803);
  nand n10588(x10588, x6481, x4673);
  nand n10589(x10589, x10588, x10587);
  nand n10590(x10590, x2258, x4543);
  nand n10591(x10591, x6481, x4413);
  nand n10592(x10592, x10591, x10590);
  nand n10593(x10593, x2261, x10583);
  nand n10594(x10594, x6494, x10586);
  nand n10595(x10595, x10594, x10593);
  nand n10596(x10596, x2261, x10589);
  nand n10597(x10597, x6494, x10592);
  nand n10598(x10598, x10597, x10596);
  nand n10599(x10599, x2264, x10595);
  nand n10600(x10600, x6501, x10598);
  nand n10601(x10601, x10600, x10599);
  nand n10602(x10602, x2258, x5327);
  nand n10603(x10603, x6481, x5197);
  nand n10604(x10604, x10603, x10602);
  nand n10605(x10605, x2258, x5067);
  nand n10606(x10606, x6481, x4937);
  nand n10607(x10607, x10606, x10605);
  nand n10608(x10608, x2258, x4807);
  nand n10609(x10609, x6481, x4677);
  nand n10610(x10610, x10609, x10608);
  nand n10611(x10611, x2258, x4547);
  nand n10612(x10612, x6481, x4417);
  nand n10613(x10613, x10612, x10611);
  nand n10614(x10614, x2261, x10604);
  nand n10615(x10615, x6494, x10607);
  nand n10616(x10616, x10615, x10614);
  nand n10617(x10617, x2261, x10610);
  nand n10618(x10618, x6494, x10613);
  nand n10619(x10619, x10618, x10617);
  nand n10620(x10620, x2264, x10616);
  nand n10621(x10621, x6501, x10619);
  nand n10622(x10622, x10621, x10620);
  nand n10623(x10623, x2258, x5331);
  nand n10624(x10624, x6481, x5201);
  nand n10625(x10625, x10624, x10623);
  nand n10626(x10626, x2258, x5071);
  nand n10627(x10627, x6481, x4941);
  nand n10628(x10628, x10627, x10626);
  nand n10629(x10629, x2258, x4811);
  nand n10630(x10630, x6481, x4681);
  nand n10631(x10631, x10630, x10629);
  nand n10632(x10632, x2258, x4551);
  nand n10633(x10633, x6481, x4421);
  nand n10634(x10634, x10633, x10632);
  nand n10635(x10635, x2261, x10625);
  nand n10636(x10636, x6494, x10628);
  nand n10637(x10637, x10636, x10635);
  nand n10638(x10638, x2261, x10631);
  nand n10639(x10639, x6494, x10634);
  nand n10640(x10640, x10639, x10638);
  nand n10641(x10641, x2264, x10637);
  nand n10642(x10642, x6501, x10640);
  nand n10643(x10643, x10642, x10641);
  nand n10644(x10644, x2258, x5335);
  nand n10645(x10645, x6481, x5205);
  nand n10646(x10646, x10645, x10644);
  nand n10647(x10647, x2258, x5075);
  nand n10648(x10648, x6481, x4945);
  nand n10649(x10649, x10648, x10647);
  nand n10650(x10650, x2258, x4815);
  nand n10651(x10651, x6481, x4685);
  nand n10652(x10652, x10651, x10650);
  nand n10653(x10653, x2258, x4555);
  nand n10654(x10654, x6481, x4425);
  nand n10655(x10655, x10654, x10653);
  nand n10656(x10656, x2261, x10646);
  nand n10657(x10657, x6494, x10649);
  nand n10658(x10658, x10657, x10656);
  nand n10659(x10659, x2261, x10652);
  nand n10660(x10660, x6494, x10655);
  nand n10661(x10661, x10660, x10659);
  nand n10662(x10662, x2264, x10658);
  nand n10663(x10663, x6501, x10661);
  nand n10664(x10664, x10663, x10662);
  nand n10665(x10665, x2258, x5339);
  nand n10666(x10666, x6481, x5209);
  nand n10667(x10667, x10666, x10665);
  nand n10668(x10668, x2258, x5079);
  nand n10669(x10669, x6481, x4949);
  nand n10670(x10670, x10669, x10668);
  nand n10671(x10671, x2258, x4819);
  nand n10672(x10672, x6481, x4689);
  nand n10673(x10673, x10672, x10671);
  nand n10674(x10674, x2258, x4559);
  nand n10675(x10675, x6481, x4429);
  nand n10676(x10676, x10675, x10674);
  nand n10677(x10677, x2261, x10667);
  nand n10678(x10678, x6494, x10670);
  nand n10679(x10679, x10678, x10677);
  nand n10680(x10680, x2261, x10673);
  nand n10681(x10681, x6494, x10676);
  nand n10682(x10682, x10681, x10680);
  nand n10683(x10683, x2264, x10679);
  nand n10684(x10684, x6501, x10682);
  nand n10685(x10685, x10684, x10683);
  nand n10686(x10686, x2258, x5343);
  nand n10687(x10687, x6481, x5213);
  nand n10688(x10688, x10687, x10686);
  nand n10689(x10689, x2258, x5083);
  nand n10690(x10690, x6481, x4953);
  nand n10691(x10691, x10690, x10689);
  nand n10692(x10692, x2258, x4823);
  nand n10693(x10693, x6481, x4693);
  nand n10694(x10694, x10693, x10692);
  nand n10695(x10695, x2258, x4563);
  nand n10696(x10696, x6481, x4433);
  nand n10697(x10697, x10696, x10695);
  nand n10698(x10698, x2261, x10688);
  nand n10699(x10699, x6494, x10691);
  nand n10700(x10700, x10699, x10698);
  nand n10701(x10701, x2261, x10694);
  nand n10702(x10702, x6494, x10697);
  nand n10703(x10703, x10702, x10701);
  nand n10704(x10704, x2264, x10700);
  nand n10705(x10705, x6501, x10703);
  nand n10706(x10706, x10705, x10704);
  nand n10707(x10707, x2258, x5347);
  nand n10708(x10708, x6481, x5217);
  nand n10709(x10709, x10708, x10707);
  nand n10710(x10710, x2258, x5087);
  nand n10711(x10711, x6481, x4957);
  nand n10712(x10712, x10711, x10710);
  nand n10713(x10713, x2258, x4827);
  nand n10714(x10714, x6481, x4697);
  nand n10715(x10715, x10714, x10713);
  nand n10716(x10716, x2258, x4567);
  nand n10717(x10717, x6481, x4437);
  nand n10718(x10718, x10717, x10716);
  nand n10719(x10719, x2261, x10709);
  nand n10720(x10720, x6494, x10712);
  nand n10721(x10721, x10720, x10719);
  nand n10722(x10722, x2261, x10715);
  nand n10723(x10723, x6494, x10718);
  nand n10724(x10724, x10723, x10722);
  nand n10725(x10725, x2264, x10721);
  nand n10726(x10726, x6501, x10724);
  nand n10727(x10727, x10726, x10725);
  nand n10728(x10728, x2258, x5351);
  nand n10729(x10729, x6481, x5221);
  nand n10730(x10730, x10729, x10728);
  nand n10731(x10731, x2258, x5091);
  nand n10732(x10732, x6481, x4961);
  nand n10733(x10733, x10732, x10731);
  nand n10734(x10734, x2258, x4831);
  nand n10735(x10735, x6481, x4701);
  nand n10736(x10736, x10735, x10734);
  nand n10737(x10737, x2258, x4571);
  nand n10738(x10738, x6481, x4441);
  nand n10739(x10739, x10738, x10737);
  nand n10740(x10740, x2261, x10730);
  nand n10741(x10741, x6494, x10733);
  nand n10742(x10742, x10741, x10740);
  nand n10743(x10743, x2261, x10736);
  nand n10744(x10744, x6494, x10739);
  nand n10745(x10745, x10744, x10743);
  nand n10746(x10746, x2264, x10742);
  nand n10747(x10747, x6501, x10745);
  nand n10748(x10748, x10747, x10746);
  nand n10749(x10749, x2258, x5355);
  nand n10750(x10750, x6481, x5225);
  nand n10751(x10751, x10750, x10749);
  nand n10752(x10752, x2258, x5095);
  nand n10753(x10753, x6481, x4965);
  nand n10754(x10754, x10753, x10752);
  nand n10755(x10755, x2258, x4835);
  nand n10756(x10756, x6481, x4705);
  nand n10757(x10757, x10756, x10755);
  nand n10758(x10758, x2258, x4575);
  nand n10759(x10759, x6481, x4445);
  nand n10760(x10760, x10759, x10758);
  nand n10761(x10761, x2261, x10751);
  nand n10762(x10762, x6494, x10754);
  nand n10763(x10763, x10762, x10761);
  nand n10764(x10764, x2261, x10757);
  nand n10765(x10765, x6494, x10760);
  nand n10766(x10766, x10765, x10764);
  nand n10767(x10767, x2264, x10763);
  nand n10768(x10768, x6501, x10766);
  nand n10769(x10769, x10768, x10767);
  nand n10770(x10770, x2258, x5359);
  nand n10771(x10771, x6481, x5229);
  nand n10772(x10772, x10771, x10770);
  nand n10773(x10773, x2258, x5099);
  nand n10774(x10774, x6481, x4969);
  nand n10775(x10775, x10774, x10773);
  nand n10776(x10776, x2258, x4839);
  nand n10777(x10777, x6481, x4709);
  nand n10778(x10778, x10777, x10776);
  nand n10779(x10779, x2258, x4579);
  nand n10780(x10780, x6481, x4449);
  nand n10781(x10781, x10780, x10779);
  nand n10782(x10782, x2261, x10772);
  nand n10783(x10783, x6494, x10775);
  nand n10784(x10784, x10783, x10782);
  nand n10785(x10785, x2261, x10778);
  nand n10786(x10786, x6494, x10781);
  nand n10787(x10787, x10786, x10785);
  nand n10788(x10788, x2264, x10784);
  nand n10789(x10789, x6501, x10787);
  nand n10790(x10790, x10789, x10788);
  nand n10791(x10791, x2258, x5363);
  nand n10792(x10792, x6481, x5233);
  nand n10793(x10793, x10792, x10791);
  nand n10794(x10794, x2258, x5103);
  nand n10795(x10795, x6481, x4973);
  nand n10796(x10796, x10795, x10794);
  nand n10797(x10797, x2258, x4843);
  nand n10798(x10798, x6481, x4713);
  nand n10799(x10799, x10798, x10797);
  nand n10800(x10800, x2258, x4583);
  nand n10801(x10801, x6481, x4453);
  nand n10802(x10802, x10801, x10800);
  nand n10803(x10803, x2261, x10793);
  nand n10804(x10804, x6494, x10796);
  nand n10805(x10805, x10804, x10803);
  nand n10806(x10806, x2261, x10799);
  nand n10807(x10807, x6494, x10802);
  nand n10808(x10808, x10807, x10806);
  nand n10809(x10809, x2264, x10805);
  nand n10810(x10810, x6501, x10808);
  nand n10811(x10811, x10810, x10809);
  nand n10812(x10812, x2258, x5367);
  nand n10813(x10813, x6481, x5237);
  nand n10814(x10814, x10813, x10812);
  nand n10815(x10815, x2258, x5107);
  nand n10816(x10816, x6481, x4977);
  nand n10817(x10817, x10816, x10815);
  nand n10818(x10818, x2258, x4847);
  nand n10819(x10819, x6481, x4717);
  nand n10820(x10820, x10819, x10818);
  nand n10821(x10821, x2258, x4587);
  nand n10822(x10822, x6481, x4457);
  nand n10823(x10823, x10822, x10821);
  nand n10824(x10824, x2261, x10814);
  nand n10825(x10825, x6494, x10817);
  nand n10826(x10826, x10825, x10824);
  nand n10827(x10827, x2261, x10820);
  nand n10828(x10828, x6494, x10823);
  nand n10829(x10829, x10828, x10827);
  nand n10830(x10830, x2264, x10826);
  nand n10831(x10831, x6501, x10829);
  nand n10832(x10832, x10831, x10830);
  nand n10833(x10833, x2258, x5371);
  nand n10834(x10834, x6481, x5241);
  nand n10835(x10835, x10834, x10833);
  nand n10836(x10836, x2258, x5111);
  nand n10837(x10837, x6481, x4981);
  nand n10838(x10838, x10837, x10836);
  nand n10839(x10839, x2258, x4851);
  nand n10840(x10840, x6481, x4721);
  nand n10841(x10841, x10840, x10839);
  nand n10842(x10842, x2258, x4591);
  nand n10843(x10843, x6481, x4461);
  nand n10844(x10844, x10843, x10842);
  nand n10845(x10845, x2261, x10835);
  nand n10846(x10846, x6494, x10838);
  nand n10847(x10847, x10846, x10845);
  nand n10848(x10848, x2261, x10841);
  nand n10849(x10849, x6494, x10844);
  nand n10850(x10850, x10849, x10848);
  nand n10851(x10851, x2264, x10847);
  nand n10852(x10852, x6501, x10850);
  nand n10853(x10853, x10852, x10851);
  nand n10854(x10854, x2258, x5375);
  nand n10855(x10855, x6481, x5245);
  nand n10856(x10856, x10855, x10854);
  nand n10857(x10857, x2258, x5115);
  nand n10858(x10858, x6481, x4985);
  nand n10859(x10859, x10858, x10857);
  nand n10860(x10860, x2258, x4855);
  nand n10861(x10861, x6481, x4725);
  nand n10862(x10862, x10861, x10860);
  nand n10863(x10863, x2258, x4595);
  nand n10864(x10864, x6481, x4465);
  nand n10865(x10865, x10864, x10863);
  nand n10866(x10866, x2261, x10856);
  nand n10867(x10867, x6494, x10859);
  nand n10868(x10868, x10867, x10866);
  nand n10869(x10869, x2261, x10862);
  nand n10870(x10870, x6494, x10865);
  nand n10871(x10871, x10870, x10869);
  nand n10872(x10872, x2264, x10868);
  nand n10873(x10873, x6501, x10871);
  nand n10874(x10874, x10873, x10872);
  nand n10875(x10875, x2258, x5379);
  nand n10876(x10876, x6481, x5249);
  nand n10877(x10877, x10876, x10875);
  nand n10878(x10878, x2258, x5119);
  nand n10879(x10879, x6481, x4989);
  nand n10880(x10880, x10879, x10878);
  nand n10881(x10881, x2258, x4859);
  nand n10882(x10882, x6481, x4729);
  nand n10883(x10883, x10882, x10881);
  nand n10884(x10884, x2258, x4599);
  nand n10885(x10885, x6481, x4469);
  nand n10886(x10886, x10885, x10884);
  nand n10887(x10887, x2261, x10877);
  nand n10888(x10888, x6494, x10880);
  nand n10889(x10889, x10888, x10887);
  nand n10890(x10890, x2261, x10883);
  nand n10891(x10891, x6494, x10886);
  nand n10892(x10892, x10891, x10890);
  nand n10893(x10893, x2264, x10889);
  nand n10894(x10894, x6501, x10892);
  nand n10895(x10895, x10894, x10893);
  nand n10896(x10896, x2258, x5383);
  nand n10897(x10897, x6481, x5253);
  nand n10898(x10898, x10897, x10896);
  nand n10899(x10899, x2258, x5123);
  nand n10900(x10900, x6481, x4993);
  nand n10901(x10901, x10900, x10899);
  nand n10902(x10902, x2258, x4863);
  nand n10903(x10903, x6481, x4733);
  nand n10904(x10904, x10903, x10902);
  nand n10905(x10905, x2258, x4603);
  nand n10906(x10906, x6481, x4473);
  nand n10907(x10907, x10906, x10905);
  nand n10908(x10908, x2261, x10898);
  nand n10909(x10909, x6494, x10901);
  nand n10910(x10910, x10909, x10908);
  nand n10911(x10911, x2261, x10904);
  nand n10912(x10912, x6494, x10907);
  nand n10913(x10913, x10912, x10911);
  nand n10914(x10914, x2264, x10910);
  nand n10915(x10915, x6501, x10913);
  nand n10916(x10916, x10915, x10914);
  nand n10917(x10917, x2258, x5387);
  nand n10918(x10918, x6481, x5257);
  nand n10919(x10919, x10918, x10917);
  nand n10920(x10920, x2258, x5127);
  nand n10921(x10921, x6481, x4997);
  nand n10922(x10922, x10921, x10920);
  nand n10923(x10923, x2258, x4867);
  nand n10924(x10924, x6481, x4737);
  nand n10925(x10925, x10924, x10923);
  nand n10926(x10926, x2258, x4607);
  nand n10927(x10927, x6481, x4477);
  nand n10928(x10928, x10927, x10926);
  nand n10929(x10929, x2261, x10919);
  nand n10930(x10930, x6494, x10922);
  nand n10931(x10931, x10930, x10929);
  nand n10932(x10932, x2261, x10925);
  nand n10933(x10933, x6494, x10928);
  nand n10934(x10934, x10933, x10932);
  nand n10935(x10935, x2264, x10931);
  nand n10936(x10936, x6501, x10934);
  nand n10937(x10937, x10936, x10935);
  nand n10938(x10938, x2258, x5391);
  nand n10939(x10939, x6481, x5261);
  nand n10940(x10940, x10939, x10938);
  nand n10941(x10941, x2258, x5131);
  nand n10942(x10942, x6481, x5001);
  nand n10943(x10943, x10942, x10941);
  nand n10944(x10944, x2258, x4871);
  nand n10945(x10945, x6481, x4741);
  nand n10946(x10946, x10945, x10944);
  nand n10947(x10947, x2258, x4611);
  nand n10948(x10948, x6481, x4481);
  nand n10949(x10949, x10948, x10947);
  nand n10950(x10950, x2261, x10940);
  nand n10951(x10951, x6494, x10943);
  nand n10952(x10952, x10951, x10950);
  nand n10953(x10953, x2261, x10946);
  nand n10954(x10954, x6494, x10949);
  nand n10955(x10955, x10954, x10953);
  nand n10956(x10956, x2264, x10952);
  nand n10957(x10957, x6501, x10955);
  nand n10958(x10958, x10957, x10956);
  nand n10959(x10959, x2258, x5395);
  nand n10960(x10960, x6481, x5265);
  nand n10961(x10961, x10960, x10959);
  nand n10962(x10962, x2258, x5135);
  nand n10963(x10963, x6481, x5005);
  nand n10964(x10964, x10963, x10962);
  nand n10965(x10965, x2258, x4875);
  nand n10966(x10966, x6481, x4745);
  nand n10967(x10967, x10966, x10965);
  nand n10968(x10968, x2258, x4615);
  nand n10969(x10969, x6481, x4485);
  nand n10970(x10970, x10969, x10968);
  nand n10971(x10971, x2261, x10961);
  nand n10972(x10972, x6494, x10964);
  nand n10973(x10973, x10972, x10971);
  nand n10974(x10974, x2261, x10967);
  nand n10975(x10975, x6494, x10970);
  nand n10976(x10976, x10975, x10974);
  nand n10977(x10977, x2264, x10973);
  nand n10978(x10978, x6501, x10976);
  nand n10979(x10979, x10978, x10977);
  nand n10980(x10980, x2258, x5399);
  nand n10981(x10981, x6481, x5269);
  nand n10982(x10982, x10981, x10980);
  nand n10983(x10983, x2258, x5139);
  nand n10984(x10984, x6481, x5009);
  nand n10985(x10985, x10984, x10983);
  nand n10986(x10986, x2258, x4879);
  nand n10987(x10987, x6481, x4749);
  nand n10988(x10988, x10987, x10986);
  nand n10989(x10989, x2258, x4619);
  nand n10990(x10990, x6481, x4489);
  nand n10991(x10991, x10990, x10989);
  nand n10992(x10992, x2261, x10982);
  nand n10993(x10993, x6494, x10985);
  nand n10994(x10994, x10993, x10992);
  nand n10995(x10995, x2261, x10988);
  nand n10996(x10996, x6494, x10991);
  nand n10997(x10997, x10996, x10995);
  nand n10998(x10998, x2264, x10994);
  nand n10999(x10999, x6501, x10997);
  nand n11000(x11000, x10999, x10998);
  nand n11001(x11001, x2258, x5403);
  nand n11002(x11002, x6481, x5273);
  nand n11003(x11003, x11002, x11001);
  nand n11004(x11004, x2258, x5143);
  nand n11005(x11005, x6481, x5013);
  nand n11006(x11006, x11005, x11004);
  nand n11007(x11007, x2258, x4883);
  nand n11008(x11008, x6481, x4753);
  nand n11009(x11009, x11008, x11007);
  nand n11010(x11010, x2258, x4623);
  nand n11011(x11011, x6481, x4493);
  nand n11012(x11012, x11011, x11010);
  nand n11013(x11013, x2261, x11003);
  nand n11014(x11014, x6494, x11006);
  nand n11015(x11015, x11014, x11013);
  nand n11016(x11016, x2261, x11009);
  nand n11017(x11017, x6494, x11012);
  nand n11018(x11018, x11017, x11016);
  nand n11019(x11019, x2264, x11015);
  nand n11020(x11020, x6501, x11018);
  nand n11021(x11021, x11020, x11019);
  nand n11022(x11022, x2258, x5407);
  nand n11023(x11023, x6481, x5277);
  nand n11024(x11024, x11023, x11022);
  nand n11025(x11025, x2258, x5147);
  nand n11026(x11026, x6481, x5017);
  nand n11027(x11027, x11026, x11025);
  nand n11028(x11028, x2258, x4887);
  nand n11029(x11029, x6481, x4757);
  nand n11030(x11030, x11029, x11028);
  nand n11031(x11031, x2258, x4627);
  nand n11032(x11032, x6481, x4497);
  nand n11033(x11033, x11032, x11031);
  nand n11034(x11034, x2261, x11024);
  nand n11035(x11035, x6494, x11027);
  nand n11036(x11036, x11035, x11034);
  nand n11037(x11037, x2261, x11030);
  nand n11038(x11038, x6494, x11033);
  nand n11039(x11039, x11038, x11037);
  nand n11040(x11040, x2264, x11036);
  nand n11041(x11041, x6501, x11039);
  nand n11042(x11042, x11041, x11040);
  nand n11043(x11043, x2258, x5411);
  nand n11044(x11044, x6481, x5281);
  nand n11045(x11045, x11044, x11043);
  nand n11046(x11046, x2258, x5151);
  nand n11047(x11047, x6481, x5021);
  nand n11048(x11048, x11047, x11046);
  nand n11049(x11049, x2258, x4891);
  nand n11050(x11050, x6481, x4761);
  nand n11051(x11051, x11050, x11049);
  nand n11052(x11052, x2258, x4631);
  nand n11053(x11053, x6481, x4501);
  nand n11054(x11054, x11053, x11052);
  nand n11055(x11055, x2261, x11045);
  nand n11056(x11056, x6494, x11048);
  nand n11057(x11057, x11056, x11055);
  nand n11058(x11058, x2261, x11051);
  nand n11059(x11059, x6494, x11054);
  nand n11060(x11060, x11059, x11058);
  nand n11061(x11061, x2264, x11057);
  nand n11062(x11062, x6501, x11060);
  nand n11063(x11063, x11062, x11061);
  nand n11064(x11064, x2258, x5415);
  nand n11065(x11065, x6481, x5285);
  nand n11066(x11066, x11065, x11064);
  nand n11067(x11067, x2258, x5155);
  nand n11068(x11068, x6481, x5025);
  nand n11069(x11069, x11068, x11067);
  nand n11070(x11070, x2258, x4895);
  nand n11071(x11071, x6481, x4765);
  nand n11072(x11072, x11071, x11070);
  nand n11073(x11073, x2258, x4635);
  nand n11074(x11074, x6481, x4505);
  nand n11075(x11075, x11074, x11073);
  nand n11076(x11076, x2261, x11066);
  nand n11077(x11077, x6494, x11069);
  nand n11078(x11078, x11077, x11076);
  nand n11079(x11079, x2261, x11072);
  nand n11080(x11080, x6494, x11075);
  nand n11081(x11081, x11080, x11079);
  nand n11082(x11082, x2264, x11078);
  nand n11083(x11083, x6501, x11081);
  nand n11084(x11084, x11083, x11082);
  nand n11085(x11085, x2258, x5419);
  nand n11086(x11086, x6481, x5289);
  nand n11087(x11087, x11086, x11085);
  nand n11088(x11088, x2258, x5159);
  nand n11089(x11089, x6481, x5029);
  nand n11090(x11090, x11089, x11088);
  nand n11091(x11091, x2258, x4899);
  nand n11092(x11092, x6481, x4769);
  nand n11093(x11093, x11092, x11091);
  nand n11094(x11094, x2258, x4639);
  nand n11095(x11095, x6481, x4509);
  nand n11096(x11096, x11095, x11094);
  nand n11097(x11097, x2261, x11087);
  nand n11098(x11098, x6494, x11090);
  nand n11099(x11099, x11098, x11097);
  nand n11100(x11100, x2261, x11093);
  nand n11101(x11101, x6494, x11096);
  nand n11102(x11102, x11101, x11100);
  nand n11103(x11103, x2264, x11099);
  nand n11104(x11104, x6501, x11102);
  nand n11105(x11105, x11104, x11103);
  nand n11106(x11106, x2258, x5423);
  nand n11107(x11107, x6481, x5293);
  nand n11108(x11108, x11107, x11106);
  nand n11109(x11109, x2258, x5163);
  nand n11110(x11110, x6481, x5033);
  nand n11111(x11111, x11110, x11109);
  nand n11112(x11112, x2258, x4903);
  nand n11113(x11113, x6481, x4773);
  nand n11114(x11114, x11113, x11112);
  nand n11115(x11115, x2258, x4643);
  nand n11116(x11116, x6481, x4513);
  nand n11117(x11117, x11116, x11115);
  nand n11118(x11118, x2261, x11108);
  nand n11119(x11119, x6494, x11111);
  nand n11120(x11120, x11119, x11118);
  nand n11121(x11121, x2261, x11114);
  nand n11122(x11122, x6494, x11117);
  nand n11123(x11123, x11122, x11121);
  nand n11124(x11124, x2264, x11120);
  nand n11125(x11125, x6501, x11123);
  nand n11126(x11126, x11125, x11124);
  nand n11127(x11127, x2258, x5427);
  nand n11128(x11128, x6481, x5297);
  nand n11129(x11129, x11128, x11127);
  nand n11130(x11130, x2258, x5167);
  nand n11131(x11131, x6481, x5037);
  nand n11132(x11132, x11131, x11130);
  nand n11133(x11133, x2258, x4907);
  nand n11134(x11134, x6481, x4777);
  nand n11135(x11135, x11134, x11133);
  nand n11136(x11136, x2258, x4647);
  nand n11137(x11137, x6481, x4517);
  nand n11138(x11138, x11137, x11136);
  nand n11139(x11139, x2261, x11129);
  nand n11140(x11140, x6494, x11132);
  nand n11141(x11141, x11140, x11139);
  nand n11142(x11142, x2261, x11135);
  nand n11143(x11143, x6494, x11138);
  nand n11144(x11144, x11143, x11142);
  nand n11145(x11145, x2264, x11141);
  nand n11146(x11146, x6501, x11144);
  nand n11147(x11147, x11146, x11145);
  nand n11148(x11148, x2258, x5431);
  nand n11149(x11149, x6481, x5301);
  nand n11150(x11150, x11149, x11148);
  nand n11151(x11151, x2258, x5171);
  nand n11152(x11152, x6481, x5041);
  nand n11153(x11153, x11152, x11151);
  nand n11154(x11154, x2258, x4911);
  nand n11155(x11155, x6481, x4781);
  nand n11156(x11156, x11155, x11154);
  nand n11157(x11157, x2258, x4651);
  nand n11158(x11158, x6481, x4521);
  nand n11159(x11159, x11158, x11157);
  nand n11160(x11160, x2261, x11150);
  nand n11161(x11161, x6494, x11153);
  nand n11162(x11162, x11161, x11160);
  nand n11163(x11163, x2261, x11156);
  nand n11164(x11164, x6494, x11159);
  nand n11165(x11165, x11164, x11163);
  nand n11166(x11166, x2264, x11162);
  nand n11167(x11167, x6501, x11165);
  nand n11168(x11168, x11167, x11166);
  nand n11169(x11169, x2258, x5435);
  nand n11170(x11170, x6481, x5305);
  nand n11171(x11171, x11170, x11169);
  nand n11172(x11172, x2258, x5175);
  nand n11173(x11173, x6481, x5045);
  nand n11174(x11174, x11173, x11172);
  nand n11175(x11175, x2258, x4915);
  nand n11176(x11176, x6481, x4785);
  nand n11177(x11177, x11176, x11175);
  nand n11178(x11178, x2258, x4655);
  nand n11179(x11179, x6481, x4525);
  nand n11180(x11180, x11179, x11178);
  nand n11181(x11181, x2261, x11171);
  nand n11182(x11182, x6494, x11174);
  nand n11183(x11183, x11182, x11181);
  nand n11184(x11184, x2261, x11177);
  nand n11185(x11185, x6494, x11180);
  nand n11186(x11186, x11185, x11184);
  nand n11187(x11187, x2264, x11183);
  nand n11188(x11188, x6501, x11186);
  nand n11189(x11189, x11188, x11187);
  nand n11190(x11190, x2269, x5311);
  nand n11191(x11191, x7156, x5181);
  nand n11192(x11192, x11191, x11190);
  nand n11193(x11193, x2269, x5051);
  nand n11194(x11194, x7156, x4921);
  nand n11195(x11195, x11194, x11193);
  nand n11196(x11196, x2269, x4791);
  nand n11197(x11197, x7156, x4661);
  nand n11198(x11198, x11197, x11196);
  nand n11199(x11199, x2269, x4531);
  nand n11200(x11200, x7156, x4399);
  nand n11201(x11201, x11200, x11199);
  nand n11202(x11202, x2272, x11192);
  nand n11203(x11203, x7169, x11195);
  nand n11204(x11204, x11203, x11202);
  nand n11205(x11205, x2272, x11198);
  nand n11206(x11206, x7169, x11201);
  nand n11207(x11207, x11206, x11205);
  nand n11208(x11208, x2275, x11204);
  nand n11209(x11209, x7176, x11207);
  nand n11210(x11210, x11209, x11208);
  nand n11211(x11211, x2269, x5315);
  nand n11212(x11212, x7156, x5185);
  nand n11213(x11213, x11212, x11211);
  nand n11214(x11214, x2269, x5055);
  nand n11215(x11215, x7156, x4925);
  nand n11216(x11216, x11215, x11214);
  nand n11217(x11217, x2269, x4795);
  nand n11218(x11218, x7156, x4665);
  nand n11219(x11219, x11218, x11217);
  nand n11220(x11220, x2269, x4535);
  nand n11221(x11221, x7156, x4405);
  nand n11222(x11222, x11221, x11220);
  nand n11223(x11223, x2272, x11213);
  nand n11224(x11224, x7169, x11216);
  nand n11225(x11225, x11224, x11223);
  nand n11226(x11226, x2272, x11219);
  nand n11227(x11227, x7169, x11222);
  nand n11228(x11228, x11227, x11226);
  nand n11229(x11229, x2275, x11225);
  nand n11230(x11230, x7176, x11228);
  nand n11231(x11231, x11230, x11229);
  nand n11232(x11232, x2269, x5319);
  nand n11233(x11233, x7156, x5189);
  nand n11234(x11234, x11233, x11232);
  nand n11235(x11235, x2269, x5059);
  nand n11236(x11236, x7156, x4929);
  nand n11237(x11237, x11236, x11235);
  nand n11238(x11238, x2269, x4799);
  nand n11239(x11239, x7156, x4669);
  nand n11240(x11240, x11239, x11238);
  nand n11241(x11241, x2269, x4539);
  nand n11242(x11242, x7156, x4409);
  nand n11243(x11243, x11242, x11241);
  nand n11244(x11244, x2272, x11234);
  nand n11245(x11245, x7169, x11237);
  nand n11246(x11246, x11245, x11244);
  nand n11247(x11247, x2272, x11240);
  nand n11248(x11248, x7169, x11243);
  nand n11249(x11249, x11248, x11247);
  nand n11250(x11250, x2275, x11246);
  nand n11251(x11251, x7176, x11249);
  nand n11252(x11252, x11251, x11250);
  nand n11253(x11253, x2269, x5323);
  nand n11254(x11254, x7156, x5193);
  nand n11255(x11255, x11254, x11253);
  nand n11256(x11256, x2269, x5063);
  nand n11257(x11257, x7156, x4933);
  nand n11258(x11258, x11257, x11256);
  nand n11259(x11259, x2269, x4803);
  nand n11260(x11260, x7156, x4673);
  nand n11261(x11261, x11260, x11259);
  nand n11262(x11262, x2269, x4543);
  nand n11263(x11263, x7156, x4413);
  nand n11264(x11264, x11263, x11262);
  nand n11265(x11265, x2272, x11255);
  nand n11266(x11266, x7169, x11258);
  nand n11267(x11267, x11266, x11265);
  nand n11268(x11268, x2272, x11261);
  nand n11269(x11269, x7169, x11264);
  nand n11270(x11270, x11269, x11268);
  nand n11271(x11271, x2275, x11267);
  nand n11272(x11272, x7176, x11270);
  nand n11273(x11273, x11272, x11271);
  nand n11274(x11274, x2269, x5327);
  nand n11275(x11275, x7156, x5197);
  nand n11276(x11276, x11275, x11274);
  nand n11277(x11277, x2269, x5067);
  nand n11278(x11278, x7156, x4937);
  nand n11279(x11279, x11278, x11277);
  nand n11280(x11280, x2269, x4807);
  nand n11281(x11281, x7156, x4677);
  nand n11282(x11282, x11281, x11280);
  nand n11283(x11283, x2269, x4547);
  nand n11284(x11284, x7156, x4417);
  nand n11285(x11285, x11284, x11283);
  nand n11286(x11286, x2272, x11276);
  nand n11287(x11287, x7169, x11279);
  nand n11288(x11288, x11287, x11286);
  nand n11289(x11289, x2272, x11282);
  nand n11290(x11290, x7169, x11285);
  nand n11291(x11291, x11290, x11289);
  nand n11292(x11292, x2275, x11288);
  nand n11293(x11293, x7176, x11291);
  nand n11294(x11294, x11293, x11292);
  nand n11295(x11295, x2269, x5331);
  nand n11296(x11296, x7156, x5201);
  nand n11297(x11297, x11296, x11295);
  nand n11298(x11298, x2269, x5071);
  nand n11299(x11299, x7156, x4941);
  nand n11300(x11300, x11299, x11298);
  nand n11301(x11301, x2269, x4811);
  nand n11302(x11302, x7156, x4681);
  nand n11303(x11303, x11302, x11301);
  nand n11304(x11304, x2269, x4551);
  nand n11305(x11305, x7156, x4421);
  nand n11306(x11306, x11305, x11304);
  nand n11307(x11307, x2272, x11297);
  nand n11308(x11308, x7169, x11300);
  nand n11309(x11309, x11308, x11307);
  nand n11310(x11310, x2272, x11303);
  nand n11311(x11311, x7169, x11306);
  nand n11312(x11312, x11311, x11310);
  nand n11313(x11313, x2275, x11309);
  nand n11314(x11314, x7176, x11312);
  nand n11315(x11315, x11314, x11313);
  nand n11316(x11316, x2269, x5335);
  nand n11317(x11317, x7156, x5205);
  nand n11318(x11318, x11317, x11316);
  nand n11319(x11319, x2269, x5075);
  nand n11320(x11320, x7156, x4945);
  nand n11321(x11321, x11320, x11319);
  nand n11322(x11322, x2269, x4815);
  nand n11323(x11323, x7156, x4685);
  nand n11324(x11324, x11323, x11322);
  nand n11325(x11325, x2269, x4555);
  nand n11326(x11326, x7156, x4425);
  nand n11327(x11327, x11326, x11325);
  nand n11328(x11328, x2272, x11318);
  nand n11329(x11329, x7169, x11321);
  nand n11330(x11330, x11329, x11328);
  nand n11331(x11331, x2272, x11324);
  nand n11332(x11332, x7169, x11327);
  nand n11333(x11333, x11332, x11331);
  nand n11334(x11334, x2275, x11330);
  nand n11335(x11335, x7176, x11333);
  nand n11336(x11336, x11335, x11334);
  nand n11337(x11337, x2269, x5339);
  nand n11338(x11338, x7156, x5209);
  nand n11339(x11339, x11338, x11337);
  nand n11340(x11340, x2269, x5079);
  nand n11341(x11341, x7156, x4949);
  nand n11342(x11342, x11341, x11340);
  nand n11343(x11343, x2269, x4819);
  nand n11344(x11344, x7156, x4689);
  nand n11345(x11345, x11344, x11343);
  nand n11346(x11346, x2269, x4559);
  nand n11347(x11347, x7156, x4429);
  nand n11348(x11348, x11347, x11346);
  nand n11349(x11349, x2272, x11339);
  nand n11350(x11350, x7169, x11342);
  nand n11351(x11351, x11350, x11349);
  nand n11352(x11352, x2272, x11345);
  nand n11353(x11353, x7169, x11348);
  nand n11354(x11354, x11353, x11352);
  nand n11355(x11355, x2275, x11351);
  nand n11356(x11356, x7176, x11354);
  nand n11357(x11357, x11356, x11355);
  nand n11358(x11358, x2269, x5343);
  nand n11359(x11359, x7156, x5213);
  nand n11360(x11360, x11359, x11358);
  nand n11361(x11361, x2269, x5083);
  nand n11362(x11362, x7156, x4953);
  nand n11363(x11363, x11362, x11361);
  nand n11364(x11364, x2269, x4823);
  nand n11365(x11365, x7156, x4693);
  nand n11366(x11366, x11365, x11364);
  nand n11367(x11367, x2269, x4563);
  nand n11368(x11368, x7156, x4433);
  nand n11369(x11369, x11368, x11367);
  nand n11370(x11370, x2272, x11360);
  nand n11371(x11371, x7169, x11363);
  nand n11372(x11372, x11371, x11370);
  nand n11373(x11373, x2272, x11366);
  nand n11374(x11374, x7169, x11369);
  nand n11375(x11375, x11374, x11373);
  nand n11376(x11376, x2275, x11372);
  nand n11377(x11377, x7176, x11375);
  nand n11378(x11378, x11377, x11376);
  nand n11379(x11379, x2269, x5347);
  nand n11380(x11380, x7156, x5217);
  nand n11381(x11381, x11380, x11379);
  nand n11382(x11382, x2269, x5087);
  nand n11383(x11383, x7156, x4957);
  nand n11384(x11384, x11383, x11382);
  nand n11385(x11385, x2269, x4827);
  nand n11386(x11386, x7156, x4697);
  nand n11387(x11387, x11386, x11385);
  nand n11388(x11388, x2269, x4567);
  nand n11389(x11389, x7156, x4437);
  nand n11390(x11390, x11389, x11388);
  nand n11391(x11391, x2272, x11381);
  nand n11392(x11392, x7169, x11384);
  nand n11393(x11393, x11392, x11391);
  nand n11394(x11394, x2272, x11387);
  nand n11395(x11395, x7169, x11390);
  nand n11396(x11396, x11395, x11394);
  nand n11397(x11397, x2275, x11393);
  nand n11398(x11398, x7176, x11396);
  nand n11399(x11399, x11398, x11397);
  nand n11400(x11400, x2269, x5351);
  nand n11401(x11401, x7156, x5221);
  nand n11402(x11402, x11401, x11400);
  nand n11403(x11403, x2269, x5091);
  nand n11404(x11404, x7156, x4961);
  nand n11405(x11405, x11404, x11403);
  nand n11406(x11406, x2269, x4831);
  nand n11407(x11407, x7156, x4701);
  nand n11408(x11408, x11407, x11406);
  nand n11409(x11409, x2269, x4571);
  nand n11410(x11410, x7156, x4441);
  nand n11411(x11411, x11410, x11409);
  nand n11412(x11412, x2272, x11402);
  nand n11413(x11413, x7169, x11405);
  nand n11414(x11414, x11413, x11412);
  nand n11415(x11415, x2272, x11408);
  nand n11416(x11416, x7169, x11411);
  nand n11417(x11417, x11416, x11415);
  nand n11418(x11418, x2275, x11414);
  nand n11419(x11419, x7176, x11417);
  nand n11420(x11420, x11419, x11418);
  nand n11421(x11421, x2269, x5355);
  nand n11422(x11422, x7156, x5225);
  nand n11423(x11423, x11422, x11421);
  nand n11424(x11424, x2269, x5095);
  nand n11425(x11425, x7156, x4965);
  nand n11426(x11426, x11425, x11424);
  nand n11427(x11427, x2269, x4835);
  nand n11428(x11428, x7156, x4705);
  nand n11429(x11429, x11428, x11427);
  nand n11430(x11430, x2269, x4575);
  nand n11431(x11431, x7156, x4445);
  nand n11432(x11432, x11431, x11430);
  nand n11433(x11433, x2272, x11423);
  nand n11434(x11434, x7169, x11426);
  nand n11435(x11435, x11434, x11433);
  nand n11436(x11436, x2272, x11429);
  nand n11437(x11437, x7169, x11432);
  nand n11438(x11438, x11437, x11436);
  nand n11439(x11439, x2275, x11435);
  nand n11440(x11440, x7176, x11438);
  nand n11441(x11441, x11440, x11439);
  nand n11442(x11442, x2269, x5359);
  nand n11443(x11443, x7156, x5229);
  nand n11444(x11444, x11443, x11442);
  nand n11445(x11445, x2269, x5099);
  nand n11446(x11446, x7156, x4969);
  nand n11447(x11447, x11446, x11445);
  nand n11448(x11448, x2269, x4839);
  nand n11449(x11449, x7156, x4709);
  nand n11450(x11450, x11449, x11448);
  nand n11451(x11451, x2269, x4579);
  nand n11452(x11452, x7156, x4449);
  nand n11453(x11453, x11452, x11451);
  nand n11454(x11454, x2272, x11444);
  nand n11455(x11455, x7169, x11447);
  nand n11456(x11456, x11455, x11454);
  nand n11457(x11457, x2272, x11450);
  nand n11458(x11458, x7169, x11453);
  nand n11459(x11459, x11458, x11457);
  nand n11460(x11460, x2275, x11456);
  nand n11461(x11461, x7176, x11459);
  nand n11462(x11462, x11461, x11460);
  nand n11463(x11463, x2269, x5363);
  nand n11464(x11464, x7156, x5233);
  nand n11465(x11465, x11464, x11463);
  nand n11466(x11466, x2269, x5103);
  nand n11467(x11467, x7156, x4973);
  nand n11468(x11468, x11467, x11466);
  nand n11469(x11469, x2269, x4843);
  nand n11470(x11470, x7156, x4713);
  nand n11471(x11471, x11470, x11469);
  nand n11472(x11472, x2269, x4583);
  nand n11473(x11473, x7156, x4453);
  nand n11474(x11474, x11473, x11472);
  nand n11475(x11475, x2272, x11465);
  nand n11476(x11476, x7169, x11468);
  nand n11477(x11477, x11476, x11475);
  nand n11478(x11478, x2272, x11471);
  nand n11479(x11479, x7169, x11474);
  nand n11480(x11480, x11479, x11478);
  nand n11481(x11481, x2275, x11477);
  nand n11482(x11482, x7176, x11480);
  nand n11483(x11483, x11482, x11481);
  nand n11484(x11484, x2269, x5367);
  nand n11485(x11485, x7156, x5237);
  nand n11486(x11486, x11485, x11484);
  nand n11487(x11487, x2269, x5107);
  nand n11488(x11488, x7156, x4977);
  nand n11489(x11489, x11488, x11487);
  nand n11490(x11490, x2269, x4847);
  nand n11491(x11491, x7156, x4717);
  nand n11492(x11492, x11491, x11490);
  nand n11493(x11493, x2269, x4587);
  nand n11494(x11494, x7156, x4457);
  nand n11495(x11495, x11494, x11493);
  nand n11496(x11496, x2272, x11486);
  nand n11497(x11497, x7169, x11489);
  nand n11498(x11498, x11497, x11496);
  nand n11499(x11499, x2272, x11492);
  nand n11500(x11500, x7169, x11495);
  nand n11501(x11501, x11500, x11499);
  nand n11502(x11502, x2275, x11498);
  nand n11503(x11503, x7176, x11501);
  nand n11504(x11504, x11503, x11502);
  nand n11505(x11505, x2269, x5371);
  nand n11506(x11506, x7156, x5241);
  nand n11507(x11507, x11506, x11505);
  nand n11508(x11508, x2269, x5111);
  nand n11509(x11509, x7156, x4981);
  nand n11510(x11510, x11509, x11508);
  nand n11511(x11511, x2269, x4851);
  nand n11512(x11512, x7156, x4721);
  nand n11513(x11513, x11512, x11511);
  nand n11514(x11514, x2269, x4591);
  nand n11515(x11515, x7156, x4461);
  nand n11516(x11516, x11515, x11514);
  nand n11517(x11517, x2272, x11507);
  nand n11518(x11518, x7169, x11510);
  nand n11519(x11519, x11518, x11517);
  nand n11520(x11520, x2272, x11513);
  nand n11521(x11521, x7169, x11516);
  nand n11522(x11522, x11521, x11520);
  nand n11523(x11523, x2275, x11519);
  nand n11524(x11524, x7176, x11522);
  nand n11525(x11525, x11524, x11523);
  nand n11526(x11526, x2269, x5375);
  nand n11527(x11527, x7156, x5245);
  nand n11528(x11528, x11527, x11526);
  nand n11529(x11529, x2269, x5115);
  nand n11530(x11530, x7156, x4985);
  nand n11531(x11531, x11530, x11529);
  nand n11532(x11532, x2269, x4855);
  nand n11533(x11533, x7156, x4725);
  nand n11534(x11534, x11533, x11532);
  nand n11535(x11535, x2269, x4595);
  nand n11536(x11536, x7156, x4465);
  nand n11537(x11537, x11536, x11535);
  nand n11538(x11538, x2272, x11528);
  nand n11539(x11539, x7169, x11531);
  nand n11540(x11540, x11539, x11538);
  nand n11541(x11541, x2272, x11534);
  nand n11542(x11542, x7169, x11537);
  nand n11543(x11543, x11542, x11541);
  nand n11544(x11544, x2275, x11540);
  nand n11545(x11545, x7176, x11543);
  nand n11546(x11546, x11545, x11544);
  nand n11547(x11547, x2269, x5379);
  nand n11548(x11548, x7156, x5249);
  nand n11549(x11549, x11548, x11547);
  nand n11550(x11550, x2269, x5119);
  nand n11551(x11551, x7156, x4989);
  nand n11552(x11552, x11551, x11550);
  nand n11553(x11553, x2269, x4859);
  nand n11554(x11554, x7156, x4729);
  nand n11555(x11555, x11554, x11553);
  nand n11556(x11556, x2269, x4599);
  nand n11557(x11557, x7156, x4469);
  nand n11558(x11558, x11557, x11556);
  nand n11559(x11559, x2272, x11549);
  nand n11560(x11560, x7169, x11552);
  nand n11561(x11561, x11560, x11559);
  nand n11562(x11562, x2272, x11555);
  nand n11563(x11563, x7169, x11558);
  nand n11564(x11564, x11563, x11562);
  nand n11565(x11565, x2275, x11561);
  nand n11566(x11566, x7176, x11564);
  nand n11567(x11567, x11566, x11565);
  nand n11568(x11568, x2269, x5383);
  nand n11569(x11569, x7156, x5253);
  nand n11570(x11570, x11569, x11568);
  nand n11571(x11571, x2269, x5123);
  nand n11572(x11572, x7156, x4993);
  nand n11573(x11573, x11572, x11571);
  nand n11574(x11574, x2269, x4863);
  nand n11575(x11575, x7156, x4733);
  nand n11576(x11576, x11575, x11574);
  nand n11577(x11577, x2269, x4603);
  nand n11578(x11578, x7156, x4473);
  nand n11579(x11579, x11578, x11577);
  nand n11580(x11580, x2272, x11570);
  nand n11581(x11581, x7169, x11573);
  nand n11582(x11582, x11581, x11580);
  nand n11583(x11583, x2272, x11576);
  nand n11584(x11584, x7169, x11579);
  nand n11585(x11585, x11584, x11583);
  nand n11586(x11586, x2275, x11582);
  nand n11587(x11587, x7176, x11585);
  nand n11588(x11588, x11587, x11586);
  nand n11589(x11589, x2269, x5387);
  nand n11590(x11590, x7156, x5257);
  nand n11591(x11591, x11590, x11589);
  nand n11592(x11592, x2269, x5127);
  nand n11593(x11593, x7156, x4997);
  nand n11594(x11594, x11593, x11592);
  nand n11595(x11595, x2269, x4867);
  nand n11596(x11596, x7156, x4737);
  nand n11597(x11597, x11596, x11595);
  nand n11598(x11598, x2269, x4607);
  nand n11599(x11599, x7156, x4477);
  nand n11600(x11600, x11599, x11598);
  nand n11601(x11601, x2272, x11591);
  nand n11602(x11602, x7169, x11594);
  nand n11603(x11603, x11602, x11601);
  nand n11604(x11604, x2272, x11597);
  nand n11605(x11605, x7169, x11600);
  nand n11606(x11606, x11605, x11604);
  nand n11607(x11607, x2275, x11603);
  nand n11608(x11608, x7176, x11606);
  nand n11609(x11609, x11608, x11607);
  nand n11610(x11610, x2269, x5391);
  nand n11611(x11611, x7156, x5261);
  nand n11612(x11612, x11611, x11610);
  nand n11613(x11613, x2269, x5131);
  nand n11614(x11614, x7156, x5001);
  nand n11615(x11615, x11614, x11613);
  nand n11616(x11616, x2269, x4871);
  nand n11617(x11617, x7156, x4741);
  nand n11618(x11618, x11617, x11616);
  nand n11619(x11619, x2269, x4611);
  nand n11620(x11620, x7156, x4481);
  nand n11621(x11621, x11620, x11619);
  nand n11622(x11622, x2272, x11612);
  nand n11623(x11623, x7169, x11615);
  nand n11624(x11624, x11623, x11622);
  nand n11625(x11625, x2272, x11618);
  nand n11626(x11626, x7169, x11621);
  nand n11627(x11627, x11626, x11625);
  nand n11628(x11628, x2275, x11624);
  nand n11629(x11629, x7176, x11627);
  nand n11630(x11630, x11629, x11628);
  nand n11631(x11631, x2269, x5395);
  nand n11632(x11632, x7156, x5265);
  nand n11633(x11633, x11632, x11631);
  nand n11634(x11634, x2269, x5135);
  nand n11635(x11635, x7156, x5005);
  nand n11636(x11636, x11635, x11634);
  nand n11637(x11637, x2269, x4875);
  nand n11638(x11638, x7156, x4745);
  nand n11639(x11639, x11638, x11637);
  nand n11640(x11640, x2269, x4615);
  nand n11641(x11641, x7156, x4485);
  nand n11642(x11642, x11641, x11640);
  nand n11643(x11643, x2272, x11633);
  nand n11644(x11644, x7169, x11636);
  nand n11645(x11645, x11644, x11643);
  nand n11646(x11646, x2272, x11639);
  nand n11647(x11647, x7169, x11642);
  nand n11648(x11648, x11647, x11646);
  nand n11649(x11649, x2275, x11645);
  nand n11650(x11650, x7176, x11648);
  nand n11651(x11651, x11650, x11649);
  nand n11652(x11652, x2269, x5399);
  nand n11653(x11653, x7156, x5269);
  nand n11654(x11654, x11653, x11652);
  nand n11655(x11655, x2269, x5139);
  nand n11656(x11656, x7156, x5009);
  nand n11657(x11657, x11656, x11655);
  nand n11658(x11658, x2269, x4879);
  nand n11659(x11659, x7156, x4749);
  nand n11660(x11660, x11659, x11658);
  nand n11661(x11661, x2269, x4619);
  nand n11662(x11662, x7156, x4489);
  nand n11663(x11663, x11662, x11661);
  nand n11664(x11664, x2272, x11654);
  nand n11665(x11665, x7169, x11657);
  nand n11666(x11666, x11665, x11664);
  nand n11667(x11667, x2272, x11660);
  nand n11668(x11668, x7169, x11663);
  nand n11669(x11669, x11668, x11667);
  nand n11670(x11670, x2275, x11666);
  nand n11671(x11671, x7176, x11669);
  nand n11672(x11672, x11671, x11670);
  nand n11673(x11673, x2269, x5403);
  nand n11674(x11674, x7156, x5273);
  nand n11675(x11675, x11674, x11673);
  nand n11676(x11676, x2269, x5143);
  nand n11677(x11677, x7156, x5013);
  nand n11678(x11678, x11677, x11676);
  nand n11679(x11679, x2269, x4883);
  nand n11680(x11680, x7156, x4753);
  nand n11681(x11681, x11680, x11679);
  nand n11682(x11682, x2269, x4623);
  nand n11683(x11683, x7156, x4493);
  nand n11684(x11684, x11683, x11682);
  nand n11685(x11685, x2272, x11675);
  nand n11686(x11686, x7169, x11678);
  nand n11687(x11687, x11686, x11685);
  nand n11688(x11688, x2272, x11681);
  nand n11689(x11689, x7169, x11684);
  nand n11690(x11690, x11689, x11688);
  nand n11691(x11691, x2275, x11687);
  nand n11692(x11692, x7176, x11690);
  nand n11693(x11693, x11692, x11691);
  nand n11694(x11694, x2269, x5407);
  nand n11695(x11695, x7156, x5277);
  nand n11696(x11696, x11695, x11694);
  nand n11697(x11697, x2269, x5147);
  nand n11698(x11698, x7156, x5017);
  nand n11699(x11699, x11698, x11697);
  nand n11700(x11700, x2269, x4887);
  nand n11701(x11701, x7156, x4757);
  nand n11702(x11702, x11701, x11700);
  nand n11703(x11703, x2269, x4627);
  nand n11704(x11704, x7156, x4497);
  nand n11705(x11705, x11704, x11703);
  nand n11706(x11706, x2272, x11696);
  nand n11707(x11707, x7169, x11699);
  nand n11708(x11708, x11707, x11706);
  nand n11709(x11709, x2272, x11702);
  nand n11710(x11710, x7169, x11705);
  nand n11711(x11711, x11710, x11709);
  nand n11712(x11712, x2275, x11708);
  nand n11713(x11713, x7176, x11711);
  nand n11714(x11714, x11713, x11712);
  nand n11715(x11715, x2269, x5411);
  nand n11716(x11716, x7156, x5281);
  nand n11717(x11717, x11716, x11715);
  nand n11718(x11718, x2269, x5151);
  nand n11719(x11719, x7156, x5021);
  nand n11720(x11720, x11719, x11718);
  nand n11721(x11721, x2269, x4891);
  nand n11722(x11722, x7156, x4761);
  nand n11723(x11723, x11722, x11721);
  nand n11724(x11724, x2269, x4631);
  nand n11725(x11725, x7156, x4501);
  nand n11726(x11726, x11725, x11724);
  nand n11727(x11727, x2272, x11717);
  nand n11728(x11728, x7169, x11720);
  nand n11729(x11729, x11728, x11727);
  nand n11730(x11730, x2272, x11723);
  nand n11731(x11731, x7169, x11726);
  nand n11732(x11732, x11731, x11730);
  nand n11733(x11733, x2275, x11729);
  nand n11734(x11734, x7176, x11732);
  nand n11735(x11735, x11734, x11733);
  nand n11736(x11736, x2269, x5415);
  nand n11737(x11737, x7156, x5285);
  nand n11738(x11738, x11737, x11736);
  nand n11739(x11739, x2269, x5155);
  nand n11740(x11740, x7156, x5025);
  nand n11741(x11741, x11740, x11739);
  nand n11742(x11742, x2269, x4895);
  nand n11743(x11743, x7156, x4765);
  nand n11744(x11744, x11743, x11742);
  nand n11745(x11745, x2269, x4635);
  nand n11746(x11746, x7156, x4505);
  nand n11747(x11747, x11746, x11745);
  nand n11748(x11748, x2272, x11738);
  nand n11749(x11749, x7169, x11741);
  nand n11750(x11750, x11749, x11748);
  nand n11751(x11751, x2272, x11744);
  nand n11752(x11752, x7169, x11747);
  nand n11753(x11753, x11752, x11751);
  nand n11754(x11754, x2275, x11750);
  nand n11755(x11755, x7176, x11753);
  nand n11756(x11756, x11755, x11754);
  nand n11757(x11757, x2269, x5419);
  nand n11758(x11758, x7156, x5289);
  nand n11759(x11759, x11758, x11757);
  nand n11760(x11760, x2269, x5159);
  nand n11761(x11761, x7156, x5029);
  nand n11762(x11762, x11761, x11760);
  nand n11763(x11763, x2269, x4899);
  nand n11764(x11764, x7156, x4769);
  nand n11765(x11765, x11764, x11763);
  nand n11766(x11766, x2269, x4639);
  nand n11767(x11767, x7156, x4509);
  nand n11768(x11768, x11767, x11766);
  nand n11769(x11769, x2272, x11759);
  nand n11770(x11770, x7169, x11762);
  nand n11771(x11771, x11770, x11769);
  nand n11772(x11772, x2272, x11765);
  nand n11773(x11773, x7169, x11768);
  nand n11774(x11774, x11773, x11772);
  nand n11775(x11775, x2275, x11771);
  nand n11776(x11776, x7176, x11774);
  nand n11777(x11777, x11776, x11775);
  nand n11778(x11778, x2269, x5423);
  nand n11779(x11779, x7156, x5293);
  nand n11780(x11780, x11779, x11778);
  nand n11781(x11781, x2269, x5163);
  nand n11782(x11782, x7156, x5033);
  nand n11783(x11783, x11782, x11781);
  nand n11784(x11784, x2269, x4903);
  nand n11785(x11785, x7156, x4773);
  nand n11786(x11786, x11785, x11784);
  nand n11787(x11787, x2269, x4643);
  nand n11788(x11788, x7156, x4513);
  nand n11789(x11789, x11788, x11787);
  nand n11790(x11790, x2272, x11780);
  nand n11791(x11791, x7169, x11783);
  nand n11792(x11792, x11791, x11790);
  nand n11793(x11793, x2272, x11786);
  nand n11794(x11794, x7169, x11789);
  nand n11795(x11795, x11794, x11793);
  nand n11796(x11796, x2275, x11792);
  nand n11797(x11797, x7176, x11795);
  nand n11798(x11798, x11797, x11796);
  nand n11799(x11799, x2269, x5427);
  nand n11800(x11800, x7156, x5297);
  nand n11801(x11801, x11800, x11799);
  nand n11802(x11802, x2269, x5167);
  nand n11803(x11803, x7156, x5037);
  nand n11804(x11804, x11803, x11802);
  nand n11805(x11805, x2269, x4907);
  nand n11806(x11806, x7156, x4777);
  nand n11807(x11807, x11806, x11805);
  nand n11808(x11808, x2269, x4647);
  nand n11809(x11809, x7156, x4517);
  nand n11810(x11810, x11809, x11808);
  nand n11811(x11811, x2272, x11801);
  nand n11812(x11812, x7169, x11804);
  nand n11813(x11813, x11812, x11811);
  nand n11814(x11814, x2272, x11807);
  nand n11815(x11815, x7169, x11810);
  nand n11816(x11816, x11815, x11814);
  nand n11817(x11817, x2275, x11813);
  nand n11818(x11818, x7176, x11816);
  nand n11819(x11819, x11818, x11817);
  nand n11820(x11820, x2269, x5431);
  nand n11821(x11821, x7156, x5301);
  nand n11822(x11822, x11821, x11820);
  nand n11823(x11823, x2269, x5171);
  nand n11824(x11824, x7156, x5041);
  nand n11825(x11825, x11824, x11823);
  nand n11826(x11826, x2269, x4911);
  nand n11827(x11827, x7156, x4781);
  nand n11828(x11828, x11827, x11826);
  nand n11829(x11829, x2269, x4651);
  nand n11830(x11830, x7156, x4521);
  nand n11831(x11831, x11830, x11829);
  nand n11832(x11832, x2272, x11822);
  nand n11833(x11833, x7169, x11825);
  nand n11834(x11834, x11833, x11832);
  nand n11835(x11835, x2272, x11828);
  nand n11836(x11836, x7169, x11831);
  nand n11837(x11837, x11836, x11835);
  nand n11838(x11838, x2275, x11834);
  nand n11839(x11839, x7176, x11837);
  nand n11840(x11840, x11839, x11838);
  nand n11841(x11841, x2269, x5435);
  nand n11842(x11842, x7156, x5305);
  nand n11843(x11843, x11842, x11841);
  nand n11844(x11844, x2269, x5175);
  nand n11845(x11845, x7156, x5045);
  nand n11846(x11846, x11845, x11844);
  nand n11847(x11847, x2269, x4915);
  nand n11848(x11848, x7156, x4785);
  nand n11849(x11849, x11848, x11847);
  nand n11850(x11850, x2269, x4655);
  nand n11851(x11851, x7156, x4525);
  nand n11852(x11852, x11851, x11850);
  nand n11853(x11853, x2272, x11843);
  nand n11854(x11854, x7169, x11846);
  nand n11855(x11855, x11854, x11853);
  nand n11856(x11856, x2272, x11849);
  nand n11857(x11857, x7169, x11852);
  nand n11858(x11858, x11857, x11856);
  nand n11859(x11859, x2275, x11855);
  nand n11860(x11860, x7176, x11858);
  nand n11861(x11861, x11860, x11859);
  nand n11862(x11862, x71202, x5311);
  nand n11863(x11863, x1448, x5181);
  nand n11864(x11864, x11863, x11862);
  nand n11865(x11865, x71202, x5051);
  nand n11866(x11866, x1448, x4921);
  nand n11867(x11867, x11866, x11865);
  nand n11868(x11868, x71202, x4791);
  nand n11869(x11869, x1448, x4661);
  nand n11870(x11870, x11869, x11868);
  nand n11871(x11871, x71202, x4531);
  nand n11872(x11872, x1448, x4399);
  nand n11873(x11873, x11872, x11871);
  nand n11874(x11874, x71205, x11864);
  nand n11875(x11875, x1461, x11867);
  nand n11876(x11876, x11875, x11874);
  nand n11877(x11877, x71205, x11870);
  nand n11878(x11878, x1461, x11873);
  nand n11879(x11879, x11878, x11877);
  nand n11880(x11880, x71210, x11876);
  nand n11881(x11881, x1468, x11879);
  nand n11882(x11882, x11881, x11880);
  nand n11883(x11883, x71202, x5315);
  nand n11884(x11884, x1448, x5185);
  nand n11885(x11885, x11884, x11883);
  nand n11886(x11886, x71202, x5055);
  nand n11887(x11887, x1448, x4925);
  nand n11888(x11888, x11887, x11886);
  nand n11889(x11889, x71202, x4795);
  nand n11890(x11890, x1448, x4665);
  nand n11891(x11891, x11890, x11889);
  nand n11892(x11892, x71202, x4535);
  nand n11893(x11893, x1448, x4405);
  nand n11894(x11894, x11893, x11892);
  nand n11895(x11895, x71205, x11885);
  nand n11896(x11896, x1461, x11888);
  nand n11897(x11897, x11896, x11895);
  nand n11898(x11898, x71205, x11891);
  nand n11899(x11899, x1461, x11894);
  nand n11900(x11900, x11899, x11898);
  nand n11901(x11901, x71210, x11897);
  nand n11902(x11902, x1468, x11900);
  nand n11903(x11903, x11902, x11901);
  nand n11904(x11904, x71202, x5319);
  nand n11905(x11905, x1448, x5189);
  nand n11906(x11906, x11905, x11904);
  nand n11907(x11907, x71202, x5059);
  nand n11908(x11908, x1448, x4929);
  nand n11909(x11909, x11908, x11907);
  nand n11910(x11910, x71202, x4799);
  nand n11911(x11911, x1448, x4669);
  nand n11912(x11912, x11911, x11910);
  nand n11913(x11913, x71202, x4539);
  nand n11914(x11914, x1448, x4409);
  nand n11915(x11915, x11914, x11913);
  nand n11916(x11916, x71205, x11906);
  nand n11917(x11917, x1461, x11909);
  nand n11918(x11918, x11917, x11916);
  nand n11919(x11919, x71205, x11912);
  nand n11920(x11920, x1461, x11915);
  nand n11921(x11921, x11920, x11919);
  nand n11922(x11922, x71210, x11918);
  nand n11923(x11923, x1468, x11921);
  nand n11924(x11924, x11923, x11922);
  nand n11925(x11925, x71202, x5323);
  nand n11926(x11926, x1448, x5193);
  nand n11927(x11927, x11926, x11925);
  nand n11928(x11928, x71202, x5063);
  nand n11929(x11929, x1448, x4933);
  nand n11930(x11930, x11929, x11928);
  nand n11931(x11931, x71202, x4803);
  nand n11932(x11932, x1448, x4673);
  nand n11933(x11933, x11932, x11931);
  nand n11934(x11934, x71202, x4543);
  nand n11935(x11935, x1448, x4413);
  nand n11936(x11936, x11935, x11934);
  nand n11937(x11937, x71205, x11927);
  nand n11938(x11938, x1461, x11930);
  nand n11939(x11939, x11938, x11937);
  nand n11940(x11940, x71205, x11933);
  nand n11941(x11941, x1461, x11936);
  nand n11942(x11942, x11941, x11940);
  nand n11943(x11943, x71210, x11939);
  nand n11944(x11944, x1468, x11942);
  nand n11945(x11945, x11944, x11943);
  nand n11946(x11946, x71202, x5327);
  nand n11947(x11947, x1448, x5197);
  nand n11948(x11948, x11947, x11946);
  nand n11949(x11949, x71202, x5067);
  nand n11950(x11950, x1448, x4937);
  nand n11951(x11951, x11950, x11949);
  nand n11952(x11952, x71202, x4807);
  nand n11953(x11953, x1448, x4677);
  nand n11954(x11954, x11953, x11952);
  nand n11955(x11955, x71202, x4547);
  nand n11956(x11956, x1448, x4417);
  nand n11957(x11957, x11956, x11955);
  nand n11958(x11958, x71205, x11948);
  nand n11959(x11959, x1461, x11951);
  nand n11960(x11960, x11959, x11958);
  nand n11961(x11961, x71205, x11954);
  nand n11962(x11962, x1461, x11957);
  nand n11963(x11963, x11962, x11961);
  nand n11964(x11964, x71210, x11960);
  nand n11965(x11965, x1468, x11963);
  nand n11966(x11966, x11965, x11964);
  nand n11967(x11967, x71202, x5331);
  nand n11968(x11968, x1448, x5201);
  nand n11969(x11969, x11968, x11967);
  nand n11970(x11970, x71202, x5071);
  nand n11971(x11971, x1448, x4941);
  nand n11972(x11972, x11971, x11970);
  nand n11973(x11973, x71202, x4811);
  nand n11974(x11974, x1448, x4681);
  nand n11975(x11975, x11974, x11973);
  nand n11976(x11976, x71202, x4551);
  nand n11977(x11977, x1448, x4421);
  nand n11978(x11978, x11977, x11976);
  nand n11979(x11979, x71205, x11969);
  nand n11980(x11980, x1461, x11972);
  nand n11981(x11981, x11980, x11979);
  nand n11982(x11982, x71205, x11975);
  nand n11983(x11983, x1461, x11978);
  nand n11984(x11984, x11983, x11982);
  nand n11985(x11985, x71210, x11981);
  nand n11986(x11986, x1468, x11984);
  nand n11987(x11987, x11986, x11985);
  nand n11988(x11988, x71202, x5335);
  nand n11989(x11989, x1448, x5205);
  nand n11990(x11990, x11989, x11988);
  nand n11991(x11991, x71202, x5075);
  nand n11992(x11992, x1448, x4945);
  nand n11993(x11993, x11992, x11991);
  nand n11994(x11994, x71202, x4815);
  nand n11995(x11995, x1448, x4685);
  nand n11996(x11996, x11995, x11994);
  nand n11997(x11997, x71202, x4555);
  nand n11998(x11998, x1448, x4425);
  nand n11999(x11999, x11998, x11997);
  nand n12000(x12000, x71205, x11990);
  nand n12001(x12001, x1461, x11993);
  nand n12002(x12002, x12001, x12000);
  nand n12003(x12003, x71205, x11996);
  nand n12004(x12004, x1461, x11999);
  nand n12005(x12005, x12004, x12003);
  nand n12006(x12006, x71210, x12002);
  nand n12007(x12007, x1468, x12005);
  nand n12008(x12008, x12007, x12006);
  nand n12009(x12009, x71202, x5339);
  nand n12010(x12010, x1448, x5209);
  nand n12011(x12011, x12010, x12009);
  nand n12012(x12012, x71202, x5079);
  nand n12013(x12013, x1448, x4949);
  nand n12014(x12014, x12013, x12012);
  nand n12015(x12015, x71202, x4819);
  nand n12016(x12016, x1448, x4689);
  nand n12017(x12017, x12016, x12015);
  nand n12018(x12018, x71202, x4559);
  nand n12019(x12019, x1448, x4429);
  nand n12020(x12020, x12019, x12018);
  nand n12021(x12021, x71205, x12011);
  nand n12022(x12022, x1461, x12014);
  nand n12023(x12023, x12022, x12021);
  nand n12024(x12024, x71205, x12017);
  nand n12025(x12025, x1461, x12020);
  nand n12026(x12026, x12025, x12024);
  nand n12027(x12027, x71210, x12023);
  nand n12028(x12028, x1468, x12026);
  nand n12029(x12029, x12028, x12027);
  nand n12030(x12030, x71202, x5343);
  nand n12031(x12031, x1448, x5213);
  nand n12032(x12032, x12031, x12030);
  nand n12033(x12033, x71202, x5083);
  nand n12034(x12034, x1448, x4953);
  nand n12035(x12035, x12034, x12033);
  nand n12036(x12036, x71202, x4823);
  nand n12037(x12037, x1448, x4693);
  nand n12038(x12038, x12037, x12036);
  nand n12039(x12039, x71202, x4563);
  nand n12040(x12040, x1448, x4433);
  nand n12041(x12041, x12040, x12039);
  nand n12042(x12042, x71205, x12032);
  nand n12043(x12043, x1461, x12035);
  nand n12044(x12044, x12043, x12042);
  nand n12045(x12045, x71205, x12038);
  nand n12046(x12046, x1461, x12041);
  nand n12047(x12047, x12046, x12045);
  nand n12048(x12048, x71210, x12044);
  nand n12049(x12049, x1468, x12047);
  nand n12050(x12050, x12049, x12048);
  nand n12051(x12051, x71202, x5347);
  nand n12052(x12052, x1448, x5217);
  nand n12053(x12053, x12052, x12051);
  nand n12054(x12054, x71202, x5087);
  nand n12055(x12055, x1448, x4957);
  nand n12056(x12056, x12055, x12054);
  nand n12057(x12057, x71202, x4827);
  nand n12058(x12058, x1448, x4697);
  nand n12059(x12059, x12058, x12057);
  nand n12060(x12060, x71202, x4567);
  nand n12061(x12061, x1448, x4437);
  nand n12062(x12062, x12061, x12060);
  nand n12063(x12063, x71205, x12053);
  nand n12064(x12064, x1461, x12056);
  nand n12065(x12065, x12064, x12063);
  nand n12066(x12066, x71205, x12059);
  nand n12067(x12067, x1461, x12062);
  nand n12068(x12068, x12067, x12066);
  nand n12069(x12069, x71210, x12065);
  nand n12070(x12070, x1468, x12068);
  nand n12071(x12071, x12070, x12069);
  nand n12072(x12072, x71202, x5351);
  nand n12073(x12073, x1448, x5221);
  nand n12074(x12074, x12073, x12072);
  nand n12075(x12075, x71202, x5091);
  nand n12076(x12076, x1448, x4961);
  nand n12077(x12077, x12076, x12075);
  nand n12078(x12078, x71202, x4831);
  nand n12079(x12079, x1448, x4701);
  nand n12080(x12080, x12079, x12078);
  nand n12081(x12081, x71202, x4571);
  nand n12082(x12082, x1448, x4441);
  nand n12083(x12083, x12082, x12081);
  nand n12084(x12084, x71205, x12074);
  nand n12085(x12085, x1461, x12077);
  nand n12086(x12086, x12085, x12084);
  nand n12087(x12087, x71205, x12080);
  nand n12088(x12088, x1461, x12083);
  nand n12089(x12089, x12088, x12087);
  nand n12090(x12090, x71210, x12086);
  nand n12091(x12091, x1468, x12089);
  nand n12092(x12092, x12091, x12090);
  nand n12093(x12093, x71202, x5355);
  nand n12094(x12094, x1448, x5225);
  nand n12095(x12095, x12094, x12093);
  nand n12096(x12096, x71202, x5095);
  nand n12097(x12097, x1448, x4965);
  nand n12098(x12098, x12097, x12096);
  nand n12099(x12099, x71202, x4835);
  nand n12100(x12100, x1448, x4705);
  nand n12101(x12101, x12100, x12099);
  nand n12102(x12102, x71202, x4575);
  nand n12103(x12103, x1448, x4445);
  nand n12104(x12104, x12103, x12102);
  nand n12105(x12105, x71205, x12095);
  nand n12106(x12106, x1461, x12098);
  nand n12107(x12107, x12106, x12105);
  nand n12108(x12108, x71205, x12101);
  nand n12109(x12109, x1461, x12104);
  nand n12110(x12110, x12109, x12108);
  nand n12111(x12111, x71210, x12107);
  nand n12112(x12112, x1468, x12110);
  nand n12113(x12113, x12112, x12111);
  nand n12114(x12114, x71202, x5359);
  nand n12115(x12115, x1448, x5229);
  nand n12116(x12116, x12115, x12114);
  nand n12117(x12117, x71202, x5099);
  nand n12118(x12118, x1448, x4969);
  nand n12119(x12119, x12118, x12117);
  nand n12120(x12120, x71202, x4839);
  nand n12121(x12121, x1448, x4709);
  nand n12122(x12122, x12121, x12120);
  nand n12123(x12123, x71202, x4579);
  nand n12124(x12124, x1448, x4449);
  nand n12125(x12125, x12124, x12123);
  nand n12126(x12126, x71205, x12116);
  nand n12127(x12127, x1461, x12119);
  nand n12128(x12128, x12127, x12126);
  nand n12129(x12129, x71205, x12122);
  nand n12130(x12130, x1461, x12125);
  nand n12131(x12131, x12130, x12129);
  nand n12132(x12132, x71210, x12128);
  nand n12133(x12133, x1468, x12131);
  nand n12134(x12134, x12133, x12132);
  nand n12135(x12135, x71202, x5363);
  nand n12136(x12136, x1448, x5233);
  nand n12137(x12137, x12136, x12135);
  nand n12138(x12138, x71202, x5103);
  nand n12139(x12139, x1448, x4973);
  nand n12140(x12140, x12139, x12138);
  nand n12141(x12141, x71202, x4843);
  nand n12142(x12142, x1448, x4713);
  nand n12143(x12143, x12142, x12141);
  nand n12144(x12144, x71202, x4583);
  nand n12145(x12145, x1448, x4453);
  nand n12146(x12146, x12145, x12144);
  nand n12147(x12147, x71205, x12137);
  nand n12148(x12148, x1461, x12140);
  nand n12149(x12149, x12148, x12147);
  nand n12150(x12150, x71205, x12143);
  nand n12151(x12151, x1461, x12146);
  nand n12152(x12152, x12151, x12150);
  nand n12153(x12153, x71210, x12149);
  nand n12154(x12154, x1468, x12152);
  nand n12155(x12155, x12154, x12153);
  nand n12156(x12156, x71202, x5367);
  nand n12157(x12157, x1448, x5237);
  nand n12158(x12158, x12157, x12156);
  nand n12159(x12159, x71202, x5107);
  nand n12160(x12160, x1448, x4977);
  nand n12161(x12161, x12160, x12159);
  nand n12162(x12162, x71202, x4847);
  nand n12163(x12163, x1448, x4717);
  nand n12164(x12164, x12163, x12162);
  nand n12165(x12165, x71202, x4587);
  nand n12166(x12166, x1448, x4457);
  nand n12167(x12167, x12166, x12165);
  nand n12168(x12168, x71205, x12158);
  nand n12169(x12169, x1461, x12161);
  nand n12170(x12170, x12169, x12168);
  nand n12171(x12171, x71205, x12164);
  nand n12172(x12172, x1461, x12167);
  nand n12173(x12173, x12172, x12171);
  nand n12174(x12174, x71210, x12170);
  nand n12175(x12175, x1468, x12173);
  nand n12176(x12176, x12175, x12174);
  nand n12177(x12177, x71202, x5371);
  nand n12178(x12178, x1448, x5241);
  nand n12179(x12179, x12178, x12177);
  nand n12180(x12180, x71202, x5111);
  nand n12181(x12181, x1448, x4981);
  nand n12182(x12182, x12181, x12180);
  nand n12183(x12183, x71202, x4851);
  nand n12184(x12184, x1448, x4721);
  nand n12185(x12185, x12184, x12183);
  nand n12186(x12186, x71202, x4591);
  nand n12187(x12187, x1448, x4461);
  nand n12188(x12188, x12187, x12186);
  nand n12189(x12189, x71205, x12179);
  nand n12190(x12190, x1461, x12182);
  nand n12191(x12191, x12190, x12189);
  nand n12192(x12192, x71205, x12185);
  nand n12193(x12193, x1461, x12188);
  nand n12194(x12194, x12193, x12192);
  nand n12195(x12195, x71210, x12191);
  nand n12196(x12196, x1468, x12194);
  nand n12197(x12197, x12196, x12195);
  nand n12198(x12198, x71202, x5375);
  nand n12199(x12199, x1448, x5245);
  nand n12200(x12200, x12199, x12198);
  nand n12201(x12201, x71202, x5115);
  nand n12202(x12202, x1448, x4985);
  nand n12203(x12203, x12202, x12201);
  nand n12204(x12204, x71202, x4855);
  nand n12205(x12205, x1448, x4725);
  nand n12206(x12206, x12205, x12204);
  nand n12207(x12207, x71202, x4595);
  nand n12208(x12208, x1448, x4465);
  nand n12209(x12209, x12208, x12207);
  nand n12210(x12210, x71205, x12200);
  nand n12211(x12211, x1461, x12203);
  nand n12212(x12212, x12211, x12210);
  nand n12213(x12213, x71205, x12206);
  nand n12214(x12214, x1461, x12209);
  nand n12215(x12215, x12214, x12213);
  nand n12216(x12216, x71210, x12212);
  nand n12217(x12217, x1468, x12215);
  nand n12218(x12218, x12217, x12216);
  nand n12219(x12219, x71202, x5379);
  nand n12220(x12220, x1448, x5249);
  nand n12221(x12221, x12220, x12219);
  nand n12222(x12222, x71202, x5119);
  nand n12223(x12223, x1448, x4989);
  nand n12224(x12224, x12223, x12222);
  nand n12225(x12225, x71202, x4859);
  nand n12226(x12226, x1448, x4729);
  nand n12227(x12227, x12226, x12225);
  nand n12228(x12228, x71202, x4599);
  nand n12229(x12229, x1448, x4469);
  nand n12230(x12230, x12229, x12228);
  nand n12231(x12231, x71205, x12221);
  nand n12232(x12232, x1461, x12224);
  nand n12233(x12233, x12232, x12231);
  nand n12234(x12234, x71205, x12227);
  nand n12235(x12235, x1461, x12230);
  nand n12236(x12236, x12235, x12234);
  nand n12237(x12237, x71210, x12233);
  nand n12238(x12238, x1468, x12236);
  nand n12239(x12239, x12238, x12237);
  nand n12240(x12240, x71202, x5383);
  nand n12241(x12241, x1448, x5253);
  nand n12242(x12242, x12241, x12240);
  nand n12243(x12243, x71202, x5123);
  nand n12244(x12244, x1448, x4993);
  nand n12245(x12245, x12244, x12243);
  nand n12246(x12246, x71202, x4863);
  nand n12247(x12247, x1448, x4733);
  nand n12248(x12248, x12247, x12246);
  nand n12249(x12249, x71202, x4603);
  nand n12250(x12250, x1448, x4473);
  nand n12251(x12251, x12250, x12249);
  nand n12252(x12252, x71205, x12242);
  nand n12253(x12253, x1461, x12245);
  nand n12254(x12254, x12253, x12252);
  nand n12255(x12255, x71205, x12248);
  nand n12256(x12256, x1461, x12251);
  nand n12257(x12257, x12256, x12255);
  nand n12258(x12258, x71210, x12254);
  nand n12259(x12259, x1468, x12257);
  nand n12260(x12260, x12259, x12258);
  nand n12261(x12261, x71202, x5387);
  nand n12262(x12262, x1448, x5257);
  nand n12263(x12263, x12262, x12261);
  nand n12264(x12264, x71202, x5127);
  nand n12265(x12265, x1448, x4997);
  nand n12266(x12266, x12265, x12264);
  nand n12267(x12267, x71202, x4867);
  nand n12268(x12268, x1448, x4737);
  nand n12269(x12269, x12268, x12267);
  nand n12270(x12270, x71202, x4607);
  nand n12271(x12271, x1448, x4477);
  nand n12272(x12272, x12271, x12270);
  nand n12273(x12273, x71205, x12263);
  nand n12274(x12274, x1461, x12266);
  nand n12275(x12275, x12274, x12273);
  nand n12276(x12276, x71205, x12269);
  nand n12277(x12277, x1461, x12272);
  nand n12278(x12278, x12277, x12276);
  nand n12279(x12279, x71210, x12275);
  nand n12280(x12280, x1468, x12278);
  nand n12281(x12281, x12280, x12279);
  nand n12282(x12282, x71202, x5391);
  nand n12283(x12283, x1448, x5261);
  nand n12284(x12284, x12283, x12282);
  nand n12285(x12285, x71202, x5131);
  nand n12286(x12286, x1448, x5001);
  nand n12287(x12287, x12286, x12285);
  nand n12288(x12288, x71202, x4871);
  nand n12289(x12289, x1448, x4741);
  nand n12290(x12290, x12289, x12288);
  nand n12291(x12291, x71202, x4611);
  nand n12292(x12292, x1448, x4481);
  nand n12293(x12293, x12292, x12291);
  nand n12294(x12294, x71205, x12284);
  nand n12295(x12295, x1461, x12287);
  nand n12296(x12296, x12295, x12294);
  nand n12297(x12297, x71205, x12290);
  nand n12298(x12298, x1461, x12293);
  nand n12299(x12299, x12298, x12297);
  nand n12300(x12300, x71210, x12296);
  nand n12301(x12301, x1468, x12299);
  nand n12302(x12302, x12301, x12300);
  nand n12303(x12303, x71202, x5395);
  nand n12304(x12304, x1448, x5265);
  nand n12305(x12305, x12304, x12303);
  nand n12306(x12306, x71202, x5135);
  nand n12307(x12307, x1448, x5005);
  nand n12308(x12308, x12307, x12306);
  nand n12309(x12309, x71202, x4875);
  nand n12310(x12310, x1448, x4745);
  nand n12311(x12311, x12310, x12309);
  nand n12312(x12312, x71202, x4615);
  nand n12313(x12313, x1448, x4485);
  nand n12314(x12314, x12313, x12312);
  nand n12315(x12315, x71205, x12305);
  nand n12316(x12316, x1461, x12308);
  nand n12317(x12317, x12316, x12315);
  nand n12318(x12318, x71205, x12311);
  nand n12319(x12319, x1461, x12314);
  nand n12320(x12320, x12319, x12318);
  nand n12321(x12321, x71210, x12317);
  nand n12322(x12322, x1468, x12320);
  nand n12323(x12323, x12322, x12321);
  nand n12324(x12324, x71202, x5399);
  nand n12325(x12325, x1448, x5269);
  nand n12326(x12326, x12325, x12324);
  nand n12327(x12327, x71202, x5139);
  nand n12328(x12328, x1448, x5009);
  nand n12329(x12329, x12328, x12327);
  nand n12330(x12330, x71202, x4879);
  nand n12331(x12331, x1448, x4749);
  nand n12332(x12332, x12331, x12330);
  nand n12333(x12333, x71202, x4619);
  nand n12334(x12334, x1448, x4489);
  nand n12335(x12335, x12334, x12333);
  nand n12336(x12336, x71205, x12326);
  nand n12337(x12337, x1461, x12329);
  nand n12338(x12338, x12337, x12336);
  nand n12339(x12339, x71205, x12332);
  nand n12340(x12340, x1461, x12335);
  nand n12341(x12341, x12340, x12339);
  nand n12342(x12342, x71210, x12338);
  nand n12343(x12343, x1468, x12341);
  nand n12344(x12344, x12343, x12342);
  nand n12345(x12345, x71202, x5403);
  nand n12346(x12346, x1448, x5273);
  nand n12347(x12347, x12346, x12345);
  nand n12348(x12348, x71202, x5143);
  nand n12349(x12349, x1448, x5013);
  nand n12350(x12350, x12349, x12348);
  nand n12351(x12351, x71202, x4883);
  nand n12352(x12352, x1448, x4753);
  nand n12353(x12353, x12352, x12351);
  nand n12354(x12354, x71202, x4623);
  nand n12355(x12355, x1448, x4493);
  nand n12356(x12356, x12355, x12354);
  nand n12357(x12357, x71205, x12347);
  nand n12358(x12358, x1461, x12350);
  nand n12359(x12359, x12358, x12357);
  nand n12360(x12360, x71205, x12353);
  nand n12361(x12361, x1461, x12356);
  nand n12362(x12362, x12361, x12360);
  nand n12363(x12363, x71210, x12359);
  nand n12364(x12364, x1468, x12362);
  nand n12365(x12365, x12364, x12363);
  nand n12366(x12366, x71202, x5407);
  nand n12367(x12367, x1448, x5277);
  nand n12368(x12368, x12367, x12366);
  nand n12369(x12369, x71202, x5147);
  nand n12370(x12370, x1448, x5017);
  nand n12371(x12371, x12370, x12369);
  nand n12372(x12372, x71202, x4887);
  nand n12373(x12373, x1448, x4757);
  nand n12374(x12374, x12373, x12372);
  nand n12375(x12375, x71202, x4627);
  nand n12376(x12376, x1448, x4497);
  nand n12377(x12377, x12376, x12375);
  nand n12378(x12378, x71205, x12368);
  nand n12379(x12379, x1461, x12371);
  nand n12380(x12380, x12379, x12378);
  nand n12381(x12381, x71205, x12374);
  nand n12382(x12382, x1461, x12377);
  nand n12383(x12383, x12382, x12381);
  nand n12384(x12384, x71210, x12380);
  nand n12385(x12385, x1468, x12383);
  nand n12386(x12386, x12385, x12384);
  nand n12387(x12387, x71202, x5411);
  nand n12388(x12388, x1448, x5281);
  nand n12389(x12389, x12388, x12387);
  nand n12390(x12390, x71202, x5151);
  nand n12391(x12391, x1448, x5021);
  nand n12392(x12392, x12391, x12390);
  nand n12393(x12393, x71202, x4891);
  nand n12394(x12394, x1448, x4761);
  nand n12395(x12395, x12394, x12393);
  nand n12396(x12396, x71202, x4631);
  nand n12397(x12397, x1448, x4501);
  nand n12398(x12398, x12397, x12396);
  nand n12399(x12399, x71205, x12389);
  nand n12400(x12400, x1461, x12392);
  nand n12401(x12401, x12400, x12399);
  nand n12402(x12402, x71205, x12395);
  nand n12403(x12403, x1461, x12398);
  nand n12404(x12404, x12403, x12402);
  nand n12405(x12405, x71210, x12401);
  nand n12406(x12406, x1468, x12404);
  nand n12407(x12407, x12406, x12405);
  nand n12408(x12408, x71202, x5415);
  nand n12409(x12409, x1448, x5285);
  nand n12410(x12410, x12409, x12408);
  nand n12411(x12411, x71202, x5155);
  nand n12412(x12412, x1448, x5025);
  nand n12413(x12413, x12412, x12411);
  nand n12414(x12414, x71202, x4895);
  nand n12415(x12415, x1448, x4765);
  nand n12416(x12416, x12415, x12414);
  nand n12417(x12417, x71202, x4635);
  nand n12418(x12418, x1448, x4505);
  nand n12419(x12419, x12418, x12417);
  nand n12420(x12420, x71205, x12410);
  nand n12421(x12421, x1461, x12413);
  nand n12422(x12422, x12421, x12420);
  nand n12423(x12423, x71205, x12416);
  nand n12424(x12424, x1461, x12419);
  nand n12425(x12425, x12424, x12423);
  nand n12426(x12426, x71210, x12422);
  nand n12427(x12427, x1468, x12425);
  nand n12428(x12428, x12427, x12426);
  nand n12429(x12429, x71202, x5419);
  nand n12430(x12430, x1448, x5289);
  nand n12431(x12431, x12430, x12429);
  nand n12432(x12432, x71202, x5159);
  nand n12433(x12433, x1448, x5029);
  nand n12434(x12434, x12433, x12432);
  nand n12435(x12435, x71202, x4899);
  nand n12436(x12436, x1448, x4769);
  nand n12437(x12437, x12436, x12435);
  nand n12438(x12438, x71202, x4639);
  nand n12439(x12439, x1448, x4509);
  nand n12440(x12440, x12439, x12438);
  nand n12441(x12441, x71205, x12431);
  nand n12442(x12442, x1461, x12434);
  nand n12443(x12443, x12442, x12441);
  nand n12444(x12444, x71205, x12437);
  nand n12445(x12445, x1461, x12440);
  nand n12446(x12446, x12445, x12444);
  nand n12447(x12447, x71210, x12443);
  nand n12448(x12448, x1468, x12446);
  nand n12449(x12449, x12448, x12447);
  nand n12450(x12450, x71202, x5423);
  nand n12451(x12451, x1448, x5293);
  nand n12452(x12452, x12451, x12450);
  nand n12453(x12453, x71202, x5163);
  nand n12454(x12454, x1448, x5033);
  nand n12455(x12455, x12454, x12453);
  nand n12456(x12456, x71202, x4903);
  nand n12457(x12457, x1448, x4773);
  nand n12458(x12458, x12457, x12456);
  nand n12459(x12459, x71202, x4643);
  nand n12460(x12460, x1448, x4513);
  nand n12461(x12461, x12460, x12459);
  nand n12462(x12462, x71205, x12452);
  nand n12463(x12463, x1461, x12455);
  nand n12464(x12464, x12463, x12462);
  nand n12465(x12465, x71205, x12458);
  nand n12466(x12466, x1461, x12461);
  nand n12467(x12467, x12466, x12465);
  nand n12468(x12468, x71210, x12464);
  nand n12469(x12469, x1468, x12467);
  nand n12470(x12470, x12469, x12468);
  nand n12471(x12471, x71202, x5427);
  nand n12472(x12472, x1448, x5297);
  nand n12473(x12473, x12472, x12471);
  nand n12474(x12474, x71202, x5167);
  nand n12475(x12475, x1448, x5037);
  nand n12476(x12476, x12475, x12474);
  nand n12477(x12477, x71202, x4907);
  nand n12478(x12478, x1448, x4777);
  nand n12479(x12479, x12478, x12477);
  nand n12480(x12480, x71202, x4647);
  nand n12481(x12481, x1448, x4517);
  nand n12482(x12482, x12481, x12480);
  nand n12483(x12483, x71205, x12473);
  nand n12484(x12484, x1461, x12476);
  nand n12485(x12485, x12484, x12483);
  nand n12486(x12486, x71205, x12479);
  nand n12487(x12487, x1461, x12482);
  nand n12488(x12488, x12487, x12486);
  nand n12489(x12489, x71210, x12485);
  nand n12490(x12490, x1468, x12488);
  nand n12491(x12491, x12490, x12489);
  nand n12492(x12492, x71202, x5431);
  nand n12493(x12493, x1448, x5301);
  nand n12494(x12494, x12493, x12492);
  nand n12495(x12495, x71202, x5171);
  nand n12496(x12496, x1448, x5041);
  nand n12497(x12497, x12496, x12495);
  nand n12498(x12498, x71202, x4911);
  nand n12499(x12499, x1448, x4781);
  nand n12500(x12500, x12499, x12498);
  nand n12501(x12501, x71202, x4651);
  nand n12502(x12502, x1448, x4521);
  nand n12503(x12503, x12502, x12501);
  nand n12504(x12504, x71205, x12494);
  nand n12505(x12505, x1461, x12497);
  nand n12506(x12506, x12505, x12504);
  nand n12507(x12507, x71205, x12500);
  nand n12508(x12508, x1461, x12503);
  nand n12509(x12509, x12508, x12507);
  nand n12510(x12510, x71210, x12506);
  nand n12511(x12511, x1468, x12509);
  nand n12512(x12512, x12511, x12510);
  nand n12513(x12513, x71202, x5435);
  nand n12514(x12514, x1448, x5305);
  nand n12515(x12515, x12514, x12513);
  nand n12516(x12516, x71202, x5175);
  nand n12517(x12517, x1448, x5045);
  nand n12518(x12518, x12517, x12516);
  nand n12519(x12519, x71202, x4915);
  nand n12520(x12520, x1448, x4785);
  nand n12521(x12521, x12520, x12519);
  nand n12522(x12522, x71202, x4655);
  nand n12523(x12523, x1448, x4525);
  nand n12524(x12524, x12523, x12522);
  nand n12525(x12525, x71205, x12515);
  nand n12526(x12526, x1461, x12518);
  nand n12527(x12527, x12526, x12525);
  nand n12528(x12528, x71205, x12521);
  nand n12529(x12529, x1461, x12524);
  nand n12530(x12530, x12529, x12528);
  nand n12531(x12531, x71210, x12527);
  nand n12532(x12532, x1468, x12530);
  nand n12533(x12533, x12532, x12531);
  nand n12534(x12534, x2258, x6355);
  nand n12535(x12535, x6481, x6225);
  nand n12536(x12536, x12535, x12534);
  nand n12537(x12537, x2258, x6095);
  nand n12538(x12538, x6481, x5965);
  nand n12539(x12539, x12538, x12537);
  nand n12540(x12540, x2258, x5835);
  nand n12541(x12541, x6481, x5705);
  nand n12542(x12542, x12541, x12540);
  nand n12543(x12543, x2258, x5575);
  nand n12544(x12544, x6481, x5443);
  nand n12545(x12545, x12544, x12543);
  nand n12546(x12546, x2261, x12536);
  nand n12547(x12547, x6494, x12539);
  nand n12548(x12548, x12547, x12546);
  nand n12549(x12549, x2261, x12542);
  nand n12550(x12550, x6494, x12545);
  nand n12551(x12551, x12550, x12549);
  nand n12552(x12552, x2264, x12548);
  nand n12553(x12553, x6501, x12551);
  nand n12554(x12554, x12553, x12552);
  nand n12555(x12555, x2258, x6359);
  nand n12556(x12556, x6481, x6229);
  nand n12557(x12557, x12556, x12555);
  nand n12558(x12558, x2258, x6099);
  nand n12559(x12559, x6481, x5969);
  nand n12560(x12560, x12559, x12558);
  nand n12561(x12561, x2258, x5839);
  nand n12562(x12562, x6481, x5709);
  nand n12563(x12563, x12562, x12561);
  nand n12564(x12564, x2258, x5579);
  nand n12565(x12565, x6481, x5449);
  nand n12566(x12566, x12565, x12564);
  nand n12567(x12567, x2261, x12557);
  nand n12568(x12568, x6494, x12560);
  nand n12569(x12569, x12568, x12567);
  nand n12570(x12570, x2261, x12563);
  nand n12571(x12571, x6494, x12566);
  nand n12572(x12572, x12571, x12570);
  nand n12573(x12573, x2264, x12569);
  nand n12574(x12574, x6501, x12572);
  nand n12575(x12575, x12574, x12573);
  nand n12576(x12576, x2258, x6363);
  nand n12577(x12577, x6481, x6233);
  nand n12578(x12578, x12577, x12576);
  nand n12579(x12579, x2258, x6103);
  nand n12580(x12580, x6481, x5973);
  nand n12581(x12581, x12580, x12579);
  nand n12582(x12582, x2258, x5843);
  nand n12583(x12583, x6481, x5713);
  nand n12584(x12584, x12583, x12582);
  nand n12585(x12585, x2258, x5583);
  nand n12586(x12586, x6481, x5453);
  nand n12587(x12587, x12586, x12585);
  nand n12588(x12588, x2261, x12578);
  nand n12589(x12589, x6494, x12581);
  nand n12590(x12590, x12589, x12588);
  nand n12591(x12591, x2261, x12584);
  nand n12592(x12592, x6494, x12587);
  nand n12593(x12593, x12592, x12591);
  nand n12594(x12594, x2264, x12590);
  nand n12595(x12595, x6501, x12593);
  nand n12596(x12596, x12595, x12594);
  nand n12597(x12597, x2258, x6367);
  nand n12598(x12598, x6481, x6237);
  nand n12599(x12599, x12598, x12597);
  nand n12600(x12600, x2258, x6107);
  nand n12601(x12601, x6481, x5977);
  nand n12602(x12602, x12601, x12600);
  nand n12603(x12603, x2258, x5847);
  nand n12604(x12604, x6481, x5717);
  nand n12605(x12605, x12604, x12603);
  nand n12606(x12606, x2258, x5587);
  nand n12607(x12607, x6481, x5457);
  nand n12608(x12608, x12607, x12606);
  nand n12609(x12609, x2261, x12599);
  nand n12610(x12610, x6494, x12602);
  nand n12611(x12611, x12610, x12609);
  nand n12612(x12612, x2261, x12605);
  nand n12613(x12613, x6494, x12608);
  nand n12614(x12614, x12613, x12612);
  nand n12615(x12615, x2264, x12611);
  nand n12616(x12616, x6501, x12614);
  nand n12617(x12617, x12616, x12615);
  nand n12618(x12618, x2258, x6371);
  nand n12619(x12619, x6481, x6241);
  nand n12620(x12620, x12619, x12618);
  nand n12621(x12621, x2258, x6111);
  nand n12622(x12622, x6481, x5981);
  nand n12623(x12623, x12622, x12621);
  nand n12624(x12624, x2258, x5851);
  nand n12625(x12625, x6481, x5721);
  nand n12626(x12626, x12625, x12624);
  nand n12627(x12627, x2258, x5591);
  nand n12628(x12628, x6481, x5461);
  nand n12629(x12629, x12628, x12627);
  nand n12630(x12630, x2261, x12620);
  nand n12631(x12631, x6494, x12623);
  nand n12632(x12632, x12631, x12630);
  nand n12633(x12633, x2261, x12626);
  nand n12634(x12634, x6494, x12629);
  nand n12635(x12635, x12634, x12633);
  nand n12636(x12636, x2264, x12632);
  nand n12637(x12637, x6501, x12635);
  nand n12638(x12638, x12637, x12636);
  nand n12639(x12639, x2258, x6375);
  nand n12640(x12640, x6481, x6245);
  nand n12641(x12641, x12640, x12639);
  nand n12642(x12642, x2258, x6115);
  nand n12643(x12643, x6481, x5985);
  nand n12644(x12644, x12643, x12642);
  nand n12645(x12645, x2258, x5855);
  nand n12646(x12646, x6481, x5725);
  nand n12647(x12647, x12646, x12645);
  nand n12648(x12648, x2258, x5595);
  nand n12649(x12649, x6481, x5465);
  nand n12650(x12650, x12649, x12648);
  nand n12651(x12651, x2261, x12641);
  nand n12652(x12652, x6494, x12644);
  nand n12653(x12653, x12652, x12651);
  nand n12654(x12654, x2261, x12647);
  nand n12655(x12655, x6494, x12650);
  nand n12656(x12656, x12655, x12654);
  nand n12657(x12657, x2264, x12653);
  nand n12658(x12658, x6501, x12656);
  nand n12659(x12659, x12658, x12657);
  nand n12660(x12660, x2258, x6379);
  nand n12661(x12661, x6481, x6249);
  nand n12662(x12662, x12661, x12660);
  nand n12663(x12663, x2258, x6119);
  nand n12664(x12664, x6481, x5989);
  nand n12665(x12665, x12664, x12663);
  nand n12666(x12666, x2258, x5859);
  nand n12667(x12667, x6481, x5729);
  nand n12668(x12668, x12667, x12666);
  nand n12669(x12669, x2258, x5599);
  nand n12670(x12670, x6481, x5469);
  nand n12671(x12671, x12670, x12669);
  nand n12672(x12672, x2261, x12662);
  nand n12673(x12673, x6494, x12665);
  nand n12674(x12674, x12673, x12672);
  nand n12675(x12675, x2261, x12668);
  nand n12676(x12676, x6494, x12671);
  nand n12677(x12677, x12676, x12675);
  nand n12678(x12678, x2264, x12674);
  nand n12679(x12679, x6501, x12677);
  nand n12680(x12680, x12679, x12678);
  nand n12681(x12681, x2258, x6383);
  nand n12682(x12682, x6481, x6253);
  nand n12683(x12683, x12682, x12681);
  nand n12684(x12684, x2258, x6123);
  nand n12685(x12685, x6481, x5993);
  nand n12686(x12686, x12685, x12684);
  nand n12687(x12687, x2258, x5863);
  nand n12688(x12688, x6481, x5733);
  nand n12689(x12689, x12688, x12687);
  nand n12690(x12690, x2258, x5603);
  nand n12691(x12691, x6481, x5473);
  nand n12692(x12692, x12691, x12690);
  nand n12693(x12693, x2261, x12683);
  nand n12694(x12694, x6494, x12686);
  nand n12695(x12695, x12694, x12693);
  nand n12696(x12696, x2261, x12689);
  nand n12697(x12697, x6494, x12692);
  nand n12698(x12698, x12697, x12696);
  nand n12699(x12699, x2264, x12695);
  nand n12700(x12700, x6501, x12698);
  nand n12701(x12701, x12700, x12699);
  nand n12702(x12702, x2258, x6387);
  nand n12703(x12703, x6481, x6257);
  nand n12704(x12704, x12703, x12702);
  nand n12705(x12705, x2258, x6127);
  nand n12706(x12706, x6481, x5997);
  nand n12707(x12707, x12706, x12705);
  nand n12708(x12708, x2258, x5867);
  nand n12709(x12709, x6481, x5737);
  nand n12710(x12710, x12709, x12708);
  nand n12711(x12711, x2258, x5607);
  nand n12712(x12712, x6481, x5477);
  nand n12713(x12713, x12712, x12711);
  nand n12714(x12714, x2261, x12704);
  nand n12715(x12715, x6494, x12707);
  nand n12716(x12716, x12715, x12714);
  nand n12717(x12717, x2261, x12710);
  nand n12718(x12718, x6494, x12713);
  nand n12719(x12719, x12718, x12717);
  nand n12720(x12720, x2264, x12716);
  nand n12721(x12721, x6501, x12719);
  nand n12722(x12722, x12721, x12720);
  nand n12723(x12723, x2258, x6391);
  nand n12724(x12724, x6481, x6261);
  nand n12725(x12725, x12724, x12723);
  nand n12726(x12726, x2258, x6131);
  nand n12727(x12727, x6481, x6001);
  nand n12728(x12728, x12727, x12726);
  nand n12729(x12729, x2258, x5871);
  nand n12730(x12730, x6481, x5741);
  nand n12731(x12731, x12730, x12729);
  nand n12732(x12732, x2258, x5611);
  nand n12733(x12733, x6481, x5481);
  nand n12734(x12734, x12733, x12732);
  nand n12735(x12735, x2261, x12725);
  nand n12736(x12736, x6494, x12728);
  nand n12737(x12737, x12736, x12735);
  nand n12738(x12738, x2261, x12731);
  nand n12739(x12739, x6494, x12734);
  nand n12740(x12740, x12739, x12738);
  nand n12741(x12741, x2264, x12737);
  nand n12742(x12742, x6501, x12740);
  nand n12743(x12743, x12742, x12741);
  nand n12744(x12744, x2258, x6395);
  nand n12745(x12745, x6481, x6265);
  nand n12746(x12746, x12745, x12744);
  nand n12747(x12747, x2258, x6135);
  nand n12748(x12748, x6481, x6005);
  nand n12749(x12749, x12748, x12747);
  nand n12750(x12750, x2258, x5875);
  nand n12751(x12751, x6481, x5745);
  nand n12752(x12752, x12751, x12750);
  nand n12753(x12753, x2258, x5615);
  nand n12754(x12754, x6481, x5485);
  nand n12755(x12755, x12754, x12753);
  nand n12756(x12756, x2261, x12746);
  nand n12757(x12757, x6494, x12749);
  nand n12758(x12758, x12757, x12756);
  nand n12759(x12759, x2261, x12752);
  nand n12760(x12760, x6494, x12755);
  nand n12761(x12761, x12760, x12759);
  nand n12762(x12762, x2264, x12758);
  nand n12763(x12763, x6501, x12761);
  nand n12764(x12764, x12763, x12762);
  nand n12765(x12765, x2258, x6399);
  nand n12766(x12766, x6481, x6269);
  nand n12767(x12767, x12766, x12765);
  nand n12768(x12768, x2258, x6139);
  nand n12769(x12769, x6481, x6009);
  nand n12770(x12770, x12769, x12768);
  nand n12771(x12771, x2258, x5879);
  nand n12772(x12772, x6481, x5749);
  nand n12773(x12773, x12772, x12771);
  nand n12774(x12774, x2258, x5619);
  nand n12775(x12775, x6481, x5489);
  nand n12776(x12776, x12775, x12774);
  nand n12777(x12777, x2261, x12767);
  nand n12778(x12778, x6494, x12770);
  nand n12779(x12779, x12778, x12777);
  nand n12780(x12780, x2261, x12773);
  nand n12781(x12781, x6494, x12776);
  nand n12782(x12782, x12781, x12780);
  nand n12783(x12783, x2264, x12779);
  nand n12784(x12784, x6501, x12782);
  nand n12785(x12785, x12784, x12783);
  nand n12786(x12786, x2258, x6403);
  nand n12787(x12787, x6481, x6273);
  nand n12788(x12788, x12787, x12786);
  nand n12789(x12789, x2258, x6143);
  nand n12790(x12790, x6481, x6013);
  nand n12791(x12791, x12790, x12789);
  nand n12792(x12792, x2258, x5883);
  nand n12793(x12793, x6481, x5753);
  nand n12794(x12794, x12793, x12792);
  nand n12795(x12795, x2258, x5623);
  nand n12796(x12796, x6481, x5493);
  nand n12797(x12797, x12796, x12795);
  nand n12798(x12798, x2261, x12788);
  nand n12799(x12799, x6494, x12791);
  nand n12800(x12800, x12799, x12798);
  nand n12801(x12801, x2261, x12794);
  nand n12802(x12802, x6494, x12797);
  nand n12803(x12803, x12802, x12801);
  nand n12804(x12804, x2264, x12800);
  nand n12805(x12805, x6501, x12803);
  nand n12806(x12806, x12805, x12804);
  nand n12807(x12807, x2258, x6407);
  nand n12808(x12808, x6481, x6277);
  nand n12809(x12809, x12808, x12807);
  nand n12810(x12810, x2258, x6147);
  nand n12811(x12811, x6481, x6017);
  nand n12812(x12812, x12811, x12810);
  nand n12813(x12813, x2258, x5887);
  nand n12814(x12814, x6481, x5757);
  nand n12815(x12815, x12814, x12813);
  nand n12816(x12816, x2258, x5627);
  nand n12817(x12817, x6481, x5497);
  nand n12818(x12818, x12817, x12816);
  nand n12819(x12819, x2261, x12809);
  nand n12820(x12820, x6494, x12812);
  nand n12821(x12821, x12820, x12819);
  nand n12822(x12822, x2261, x12815);
  nand n12823(x12823, x6494, x12818);
  nand n12824(x12824, x12823, x12822);
  nand n12825(x12825, x2264, x12821);
  nand n12826(x12826, x6501, x12824);
  nand n12827(x12827, x12826, x12825);
  nand n12828(x12828, x2258, x6411);
  nand n12829(x12829, x6481, x6281);
  nand n12830(x12830, x12829, x12828);
  nand n12831(x12831, x2258, x6151);
  nand n12832(x12832, x6481, x6021);
  nand n12833(x12833, x12832, x12831);
  nand n12834(x12834, x2258, x5891);
  nand n12835(x12835, x6481, x5761);
  nand n12836(x12836, x12835, x12834);
  nand n12837(x12837, x2258, x5631);
  nand n12838(x12838, x6481, x5501);
  nand n12839(x12839, x12838, x12837);
  nand n12840(x12840, x2261, x12830);
  nand n12841(x12841, x6494, x12833);
  nand n12842(x12842, x12841, x12840);
  nand n12843(x12843, x2261, x12836);
  nand n12844(x12844, x6494, x12839);
  nand n12845(x12845, x12844, x12843);
  nand n12846(x12846, x2264, x12842);
  nand n12847(x12847, x6501, x12845);
  nand n12848(x12848, x12847, x12846);
  nand n12849(x12849, x2258, x6415);
  nand n12850(x12850, x6481, x6285);
  nand n12851(x12851, x12850, x12849);
  nand n12852(x12852, x2258, x6155);
  nand n12853(x12853, x6481, x6025);
  nand n12854(x12854, x12853, x12852);
  nand n12855(x12855, x2258, x5895);
  nand n12856(x12856, x6481, x5765);
  nand n12857(x12857, x12856, x12855);
  nand n12858(x12858, x2258, x5635);
  nand n12859(x12859, x6481, x5505);
  nand n12860(x12860, x12859, x12858);
  nand n12861(x12861, x2261, x12851);
  nand n12862(x12862, x6494, x12854);
  nand n12863(x12863, x12862, x12861);
  nand n12864(x12864, x2261, x12857);
  nand n12865(x12865, x6494, x12860);
  nand n12866(x12866, x12865, x12864);
  nand n12867(x12867, x2264, x12863);
  nand n12868(x12868, x6501, x12866);
  nand n12869(x12869, x12868, x12867);
  nand n12870(x12870, x2258, x6419);
  nand n12871(x12871, x6481, x6289);
  nand n12872(x12872, x12871, x12870);
  nand n12873(x12873, x2258, x6159);
  nand n12874(x12874, x6481, x6029);
  nand n12875(x12875, x12874, x12873);
  nand n12876(x12876, x2258, x5899);
  nand n12877(x12877, x6481, x5769);
  nand n12878(x12878, x12877, x12876);
  nand n12879(x12879, x2258, x5639);
  nand n12880(x12880, x6481, x5509);
  nand n12881(x12881, x12880, x12879);
  nand n12882(x12882, x2261, x12872);
  nand n12883(x12883, x6494, x12875);
  nand n12884(x12884, x12883, x12882);
  nand n12885(x12885, x2261, x12878);
  nand n12886(x12886, x6494, x12881);
  nand n12887(x12887, x12886, x12885);
  nand n12888(x12888, x2264, x12884);
  nand n12889(x12889, x6501, x12887);
  nand n12890(x12890, x12889, x12888);
  nand n12891(x12891, x2258, x6423);
  nand n12892(x12892, x6481, x6293);
  nand n12893(x12893, x12892, x12891);
  nand n12894(x12894, x2258, x6163);
  nand n12895(x12895, x6481, x6033);
  nand n12896(x12896, x12895, x12894);
  nand n12897(x12897, x2258, x5903);
  nand n12898(x12898, x6481, x5773);
  nand n12899(x12899, x12898, x12897);
  nand n12900(x12900, x2258, x5643);
  nand n12901(x12901, x6481, x5513);
  nand n12902(x12902, x12901, x12900);
  nand n12903(x12903, x2261, x12893);
  nand n12904(x12904, x6494, x12896);
  nand n12905(x12905, x12904, x12903);
  nand n12906(x12906, x2261, x12899);
  nand n12907(x12907, x6494, x12902);
  nand n12908(x12908, x12907, x12906);
  nand n12909(x12909, x2264, x12905);
  nand n12910(x12910, x6501, x12908);
  nand n12911(x12911, x12910, x12909);
  nand n12912(x12912, x2258, x6427);
  nand n12913(x12913, x6481, x6297);
  nand n12914(x12914, x12913, x12912);
  nand n12915(x12915, x2258, x6167);
  nand n12916(x12916, x6481, x6037);
  nand n12917(x12917, x12916, x12915);
  nand n12918(x12918, x2258, x5907);
  nand n12919(x12919, x6481, x5777);
  nand n12920(x12920, x12919, x12918);
  nand n12921(x12921, x2258, x5647);
  nand n12922(x12922, x6481, x5517);
  nand n12923(x12923, x12922, x12921);
  nand n12924(x12924, x2261, x12914);
  nand n12925(x12925, x6494, x12917);
  nand n12926(x12926, x12925, x12924);
  nand n12927(x12927, x2261, x12920);
  nand n12928(x12928, x6494, x12923);
  nand n12929(x12929, x12928, x12927);
  nand n12930(x12930, x2264, x12926);
  nand n12931(x12931, x6501, x12929);
  nand n12932(x12932, x12931, x12930);
  nand n12933(x12933, x2258, x6431);
  nand n12934(x12934, x6481, x6301);
  nand n12935(x12935, x12934, x12933);
  nand n12936(x12936, x2258, x6171);
  nand n12937(x12937, x6481, x6041);
  nand n12938(x12938, x12937, x12936);
  nand n12939(x12939, x2258, x5911);
  nand n12940(x12940, x6481, x5781);
  nand n12941(x12941, x12940, x12939);
  nand n12942(x12942, x2258, x5651);
  nand n12943(x12943, x6481, x5521);
  nand n12944(x12944, x12943, x12942);
  nand n12945(x12945, x2261, x12935);
  nand n12946(x12946, x6494, x12938);
  nand n12947(x12947, x12946, x12945);
  nand n12948(x12948, x2261, x12941);
  nand n12949(x12949, x6494, x12944);
  nand n12950(x12950, x12949, x12948);
  nand n12951(x12951, x2264, x12947);
  nand n12952(x12952, x6501, x12950);
  nand n12953(x12953, x12952, x12951);
  nand n12954(x12954, x2258, x6435);
  nand n12955(x12955, x6481, x6305);
  nand n12956(x12956, x12955, x12954);
  nand n12957(x12957, x2258, x6175);
  nand n12958(x12958, x6481, x6045);
  nand n12959(x12959, x12958, x12957);
  nand n12960(x12960, x2258, x5915);
  nand n12961(x12961, x6481, x5785);
  nand n12962(x12962, x12961, x12960);
  nand n12963(x12963, x2258, x5655);
  nand n12964(x12964, x6481, x5525);
  nand n12965(x12965, x12964, x12963);
  nand n12966(x12966, x2261, x12956);
  nand n12967(x12967, x6494, x12959);
  nand n12968(x12968, x12967, x12966);
  nand n12969(x12969, x2261, x12962);
  nand n12970(x12970, x6494, x12965);
  nand n12971(x12971, x12970, x12969);
  nand n12972(x12972, x2264, x12968);
  nand n12973(x12973, x6501, x12971);
  nand n12974(x12974, x12973, x12972);
  nand n12975(x12975, x2258, x6439);
  nand n12976(x12976, x6481, x6309);
  nand n12977(x12977, x12976, x12975);
  nand n12978(x12978, x2258, x6179);
  nand n12979(x12979, x6481, x6049);
  nand n12980(x12980, x12979, x12978);
  nand n12981(x12981, x2258, x5919);
  nand n12982(x12982, x6481, x5789);
  nand n12983(x12983, x12982, x12981);
  nand n12984(x12984, x2258, x5659);
  nand n12985(x12985, x6481, x5529);
  nand n12986(x12986, x12985, x12984);
  nand n12987(x12987, x2261, x12977);
  nand n12988(x12988, x6494, x12980);
  nand n12989(x12989, x12988, x12987);
  nand n12990(x12990, x2261, x12983);
  nand n12991(x12991, x6494, x12986);
  nand n12992(x12992, x12991, x12990);
  nand n12993(x12993, x2264, x12989);
  nand n12994(x12994, x6501, x12992);
  nand n12995(x12995, x12994, x12993);
  nand n12996(x12996, x2258, x6443);
  nand n12997(x12997, x6481, x6313);
  nand n12998(x12998, x12997, x12996);
  nand n12999(x12999, x2258, x6183);
  nand n13000(x13000, x6481, x6053);
  nand n13001(x13001, x13000, x12999);
  nand n13002(x13002, x2258, x5923);
  nand n13003(x13003, x6481, x5793);
  nand n13004(x13004, x13003, x13002);
  nand n13005(x13005, x2258, x5663);
  nand n13006(x13006, x6481, x5533);
  nand n13007(x13007, x13006, x13005);
  nand n13008(x13008, x2261, x12998);
  nand n13009(x13009, x6494, x13001);
  nand n13010(x13010, x13009, x13008);
  nand n13011(x13011, x2261, x13004);
  nand n13012(x13012, x6494, x13007);
  nand n13013(x13013, x13012, x13011);
  nand n13014(x13014, x2264, x13010);
  nand n13015(x13015, x6501, x13013);
  nand n13016(x13016, x13015, x13014);
  nand n13017(x13017, x2258, x6447);
  nand n13018(x13018, x6481, x6317);
  nand n13019(x13019, x13018, x13017);
  nand n13020(x13020, x2258, x6187);
  nand n13021(x13021, x6481, x6057);
  nand n13022(x13022, x13021, x13020);
  nand n13023(x13023, x2258, x5927);
  nand n13024(x13024, x6481, x5797);
  nand n13025(x13025, x13024, x13023);
  nand n13026(x13026, x2258, x5667);
  nand n13027(x13027, x6481, x5537);
  nand n13028(x13028, x13027, x13026);
  nand n13029(x13029, x2261, x13019);
  nand n13030(x13030, x6494, x13022);
  nand n13031(x13031, x13030, x13029);
  nand n13032(x13032, x2261, x13025);
  nand n13033(x13033, x6494, x13028);
  nand n13034(x13034, x13033, x13032);
  nand n13035(x13035, x2264, x13031);
  nand n13036(x13036, x6501, x13034);
  nand n13037(x13037, x13036, x13035);
  nand n13038(x13038, x2258, x6451);
  nand n13039(x13039, x6481, x6321);
  nand n13040(x13040, x13039, x13038);
  nand n13041(x13041, x2258, x6191);
  nand n13042(x13042, x6481, x6061);
  nand n13043(x13043, x13042, x13041);
  nand n13044(x13044, x2258, x5931);
  nand n13045(x13045, x6481, x5801);
  nand n13046(x13046, x13045, x13044);
  nand n13047(x13047, x2258, x5671);
  nand n13048(x13048, x6481, x5541);
  nand n13049(x13049, x13048, x13047);
  nand n13050(x13050, x2261, x13040);
  nand n13051(x13051, x6494, x13043);
  nand n13052(x13052, x13051, x13050);
  nand n13053(x13053, x2261, x13046);
  nand n13054(x13054, x6494, x13049);
  nand n13055(x13055, x13054, x13053);
  nand n13056(x13056, x2264, x13052);
  nand n13057(x13057, x6501, x13055);
  nand n13058(x13058, x13057, x13056);
  nand n13059(x13059, x2258, x6455);
  nand n13060(x13060, x6481, x6325);
  nand n13061(x13061, x13060, x13059);
  nand n13062(x13062, x2258, x6195);
  nand n13063(x13063, x6481, x6065);
  nand n13064(x13064, x13063, x13062);
  nand n13065(x13065, x2258, x5935);
  nand n13066(x13066, x6481, x5805);
  nand n13067(x13067, x13066, x13065);
  nand n13068(x13068, x2258, x5675);
  nand n13069(x13069, x6481, x5545);
  nand n13070(x13070, x13069, x13068);
  nand n13071(x13071, x2261, x13061);
  nand n13072(x13072, x6494, x13064);
  nand n13073(x13073, x13072, x13071);
  nand n13074(x13074, x2261, x13067);
  nand n13075(x13075, x6494, x13070);
  nand n13076(x13076, x13075, x13074);
  nand n13077(x13077, x2264, x13073);
  nand n13078(x13078, x6501, x13076);
  nand n13079(x13079, x13078, x13077);
  nand n13080(x13080, x2258, x6459);
  nand n13081(x13081, x6481, x6329);
  nand n13082(x13082, x13081, x13080);
  nand n13083(x13083, x2258, x6199);
  nand n13084(x13084, x6481, x6069);
  nand n13085(x13085, x13084, x13083);
  nand n13086(x13086, x2258, x5939);
  nand n13087(x13087, x6481, x5809);
  nand n13088(x13088, x13087, x13086);
  nand n13089(x13089, x2258, x5679);
  nand n13090(x13090, x6481, x5549);
  nand n13091(x13091, x13090, x13089);
  nand n13092(x13092, x2261, x13082);
  nand n13093(x13093, x6494, x13085);
  nand n13094(x13094, x13093, x13092);
  nand n13095(x13095, x2261, x13088);
  nand n13096(x13096, x6494, x13091);
  nand n13097(x13097, x13096, x13095);
  nand n13098(x13098, x2264, x13094);
  nand n13099(x13099, x6501, x13097);
  nand n13100(x13100, x13099, x13098);
  nand n13101(x13101, x2258, x6463);
  nand n13102(x13102, x6481, x6333);
  nand n13103(x13103, x13102, x13101);
  nand n13104(x13104, x2258, x6203);
  nand n13105(x13105, x6481, x6073);
  nand n13106(x13106, x13105, x13104);
  nand n13107(x13107, x2258, x5943);
  nand n13108(x13108, x6481, x5813);
  nand n13109(x13109, x13108, x13107);
  nand n13110(x13110, x2258, x5683);
  nand n13111(x13111, x6481, x5553);
  nand n13112(x13112, x13111, x13110);
  nand n13113(x13113, x2261, x13103);
  nand n13114(x13114, x6494, x13106);
  nand n13115(x13115, x13114, x13113);
  nand n13116(x13116, x2261, x13109);
  nand n13117(x13117, x6494, x13112);
  nand n13118(x13118, x13117, x13116);
  nand n13119(x13119, x2264, x13115);
  nand n13120(x13120, x6501, x13118);
  nand n13121(x13121, x13120, x13119);
  nand n13122(x13122, x2258, x6467);
  nand n13123(x13123, x6481, x6337);
  nand n13124(x13124, x13123, x13122);
  nand n13125(x13125, x2258, x6207);
  nand n13126(x13126, x6481, x6077);
  nand n13127(x13127, x13126, x13125);
  nand n13128(x13128, x2258, x5947);
  nand n13129(x13129, x6481, x5817);
  nand n13130(x13130, x13129, x13128);
  nand n13131(x13131, x2258, x5687);
  nand n13132(x13132, x6481, x5557);
  nand n13133(x13133, x13132, x13131);
  nand n13134(x13134, x2261, x13124);
  nand n13135(x13135, x6494, x13127);
  nand n13136(x13136, x13135, x13134);
  nand n13137(x13137, x2261, x13130);
  nand n13138(x13138, x6494, x13133);
  nand n13139(x13139, x13138, x13137);
  nand n13140(x13140, x2264, x13136);
  nand n13141(x13141, x6501, x13139);
  nand n13142(x13142, x13141, x13140);
  nand n13143(x13143, x2258, x6471);
  nand n13144(x13144, x6481, x6341);
  nand n13145(x13145, x13144, x13143);
  nand n13146(x13146, x2258, x6211);
  nand n13147(x13147, x6481, x6081);
  nand n13148(x13148, x13147, x13146);
  nand n13149(x13149, x2258, x5951);
  nand n13150(x13150, x6481, x5821);
  nand n13151(x13151, x13150, x13149);
  nand n13152(x13152, x2258, x5691);
  nand n13153(x13153, x6481, x5561);
  nand n13154(x13154, x13153, x13152);
  nand n13155(x13155, x2261, x13145);
  nand n13156(x13156, x6494, x13148);
  nand n13157(x13157, x13156, x13155);
  nand n13158(x13158, x2261, x13151);
  nand n13159(x13159, x6494, x13154);
  nand n13160(x13160, x13159, x13158);
  nand n13161(x13161, x2264, x13157);
  nand n13162(x13162, x6501, x13160);
  nand n13163(x13163, x13162, x13161);
  nand n13164(x13164, x2258, x6475);
  nand n13165(x13165, x6481, x6345);
  nand n13166(x13166, x13165, x13164);
  nand n13167(x13167, x2258, x6215);
  nand n13168(x13168, x6481, x6085);
  nand n13169(x13169, x13168, x13167);
  nand n13170(x13170, x2258, x5955);
  nand n13171(x13171, x6481, x5825);
  nand n13172(x13172, x13171, x13170);
  nand n13173(x13173, x2258, x5695);
  nand n13174(x13174, x6481, x5565);
  nand n13175(x13175, x13174, x13173);
  nand n13176(x13176, x2261, x13166);
  nand n13177(x13177, x6494, x13169);
  nand n13178(x13178, x13177, x13176);
  nand n13179(x13179, x2261, x13172);
  nand n13180(x13180, x6494, x13175);
  nand n13181(x13181, x13180, x13179);
  nand n13182(x13182, x2264, x13178);
  nand n13183(x13183, x6501, x13181);
  nand n13184(x13184, x13183, x13182);
  nand n13185(x13185, x2258, x6479);
  nand n13186(x13186, x6481, x6349);
  nand n13187(x13187, x13186, x13185);
  nand n13188(x13188, x2258, x6219);
  nand n13189(x13189, x6481, x6089);
  nand n13190(x13190, x13189, x13188);
  nand n13191(x13191, x2258, x5959);
  nand n13192(x13192, x6481, x5829);
  nand n13193(x13193, x13192, x13191);
  nand n13194(x13194, x2258, x5699);
  nand n13195(x13195, x6481, x5569);
  nand n13196(x13196, x13195, x13194);
  nand n13197(x13197, x2261, x13187);
  nand n13198(x13198, x6494, x13190);
  nand n13199(x13199, x13198, x13197);
  nand n13200(x13200, x2261, x13193);
  nand n13201(x13201, x6494, x13196);
  nand n13202(x13202, x13201, x13200);
  nand n13203(x13203, x2264, x13199);
  nand n13204(x13204, x6501, x13202);
  nand n13205(x13205, x13204, x13203);
  nand n13206(x13206, x2269, x6355);
  nand n13207(x13207, x7156, x6225);
  nand n13208(x13208, x13207, x13206);
  nand n13209(x13209, x2269, x6095);
  nand n13210(x13210, x7156, x5965);
  nand n13211(x13211, x13210, x13209);
  nand n13212(x13212, x2269, x5835);
  nand n13213(x13213, x7156, x5705);
  nand n13214(x13214, x13213, x13212);
  nand n13215(x13215, x2269, x5575);
  nand n13216(x13216, x7156, x5443);
  nand n13217(x13217, x13216, x13215);
  nand n13218(x13218, x2272, x13208);
  nand n13219(x13219, x7169, x13211);
  nand n13220(x13220, x13219, x13218);
  nand n13221(x13221, x2272, x13214);
  nand n13222(x13222, x7169, x13217);
  nand n13223(x13223, x13222, x13221);
  nand n13224(x13224, x2275, x13220);
  nand n13225(x13225, x7176, x13223);
  nand n13226(x13226, x13225, x13224);
  nand n13227(x13227, x2269, x6359);
  nand n13228(x13228, x7156, x6229);
  nand n13229(x13229, x13228, x13227);
  nand n13230(x13230, x2269, x6099);
  nand n13231(x13231, x7156, x5969);
  nand n13232(x13232, x13231, x13230);
  nand n13233(x13233, x2269, x5839);
  nand n13234(x13234, x7156, x5709);
  nand n13235(x13235, x13234, x13233);
  nand n13236(x13236, x2269, x5579);
  nand n13237(x13237, x7156, x5449);
  nand n13238(x13238, x13237, x13236);
  nand n13239(x13239, x2272, x13229);
  nand n13240(x13240, x7169, x13232);
  nand n13241(x13241, x13240, x13239);
  nand n13242(x13242, x2272, x13235);
  nand n13243(x13243, x7169, x13238);
  nand n13244(x13244, x13243, x13242);
  nand n13245(x13245, x2275, x13241);
  nand n13246(x13246, x7176, x13244);
  nand n13247(x13247, x13246, x13245);
  nand n13248(x13248, x2269, x6363);
  nand n13249(x13249, x7156, x6233);
  nand n13250(x13250, x13249, x13248);
  nand n13251(x13251, x2269, x6103);
  nand n13252(x13252, x7156, x5973);
  nand n13253(x13253, x13252, x13251);
  nand n13254(x13254, x2269, x5843);
  nand n13255(x13255, x7156, x5713);
  nand n13256(x13256, x13255, x13254);
  nand n13257(x13257, x2269, x5583);
  nand n13258(x13258, x7156, x5453);
  nand n13259(x13259, x13258, x13257);
  nand n13260(x13260, x2272, x13250);
  nand n13261(x13261, x7169, x13253);
  nand n13262(x13262, x13261, x13260);
  nand n13263(x13263, x2272, x13256);
  nand n13264(x13264, x7169, x13259);
  nand n13265(x13265, x13264, x13263);
  nand n13266(x13266, x2275, x13262);
  nand n13267(x13267, x7176, x13265);
  nand n13268(x13268, x13267, x13266);
  nand n13269(x13269, x2269, x6367);
  nand n13270(x13270, x7156, x6237);
  nand n13271(x13271, x13270, x13269);
  nand n13272(x13272, x2269, x6107);
  nand n13273(x13273, x7156, x5977);
  nand n13274(x13274, x13273, x13272);
  nand n13275(x13275, x2269, x5847);
  nand n13276(x13276, x7156, x5717);
  nand n13277(x13277, x13276, x13275);
  nand n13278(x13278, x2269, x5587);
  nand n13279(x13279, x7156, x5457);
  nand n13280(x13280, x13279, x13278);
  nand n13281(x13281, x2272, x13271);
  nand n13282(x13282, x7169, x13274);
  nand n13283(x13283, x13282, x13281);
  nand n13284(x13284, x2272, x13277);
  nand n13285(x13285, x7169, x13280);
  nand n13286(x13286, x13285, x13284);
  nand n13287(x13287, x2275, x13283);
  nand n13288(x13288, x7176, x13286);
  nand n13289(x13289, x13288, x13287);
  nand n13290(x13290, x2269, x6371);
  nand n13291(x13291, x7156, x6241);
  nand n13292(x13292, x13291, x13290);
  nand n13293(x13293, x2269, x6111);
  nand n13294(x13294, x7156, x5981);
  nand n13295(x13295, x13294, x13293);
  nand n13296(x13296, x2269, x5851);
  nand n13297(x13297, x7156, x5721);
  nand n13298(x13298, x13297, x13296);
  nand n13299(x13299, x2269, x5591);
  nand n13300(x13300, x7156, x5461);
  nand n13301(x13301, x13300, x13299);
  nand n13302(x13302, x2272, x13292);
  nand n13303(x13303, x7169, x13295);
  nand n13304(x13304, x13303, x13302);
  nand n13305(x13305, x2272, x13298);
  nand n13306(x13306, x7169, x13301);
  nand n13307(x13307, x13306, x13305);
  nand n13308(x13308, x2275, x13304);
  nand n13309(x13309, x7176, x13307);
  nand n13310(x13310, x13309, x13308);
  nand n13311(x13311, x2269, x6375);
  nand n13312(x13312, x7156, x6245);
  nand n13313(x13313, x13312, x13311);
  nand n13314(x13314, x2269, x6115);
  nand n13315(x13315, x7156, x5985);
  nand n13316(x13316, x13315, x13314);
  nand n13317(x13317, x2269, x5855);
  nand n13318(x13318, x7156, x5725);
  nand n13319(x13319, x13318, x13317);
  nand n13320(x13320, x2269, x5595);
  nand n13321(x13321, x7156, x5465);
  nand n13322(x13322, x13321, x13320);
  nand n13323(x13323, x2272, x13313);
  nand n13324(x13324, x7169, x13316);
  nand n13325(x13325, x13324, x13323);
  nand n13326(x13326, x2272, x13319);
  nand n13327(x13327, x7169, x13322);
  nand n13328(x13328, x13327, x13326);
  nand n13329(x13329, x2275, x13325);
  nand n13330(x13330, x7176, x13328);
  nand n13331(x13331, x13330, x13329);
  nand n13332(x13332, x2269, x6379);
  nand n13333(x13333, x7156, x6249);
  nand n13334(x13334, x13333, x13332);
  nand n13335(x13335, x2269, x6119);
  nand n13336(x13336, x7156, x5989);
  nand n13337(x13337, x13336, x13335);
  nand n13338(x13338, x2269, x5859);
  nand n13339(x13339, x7156, x5729);
  nand n13340(x13340, x13339, x13338);
  nand n13341(x13341, x2269, x5599);
  nand n13342(x13342, x7156, x5469);
  nand n13343(x13343, x13342, x13341);
  nand n13344(x13344, x2272, x13334);
  nand n13345(x13345, x7169, x13337);
  nand n13346(x13346, x13345, x13344);
  nand n13347(x13347, x2272, x13340);
  nand n13348(x13348, x7169, x13343);
  nand n13349(x13349, x13348, x13347);
  nand n13350(x13350, x2275, x13346);
  nand n13351(x13351, x7176, x13349);
  nand n13352(x13352, x13351, x13350);
  nand n13353(x13353, x2269, x6383);
  nand n13354(x13354, x7156, x6253);
  nand n13355(x13355, x13354, x13353);
  nand n13356(x13356, x2269, x6123);
  nand n13357(x13357, x7156, x5993);
  nand n13358(x13358, x13357, x13356);
  nand n13359(x13359, x2269, x5863);
  nand n13360(x13360, x7156, x5733);
  nand n13361(x13361, x13360, x13359);
  nand n13362(x13362, x2269, x5603);
  nand n13363(x13363, x7156, x5473);
  nand n13364(x13364, x13363, x13362);
  nand n13365(x13365, x2272, x13355);
  nand n13366(x13366, x7169, x13358);
  nand n13367(x13367, x13366, x13365);
  nand n13368(x13368, x2272, x13361);
  nand n13369(x13369, x7169, x13364);
  nand n13370(x13370, x13369, x13368);
  nand n13371(x13371, x2275, x13367);
  nand n13372(x13372, x7176, x13370);
  nand n13373(x13373, x13372, x13371);
  nand n13374(x13374, x2269, x6387);
  nand n13375(x13375, x7156, x6257);
  nand n13376(x13376, x13375, x13374);
  nand n13377(x13377, x2269, x6127);
  nand n13378(x13378, x7156, x5997);
  nand n13379(x13379, x13378, x13377);
  nand n13380(x13380, x2269, x5867);
  nand n13381(x13381, x7156, x5737);
  nand n13382(x13382, x13381, x13380);
  nand n13383(x13383, x2269, x5607);
  nand n13384(x13384, x7156, x5477);
  nand n13385(x13385, x13384, x13383);
  nand n13386(x13386, x2272, x13376);
  nand n13387(x13387, x7169, x13379);
  nand n13388(x13388, x13387, x13386);
  nand n13389(x13389, x2272, x13382);
  nand n13390(x13390, x7169, x13385);
  nand n13391(x13391, x13390, x13389);
  nand n13392(x13392, x2275, x13388);
  nand n13393(x13393, x7176, x13391);
  nand n13394(x13394, x13393, x13392);
  nand n13395(x13395, x2269, x6391);
  nand n13396(x13396, x7156, x6261);
  nand n13397(x13397, x13396, x13395);
  nand n13398(x13398, x2269, x6131);
  nand n13399(x13399, x7156, x6001);
  nand n13400(x13400, x13399, x13398);
  nand n13401(x13401, x2269, x5871);
  nand n13402(x13402, x7156, x5741);
  nand n13403(x13403, x13402, x13401);
  nand n13404(x13404, x2269, x5611);
  nand n13405(x13405, x7156, x5481);
  nand n13406(x13406, x13405, x13404);
  nand n13407(x13407, x2272, x13397);
  nand n13408(x13408, x7169, x13400);
  nand n13409(x13409, x13408, x13407);
  nand n13410(x13410, x2272, x13403);
  nand n13411(x13411, x7169, x13406);
  nand n13412(x13412, x13411, x13410);
  nand n13413(x13413, x2275, x13409);
  nand n13414(x13414, x7176, x13412);
  nand n13415(x13415, x13414, x13413);
  nand n13416(x13416, x2269, x6395);
  nand n13417(x13417, x7156, x6265);
  nand n13418(x13418, x13417, x13416);
  nand n13419(x13419, x2269, x6135);
  nand n13420(x13420, x7156, x6005);
  nand n13421(x13421, x13420, x13419);
  nand n13422(x13422, x2269, x5875);
  nand n13423(x13423, x7156, x5745);
  nand n13424(x13424, x13423, x13422);
  nand n13425(x13425, x2269, x5615);
  nand n13426(x13426, x7156, x5485);
  nand n13427(x13427, x13426, x13425);
  nand n13428(x13428, x2272, x13418);
  nand n13429(x13429, x7169, x13421);
  nand n13430(x13430, x13429, x13428);
  nand n13431(x13431, x2272, x13424);
  nand n13432(x13432, x7169, x13427);
  nand n13433(x13433, x13432, x13431);
  nand n13434(x13434, x2275, x13430);
  nand n13435(x13435, x7176, x13433);
  nand n13436(x13436, x13435, x13434);
  nand n13437(x13437, x2269, x6399);
  nand n13438(x13438, x7156, x6269);
  nand n13439(x13439, x13438, x13437);
  nand n13440(x13440, x2269, x6139);
  nand n13441(x13441, x7156, x6009);
  nand n13442(x13442, x13441, x13440);
  nand n13443(x13443, x2269, x5879);
  nand n13444(x13444, x7156, x5749);
  nand n13445(x13445, x13444, x13443);
  nand n13446(x13446, x2269, x5619);
  nand n13447(x13447, x7156, x5489);
  nand n13448(x13448, x13447, x13446);
  nand n13449(x13449, x2272, x13439);
  nand n13450(x13450, x7169, x13442);
  nand n13451(x13451, x13450, x13449);
  nand n13452(x13452, x2272, x13445);
  nand n13453(x13453, x7169, x13448);
  nand n13454(x13454, x13453, x13452);
  nand n13455(x13455, x2275, x13451);
  nand n13456(x13456, x7176, x13454);
  nand n13457(x13457, x13456, x13455);
  nand n13458(x13458, x2269, x6403);
  nand n13459(x13459, x7156, x6273);
  nand n13460(x13460, x13459, x13458);
  nand n13461(x13461, x2269, x6143);
  nand n13462(x13462, x7156, x6013);
  nand n13463(x13463, x13462, x13461);
  nand n13464(x13464, x2269, x5883);
  nand n13465(x13465, x7156, x5753);
  nand n13466(x13466, x13465, x13464);
  nand n13467(x13467, x2269, x5623);
  nand n13468(x13468, x7156, x5493);
  nand n13469(x13469, x13468, x13467);
  nand n13470(x13470, x2272, x13460);
  nand n13471(x13471, x7169, x13463);
  nand n13472(x13472, x13471, x13470);
  nand n13473(x13473, x2272, x13466);
  nand n13474(x13474, x7169, x13469);
  nand n13475(x13475, x13474, x13473);
  nand n13476(x13476, x2275, x13472);
  nand n13477(x13477, x7176, x13475);
  nand n13478(x13478, x13477, x13476);
  nand n13479(x13479, x2269, x6407);
  nand n13480(x13480, x7156, x6277);
  nand n13481(x13481, x13480, x13479);
  nand n13482(x13482, x2269, x6147);
  nand n13483(x13483, x7156, x6017);
  nand n13484(x13484, x13483, x13482);
  nand n13485(x13485, x2269, x5887);
  nand n13486(x13486, x7156, x5757);
  nand n13487(x13487, x13486, x13485);
  nand n13488(x13488, x2269, x5627);
  nand n13489(x13489, x7156, x5497);
  nand n13490(x13490, x13489, x13488);
  nand n13491(x13491, x2272, x13481);
  nand n13492(x13492, x7169, x13484);
  nand n13493(x13493, x13492, x13491);
  nand n13494(x13494, x2272, x13487);
  nand n13495(x13495, x7169, x13490);
  nand n13496(x13496, x13495, x13494);
  nand n13497(x13497, x2275, x13493);
  nand n13498(x13498, x7176, x13496);
  nand n13499(x13499, x13498, x13497);
  nand n13500(x13500, x2269, x6411);
  nand n13501(x13501, x7156, x6281);
  nand n13502(x13502, x13501, x13500);
  nand n13503(x13503, x2269, x6151);
  nand n13504(x13504, x7156, x6021);
  nand n13505(x13505, x13504, x13503);
  nand n13506(x13506, x2269, x5891);
  nand n13507(x13507, x7156, x5761);
  nand n13508(x13508, x13507, x13506);
  nand n13509(x13509, x2269, x5631);
  nand n13510(x13510, x7156, x5501);
  nand n13511(x13511, x13510, x13509);
  nand n13512(x13512, x2272, x13502);
  nand n13513(x13513, x7169, x13505);
  nand n13514(x13514, x13513, x13512);
  nand n13515(x13515, x2272, x13508);
  nand n13516(x13516, x7169, x13511);
  nand n13517(x13517, x13516, x13515);
  nand n13518(x13518, x2275, x13514);
  nand n13519(x13519, x7176, x13517);
  nand n13520(x13520, x13519, x13518);
  nand n13521(x13521, x2269, x6415);
  nand n13522(x13522, x7156, x6285);
  nand n13523(x13523, x13522, x13521);
  nand n13524(x13524, x2269, x6155);
  nand n13525(x13525, x7156, x6025);
  nand n13526(x13526, x13525, x13524);
  nand n13527(x13527, x2269, x5895);
  nand n13528(x13528, x7156, x5765);
  nand n13529(x13529, x13528, x13527);
  nand n13530(x13530, x2269, x5635);
  nand n13531(x13531, x7156, x5505);
  nand n13532(x13532, x13531, x13530);
  nand n13533(x13533, x2272, x13523);
  nand n13534(x13534, x7169, x13526);
  nand n13535(x13535, x13534, x13533);
  nand n13536(x13536, x2272, x13529);
  nand n13537(x13537, x7169, x13532);
  nand n13538(x13538, x13537, x13536);
  nand n13539(x13539, x2275, x13535);
  nand n13540(x13540, x7176, x13538);
  nand n13541(x13541, x13540, x13539);
  nand n13542(x13542, x2269, x6419);
  nand n13543(x13543, x7156, x6289);
  nand n13544(x13544, x13543, x13542);
  nand n13545(x13545, x2269, x6159);
  nand n13546(x13546, x7156, x6029);
  nand n13547(x13547, x13546, x13545);
  nand n13548(x13548, x2269, x5899);
  nand n13549(x13549, x7156, x5769);
  nand n13550(x13550, x13549, x13548);
  nand n13551(x13551, x2269, x5639);
  nand n13552(x13552, x7156, x5509);
  nand n13553(x13553, x13552, x13551);
  nand n13554(x13554, x2272, x13544);
  nand n13555(x13555, x7169, x13547);
  nand n13556(x13556, x13555, x13554);
  nand n13557(x13557, x2272, x13550);
  nand n13558(x13558, x7169, x13553);
  nand n13559(x13559, x13558, x13557);
  nand n13560(x13560, x2275, x13556);
  nand n13561(x13561, x7176, x13559);
  nand n13562(x13562, x13561, x13560);
  nand n13563(x13563, x2269, x6423);
  nand n13564(x13564, x7156, x6293);
  nand n13565(x13565, x13564, x13563);
  nand n13566(x13566, x2269, x6163);
  nand n13567(x13567, x7156, x6033);
  nand n13568(x13568, x13567, x13566);
  nand n13569(x13569, x2269, x5903);
  nand n13570(x13570, x7156, x5773);
  nand n13571(x13571, x13570, x13569);
  nand n13572(x13572, x2269, x5643);
  nand n13573(x13573, x7156, x5513);
  nand n13574(x13574, x13573, x13572);
  nand n13575(x13575, x2272, x13565);
  nand n13576(x13576, x7169, x13568);
  nand n13577(x13577, x13576, x13575);
  nand n13578(x13578, x2272, x13571);
  nand n13579(x13579, x7169, x13574);
  nand n13580(x13580, x13579, x13578);
  nand n13581(x13581, x2275, x13577);
  nand n13582(x13582, x7176, x13580);
  nand n13583(x13583, x13582, x13581);
  nand n13584(x13584, x2269, x6427);
  nand n13585(x13585, x7156, x6297);
  nand n13586(x13586, x13585, x13584);
  nand n13587(x13587, x2269, x6167);
  nand n13588(x13588, x7156, x6037);
  nand n13589(x13589, x13588, x13587);
  nand n13590(x13590, x2269, x5907);
  nand n13591(x13591, x7156, x5777);
  nand n13592(x13592, x13591, x13590);
  nand n13593(x13593, x2269, x5647);
  nand n13594(x13594, x7156, x5517);
  nand n13595(x13595, x13594, x13593);
  nand n13596(x13596, x2272, x13586);
  nand n13597(x13597, x7169, x13589);
  nand n13598(x13598, x13597, x13596);
  nand n13599(x13599, x2272, x13592);
  nand n13600(x13600, x7169, x13595);
  nand n13601(x13601, x13600, x13599);
  nand n13602(x13602, x2275, x13598);
  nand n13603(x13603, x7176, x13601);
  nand n13604(x13604, x13603, x13602);
  nand n13605(x13605, x2269, x6431);
  nand n13606(x13606, x7156, x6301);
  nand n13607(x13607, x13606, x13605);
  nand n13608(x13608, x2269, x6171);
  nand n13609(x13609, x7156, x6041);
  nand n13610(x13610, x13609, x13608);
  nand n13611(x13611, x2269, x5911);
  nand n13612(x13612, x7156, x5781);
  nand n13613(x13613, x13612, x13611);
  nand n13614(x13614, x2269, x5651);
  nand n13615(x13615, x7156, x5521);
  nand n13616(x13616, x13615, x13614);
  nand n13617(x13617, x2272, x13607);
  nand n13618(x13618, x7169, x13610);
  nand n13619(x13619, x13618, x13617);
  nand n13620(x13620, x2272, x13613);
  nand n13621(x13621, x7169, x13616);
  nand n13622(x13622, x13621, x13620);
  nand n13623(x13623, x2275, x13619);
  nand n13624(x13624, x7176, x13622);
  nand n13625(x13625, x13624, x13623);
  nand n13626(x13626, x2269, x6435);
  nand n13627(x13627, x7156, x6305);
  nand n13628(x13628, x13627, x13626);
  nand n13629(x13629, x2269, x6175);
  nand n13630(x13630, x7156, x6045);
  nand n13631(x13631, x13630, x13629);
  nand n13632(x13632, x2269, x5915);
  nand n13633(x13633, x7156, x5785);
  nand n13634(x13634, x13633, x13632);
  nand n13635(x13635, x2269, x5655);
  nand n13636(x13636, x7156, x5525);
  nand n13637(x13637, x13636, x13635);
  nand n13638(x13638, x2272, x13628);
  nand n13639(x13639, x7169, x13631);
  nand n13640(x13640, x13639, x13638);
  nand n13641(x13641, x2272, x13634);
  nand n13642(x13642, x7169, x13637);
  nand n13643(x13643, x13642, x13641);
  nand n13644(x13644, x2275, x13640);
  nand n13645(x13645, x7176, x13643);
  nand n13646(x13646, x13645, x13644);
  nand n13647(x13647, x2269, x6439);
  nand n13648(x13648, x7156, x6309);
  nand n13649(x13649, x13648, x13647);
  nand n13650(x13650, x2269, x6179);
  nand n13651(x13651, x7156, x6049);
  nand n13652(x13652, x13651, x13650);
  nand n13653(x13653, x2269, x5919);
  nand n13654(x13654, x7156, x5789);
  nand n13655(x13655, x13654, x13653);
  nand n13656(x13656, x2269, x5659);
  nand n13657(x13657, x7156, x5529);
  nand n13658(x13658, x13657, x13656);
  nand n13659(x13659, x2272, x13649);
  nand n13660(x13660, x7169, x13652);
  nand n13661(x13661, x13660, x13659);
  nand n13662(x13662, x2272, x13655);
  nand n13663(x13663, x7169, x13658);
  nand n13664(x13664, x13663, x13662);
  nand n13665(x13665, x2275, x13661);
  nand n13666(x13666, x7176, x13664);
  nand n13667(x13667, x13666, x13665);
  nand n13668(x13668, x2269, x6443);
  nand n13669(x13669, x7156, x6313);
  nand n13670(x13670, x13669, x13668);
  nand n13671(x13671, x2269, x6183);
  nand n13672(x13672, x7156, x6053);
  nand n13673(x13673, x13672, x13671);
  nand n13674(x13674, x2269, x5923);
  nand n13675(x13675, x7156, x5793);
  nand n13676(x13676, x13675, x13674);
  nand n13677(x13677, x2269, x5663);
  nand n13678(x13678, x7156, x5533);
  nand n13679(x13679, x13678, x13677);
  nand n13680(x13680, x2272, x13670);
  nand n13681(x13681, x7169, x13673);
  nand n13682(x13682, x13681, x13680);
  nand n13683(x13683, x2272, x13676);
  nand n13684(x13684, x7169, x13679);
  nand n13685(x13685, x13684, x13683);
  nand n13686(x13686, x2275, x13682);
  nand n13687(x13687, x7176, x13685);
  nand n13688(x13688, x13687, x13686);
  nand n13689(x13689, x2269, x6447);
  nand n13690(x13690, x7156, x6317);
  nand n13691(x13691, x13690, x13689);
  nand n13692(x13692, x2269, x6187);
  nand n13693(x13693, x7156, x6057);
  nand n13694(x13694, x13693, x13692);
  nand n13695(x13695, x2269, x5927);
  nand n13696(x13696, x7156, x5797);
  nand n13697(x13697, x13696, x13695);
  nand n13698(x13698, x2269, x5667);
  nand n13699(x13699, x7156, x5537);
  nand n13700(x13700, x13699, x13698);
  nand n13701(x13701, x2272, x13691);
  nand n13702(x13702, x7169, x13694);
  nand n13703(x13703, x13702, x13701);
  nand n13704(x13704, x2272, x13697);
  nand n13705(x13705, x7169, x13700);
  nand n13706(x13706, x13705, x13704);
  nand n13707(x13707, x2275, x13703);
  nand n13708(x13708, x7176, x13706);
  nand n13709(x13709, x13708, x13707);
  nand n13710(x13710, x2269, x6451);
  nand n13711(x13711, x7156, x6321);
  nand n13712(x13712, x13711, x13710);
  nand n13713(x13713, x2269, x6191);
  nand n13714(x13714, x7156, x6061);
  nand n13715(x13715, x13714, x13713);
  nand n13716(x13716, x2269, x5931);
  nand n13717(x13717, x7156, x5801);
  nand n13718(x13718, x13717, x13716);
  nand n13719(x13719, x2269, x5671);
  nand n13720(x13720, x7156, x5541);
  nand n13721(x13721, x13720, x13719);
  nand n13722(x13722, x2272, x13712);
  nand n13723(x13723, x7169, x13715);
  nand n13724(x13724, x13723, x13722);
  nand n13725(x13725, x2272, x13718);
  nand n13726(x13726, x7169, x13721);
  nand n13727(x13727, x13726, x13725);
  nand n13728(x13728, x2275, x13724);
  nand n13729(x13729, x7176, x13727);
  nand n13730(x13730, x13729, x13728);
  nand n13731(x13731, x2269, x6455);
  nand n13732(x13732, x7156, x6325);
  nand n13733(x13733, x13732, x13731);
  nand n13734(x13734, x2269, x6195);
  nand n13735(x13735, x7156, x6065);
  nand n13736(x13736, x13735, x13734);
  nand n13737(x13737, x2269, x5935);
  nand n13738(x13738, x7156, x5805);
  nand n13739(x13739, x13738, x13737);
  nand n13740(x13740, x2269, x5675);
  nand n13741(x13741, x7156, x5545);
  nand n13742(x13742, x13741, x13740);
  nand n13743(x13743, x2272, x13733);
  nand n13744(x13744, x7169, x13736);
  nand n13745(x13745, x13744, x13743);
  nand n13746(x13746, x2272, x13739);
  nand n13747(x13747, x7169, x13742);
  nand n13748(x13748, x13747, x13746);
  nand n13749(x13749, x2275, x13745);
  nand n13750(x13750, x7176, x13748);
  nand n13751(x13751, x13750, x13749);
  nand n13752(x13752, x2269, x6459);
  nand n13753(x13753, x7156, x6329);
  nand n13754(x13754, x13753, x13752);
  nand n13755(x13755, x2269, x6199);
  nand n13756(x13756, x7156, x6069);
  nand n13757(x13757, x13756, x13755);
  nand n13758(x13758, x2269, x5939);
  nand n13759(x13759, x7156, x5809);
  nand n13760(x13760, x13759, x13758);
  nand n13761(x13761, x2269, x5679);
  nand n13762(x13762, x7156, x5549);
  nand n13763(x13763, x13762, x13761);
  nand n13764(x13764, x2272, x13754);
  nand n13765(x13765, x7169, x13757);
  nand n13766(x13766, x13765, x13764);
  nand n13767(x13767, x2272, x13760);
  nand n13768(x13768, x7169, x13763);
  nand n13769(x13769, x13768, x13767);
  nand n13770(x13770, x2275, x13766);
  nand n13771(x13771, x7176, x13769);
  nand n13772(x13772, x13771, x13770);
  nand n13773(x13773, x2269, x6463);
  nand n13774(x13774, x7156, x6333);
  nand n13775(x13775, x13774, x13773);
  nand n13776(x13776, x2269, x6203);
  nand n13777(x13777, x7156, x6073);
  nand n13778(x13778, x13777, x13776);
  nand n13779(x13779, x2269, x5943);
  nand n13780(x13780, x7156, x5813);
  nand n13781(x13781, x13780, x13779);
  nand n13782(x13782, x2269, x5683);
  nand n13783(x13783, x7156, x5553);
  nand n13784(x13784, x13783, x13782);
  nand n13785(x13785, x2272, x13775);
  nand n13786(x13786, x7169, x13778);
  nand n13787(x13787, x13786, x13785);
  nand n13788(x13788, x2272, x13781);
  nand n13789(x13789, x7169, x13784);
  nand n13790(x13790, x13789, x13788);
  nand n13791(x13791, x2275, x13787);
  nand n13792(x13792, x7176, x13790);
  nand n13793(x13793, x13792, x13791);
  nand n13794(x13794, x2269, x6467);
  nand n13795(x13795, x7156, x6337);
  nand n13796(x13796, x13795, x13794);
  nand n13797(x13797, x2269, x6207);
  nand n13798(x13798, x7156, x6077);
  nand n13799(x13799, x13798, x13797);
  nand n13800(x13800, x2269, x5947);
  nand n13801(x13801, x7156, x5817);
  nand n13802(x13802, x13801, x13800);
  nand n13803(x13803, x2269, x5687);
  nand n13804(x13804, x7156, x5557);
  nand n13805(x13805, x13804, x13803);
  nand n13806(x13806, x2272, x13796);
  nand n13807(x13807, x7169, x13799);
  nand n13808(x13808, x13807, x13806);
  nand n13809(x13809, x2272, x13802);
  nand n13810(x13810, x7169, x13805);
  nand n13811(x13811, x13810, x13809);
  nand n13812(x13812, x2275, x13808);
  nand n13813(x13813, x7176, x13811);
  nand n13814(x13814, x13813, x13812);
  nand n13815(x13815, x2269, x6471);
  nand n13816(x13816, x7156, x6341);
  nand n13817(x13817, x13816, x13815);
  nand n13818(x13818, x2269, x6211);
  nand n13819(x13819, x7156, x6081);
  nand n13820(x13820, x13819, x13818);
  nand n13821(x13821, x2269, x5951);
  nand n13822(x13822, x7156, x5821);
  nand n13823(x13823, x13822, x13821);
  nand n13824(x13824, x2269, x5691);
  nand n13825(x13825, x7156, x5561);
  nand n13826(x13826, x13825, x13824);
  nand n13827(x13827, x2272, x13817);
  nand n13828(x13828, x7169, x13820);
  nand n13829(x13829, x13828, x13827);
  nand n13830(x13830, x2272, x13823);
  nand n13831(x13831, x7169, x13826);
  nand n13832(x13832, x13831, x13830);
  nand n13833(x13833, x2275, x13829);
  nand n13834(x13834, x7176, x13832);
  nand n13835(x13835, x13834, x13833);
  nand n13836(x13836, x2269, x6475);
  nand n13837(x13837, x7156, x6345);
  nand n13838(x13838, x13837, x13836);
  nand n13839(x13839, x2269, x6215);
  nand n13840(x13840, x7156, x6085);
  nand n13841(x13841, x13840, x13839);
  nand n13842(x13842, x2269, x5955);
  nand n13843(x13843, x7156, x5825);
  nand n13844(x13844, x13843, x13842);
  nand n13845(x13845, x2269, x5695);
  nand n13846(x13846, x7156, x5565);
  nand n13847(x13847, x13846, x13845);
  nand n13848(x13848, x2272, x13838);
  nand n13849(x13849, x7169, x13841);
  nand n13850(x13850, x13849, x13848);
  nand n13851(x13851, x2272, x13844);
  nand n13852(x13852, x7169, x13847);
  nand n13853(x13853, x13852, x13851);
  nand n13854(x13854, x2275, x13850);
  nand n13855(x13855, x7176, x13853);
  nand n13856(x13856, x13855, x13854);
  nand n13857(x13857, x2269, x6479);
  nand n13858(x13858, x7156, x6349);
  nand n13859(x13859, x13858, x13857);
  nand n13860(x13860, x2269, x6219);
  nand n13861(x13861, x7156, x6089);
  nand n13862(x13862, x13861, x13860);
  nand n13863(x13863, x2269, x5959);
  nand n13864(x13864, x7156, x5829);
  nand n13865(x13865, x13864, x13863);
  nand n13866(x13866, x2269, x5699);
  nand n13867(x13867, x7156, x5569);
  nand n13868(x13868, x13867, x13866);
  nand n13869(x13869, x2272, x13859);
  nand n13870(x13870, x7169, x13862);
  nand n13871(x13871, x13870, x13869);
  nand n13872(x13872, x2272, x13865);
  nand n13873(x13873, x7169, x13868);
  nand n13874(x13874, x13873, x13872);
  nand n13875(x13875, x2275, x13871);
  nand n13876(x13876, x7176, x13874);
  nand n13877(x13877, x13876, x13875);
  nand n13878(x13878, x71202, x6355);
  nand n13879(x13879, x1448, x6225);
  nand n13880(x13880, x13879, x13878);
  nand n13881(x13881, x71202, x6095);
  nand n13882(x13882, x1448, x5965);
  nand n13883(x13883, x13882, x13881);
  nand n13884(x13884, x71202, x5835);
  nand n13885(x13885, x1448, x5705);
  nand n13886(x13886, x13885, x13884);
  nand n13887(x13887, x71202, x5575);
  nand n13888(x13888, x1448, x5443);
  nand n13889(x13889, x13888, x13887);
  nand n13890(x13890, x71205, x13880);
  nand n13891(x13891, x1461, x13883);
  nand n13892(x13892, x13891, x13890);
  nand n13893(x13893, x71205, x13886);
  nand n13894(x13894, x1461, x13889);
  nand n13895(x13895, x13894, x13893);
  nand n13896(x13896, x71210, x13892);
  nand n13897(x13897, x1468, x13895);
  nand n13898(x13898, x13897, x13896);
  nand n13899(x13899, x71202, x6359);
  nand n13900(x13900, x1448, x6229);
  nand n13901(x13901, x13900, x13899);
  nand n13902(x13902, x71202, x6099);
  nand n13903(x13903, x1448, x5969);
  nand n13904(x13904, x13903, x13902);
  nand n13905(x13905, x71202, x5839);
  nand n13906(x13906, x1448, x5709);
  nand n13907(x13907, x13906, x13905);
  nand n13908(x13908, x71202, x5579);
  nand n13909(x13909, x1448, x5449);
  nand n13910(x13910, x13909, x13908);
  nand n13911(x13911, x71205, x13901);
  nand n13912(x13912, x1461, x13904);
  nand n13913(x13913, x13912, x13911);
  nand n13914(x13914, x71205, x13907);
  nand n13915(x13915, x1461, x13910);
  nand n13916(x13916, x13915, x13914);
  nand n13917(x13917, x71210, x13913);
  nand n13918(x13918, x1468, x13916);
  nand n13919(x13919, x13918, x13917);
  nand n13920(x13920, x71202, x6363);
  nand n13921(x13921, x1448, x6233);
  nand n13922(x13922, x13921, x13920);
  nand n13923(x13923, x71202, x6103);
  nand n13924(x13924, x1448, x5973);
  nand n13925(x13925, x13924, x13923);
  nand n13926(x13926, x71202, x5843);
  nand n13927(x13927, x1448, x5713);
  nand n13928(x13928, x13927, x13926);
  nand n13929(x13929, x71202, x5583);
  nand n13930(x13930, x1448, x5453);
  nand n13931(x13931, x13930, x13929);
  nand n13932(x13932, x71205, x13922);
  nand n13933(x13933, x1461, x13925);
  nand n13934(x13934, x13933, x13932);
  nand n13935(x13935, x71205, x13928);
  nand n13936(x13936, x1461, x13931);
  nand n13937(x13937, x13936, x13935);
  nand n13938(x13938, x71210, x13934);
  nand n13939(x13939, x1468, x13937);
  nand n13940(x13940, x13939, x13938);
  nand n13941(x13941, x71202, x6367);
  nand n13942(x13942, x1448, x6237);
  nand n13943(x13943, x13942, x13941);
  nand n13944(x13944, x71202, x6107);
  nand n13945(x13945, x1448, x5977);
  nand n13946(x13946, x13945, x13944);
  nand n13947(x13947, x71202, x5847);
  nand n13948(x13948, x1448, x5717);
  nand n13949(x13949, x13948, x13947);
  nand n13950(x13950, x71202, x5587);
  nand n13951(x13951, x1448, x5457);
  nand n13952(x13952, x13951, x13950);
  nand n13953(x13953, x71205, x13943);
  nand n13954(x13954, x1461, x13946);
  nand n13955(x13955, x13954, x13953);
  nand n13956(x13956, x71205, x13949);
  nand n13957(x13957, x1461, x13952);
  nand n13958(x13958, x13957, x13956);
  nand n13959(x13959, x71210, x13955);
  nand n13960(x13960, x1468, x13958);
  nand n13961(x13961, x13960, x13959);
  nand n13962(x13962, x71202, x6371);
  nand n13963(x13963, x1448, x6241);
  nand n13964(x13964, x13963, x13962);
  nand n13965(x13965, x71202, x6111);
  nand n13966(x13966, x1448, x5981);
  nand n13967(x13967, x13966, x13965);
  nand n13968(x13968, x71202, x5851);
  nand n13969(x13969, x1448, x5721);
  nand n13970(x13970, x13969, x13968);
  nand n13971(x13971, x71202, x5591);
  nand n13972(x13972, x1448, x5461);
  nand n13973(x13973, x13972, x13971);
  nand n13974(x13974, x71205, x13964);
  nand n13975(x13975, x1461, x13967);
  nand n13976(x13976, x13975, x13974);
  nand n13977(x13977, x71205, x13970);
  nand n13978(x13978, x1461, x13973);
  nand n13979(x13979, x13978, x13977);
  nand n13980(x13980, x71210, x13976);
  nand n13981(x13981, x1468, x13979);
  nand n13982(x13982, x13981, x13980);
  nand n13983(x13983, x71202, x6375);
  nand n13984(x13984, x1448, x6245);
  nand n13985(x13985, x13984, x13983);
  nand n13986(x13986, x71202, x6115);
  nand n13987(x13987, x1448, x5985);
  nand n13988(x13988, x13987, x13986);
  nand n13989(x13989, x71202, x5855);
  nand n13990(x13990, x1448, x5725);
  nand n13991(x13991, x13990, x13989);
  nand n13992(x13992, x71202, x5595);
  nand n13993(x13993, x1448, x5465);
  nand n13994(x13994, x13993, x13992);
  nand n13995(x13995, x71205, x13985);
  nand n13996(x13996, x1461, x13988);
  nand n13997(x13997, x13996, x13995);
  nand n13998(x13998, x71205, x13991);
  nand n13999(x13999, x1461, x13994);
  nand n14000(x14000, x13999, x13998);
  nand n14001(x14001, x71210, x13997);
  nand n14002(x14002, x1468, x14000);
  nand n14003(x14003, x14002, x14001);
  nand n14004(x14004, x71202, x6379);
  nand n14005(x14005, x1448, x6249);
  nand n14006(x14006, x14005, x14004);
  nand n14007(x14007, x71202, x6119);
  nand n14008(x14008, x1448, x5989);
  nand n14009(x14009, x14008, x14007);
  nand n14010(x14010, x71202, x5859);
  nand n14011(x14011, x1448, x5729);
  nand n14012(x14012, x14011, x14010);
  nand n14013(x14013, x71202, x5599);
  nand n14014(x14014, x1448, x5469);
  nand n14015(x14015, x14014, x14013);
  nand n14016(x14016, x71205, x14006);
  nand n14017(x14017, x1461, x14009);
  nand n14018(x14018, x14017, x14016);
  nand n14019(x14019, x71205, x14012);
  nand n14020(x14020, x1461, x14015);
  nand n14021(x14021, x14020, x14019);
  nand n14022(x14022, x71210, x14018);
  nand n14023(x14023, x1468, x14021);
  nand n14024(x14024, x14023, x14022);
  nand n14025(x14025, x71202, x6383);
  nand n14026(x14026, x1448, x6253);
  nand n14027(x14027, x14026, x14025);
  nand n14028(x14028, x71202, x6123);
  nand n14029(x14029, x1448, x5993);
  nand n14030(x14030, x14029, x14028);
  nand n14031(x14031, x71202, x5863);
  nand n14032(x14032, x1448, x5733);
  nand n14033(x14033, x14032, x14031);
  nand n14034(x14034, x71202, x5603);
  nand n14035(x14035, x1448, x5473);
  nand n14036(x14036, x14035, x14034);
  nand n14037(x14037, x71205, x14027);
  nand n14038(x14038, x1461, x14030);
  nand n14039(x14039, x14038, x14037);
  nand n14040(x14040, x71205, x14033);
  nand n14041(x14041, x1461, x14036);
  nand n14042(x14042, x14041, x14040);
  nand n14043(x14043, x71210, x14039);
  nand n14044(x14044, x1468, x14042);
  nand n14045(x14045, x14044, x14043);
  nand n14046(x14046, x71202, x6387);
  nand n14047(x14047, x1448, x6257);
  nand n14048(x14048, x14047, x14046);
  nand n14049(x14049, x71202, x6127);
  nand n14050(x14050, x1448, x5997);
  nand n14051(x14051, x14050, x14049);
  nand n14052(x14052, x71202, x5867);
  nand n14053(x14053, x1448, x5737);
  nand n14054(x14054, x14053, x14052);
  nand n14055(x14055, x71202, x5607);
  nand n14056(x14056, x1448, x5477);
  nand n14057(x14057, x14056, x14055);
  nand n14058(x14058, x71205, x14048);
  nand n14059(x14059, x1461, x14051);
  nand n14060(x14060, x14059, x14058);
  nand n14061(x14061, x71205, x14054);
  nand n14062(x14062, x1461, x14057);
  nand n14063(x14063, x14062, x14061);
  nand n14064(x14064, x71210, x14060);
  nand n14065(x14065, x1468, x14063);
  nand n14066(x14066, x14065, x14064);
  nand n14067(x14067, x71202, x6391);
  nand n14068(x14068, x1448, x6261);
  nand n14069(x14069, x14068, x14067);
  nand n14070(x14070, x71202, x6131);
  nand n14071(x14071, x1448, x6001);
  nand n14072(x14072, x14071, x14070);
  nand n14073(x14073, x71202, x5871);
  nand n14074(x14074, x1448, x5741);
  nand n14075(x14075, x14074, x14073);
  nand n14076(x14076, x71202, x5611);
  nand n14077(x14077, x1448, x5481);
  nand n14078(x14078, x14077, x14076);
  nand n14079(x14079, x71205, x14069);
  nand n14080(x14080, x1461, x14072);
  nand n14081(x14081, x14080, x14079);
  nand n14082(x14082, x71205, x14075);
  nand n14083(x14083, x1461, x14078);
  nand n14084(x14084, x14083, x14082);
  nand n14085(x14085, x71210, x14081);
  nand n14086(x14086, x1468, x14084);
  nand n14087(x14087, x14086, x14085);
  nand n14088(x14088, x71202, x6395);
  nand n14089(x14089, x1448, x6265);
  nand n14090(x14090, x14089, x14088);
  nand n14091(x14091, x71202, x6135);
  nand n14092(x14092, x1448, x6005);
  nand n14093(x14093, x14092, x14091);
  nand n14094(x14094, x71202, x5875);
  nand n14095(x14095, x1448, x5745);
  nand n14096(x14096, x14095, x14094);
  nand n14097(x14097, x71202, x5615);
  nand n14098(x14098, x1448, x5485);
  nand n14099(x14099, x14098, x14097);
  nand n14100(x14100, x71205, x14090);
  nand n14101(x14101, x1461, x14093);
  nand n14102(x14102, x14101, x14100);
  nand n14103(x14103, x71205, x14096);
  nand n14104(x14104, x1461, x14099);
  nand n14105(x14105, x14104, x14103);
  nand n14106(x14106, x71210, x14102);
  nand n14107(x14107, x1468, x14105);
  nand n14108(x14108, x14107, x14106);
  nand n14109(x14109, x71202, x6399);
  nand n14110(x14110, x1448, x6269);
  nand n14111(x14111, x14110, x14109);
  nand n14112(x14112, x71202, x6139);
  nand n14113(x14113, x1448, x6009);
  nand n14114(x14114, x14113, x14112);
  nand n14115(x14115, x71202, x5879);
  nand n14116(x14116, x1448, x5749);
  nand n14117(x14117, x14116, x14115);
  nand n14118(x14118, x71202, x5619);
  nand n14119(x14119, x1448, x5489);
  nand n14120(x14120, x14119, x14118);
  nand n14121(x14121, x71205, x14111);
  nand n14122(x14122, x1461, x14114);
  nand n14123(x14123, x14122, x14121);
  nand n14124(x14124, x71205, x14117);
  nand n14125(x14125, x1461, x14120);
  nand n14126(x14126, x14125, x14124);
  nand n14127(x14127, x71210, x14123);
  nand n14128(x14128, x1468, x14126);
  nand n14129(x14129, x14128, x14127);
  nand n14130(x14130, x71202, x6403);
  nand n14131(x14131, x1448, x6273);
  nand n14132(x14132, x14131, x14130);
  nand n14133(x14133, x71202, x6143);
  nand n14134(x14134, x1448, x6013);
  nand n14135(x14135, x14134, x14133);
  nand n14136(x14136, x71202, x5883);
  nand n14137(x14137, x1448, x5753);
  nand n14138(x14138, x14137, x14136);
  nand n14139(x14139, x71202, x5623);
  nand n14140(x14140, x1448, x5493);
  nand n14141(x14141, x14140, x14139);
  nand n14142(x14142, x71205, x14132);
  nand n14143(x14143, x1461, x14135);
  nand n14144(x14144, x14143, x14142);
  nand n14145(x14145, x71205, x14138);
  nand n14146(x14146, x1461, x14141);
  nand n14147(x14147, x14146, x14145);
  nand n14148(x14148, x71210, x14144);
  nand n14149(x14149, x1468, x14147);
  nand n14150(x14150, x14149, x14148);
  nand n14151(x14151, x71202, x6407);
  nand n14152(x14152, x1448, x6277);
  nand n14153(x14153, x14152, x14151);
  nand n14154(x14154, x71202, x6147);
  nand n14155(x14155, x1448, x6017);
  nand n14156(x14156, x14155, x14154);
  nand n14157(x14157, x71202, x5887);
  nand n14158(x14158, x1448, x5757);
  nand n14159(x14159, x14158, x14157);
  nand n14160(x14160, x71202, x5627);
  nand n14161(x14161, x1448, x5497);
  nand n14162(x14162, x14161, x14160);
  nand n14163(x14163, x71205, x14153);
  nand n14164(x14164, x1461, x14156);
  nand n14165(x14165, x14164, x14163);
  nand n14166(x14166, x71205, x14159);
  nand n14167(x14167, x1461, x14162);
  nand n14168(x14168, x14167, x14166);
  nand n14169(x14169, x71210, x14165);
  nand n14170(x14170, x1468, x14168);
  nand n14171(x14171, x14170, x14169);
  nand n14172(x14172, x71202, x6411);
  nand n14173(x14173, x1448, x6281);
  nand n14174(x14174, x14173, x14172);
  nand n14175(x14175, x71202, x6151);
  nand n14176(x14176, x1448, x6021);
  nand n14177(x14177, x14176, x14175);
  nand n14178(x14178, x71202, x5891);
  nand n14179(x14179, x1448, x5761);
  nand n14180(x14180, x14179, x14178);
  nand n14181(x14181, x71202, x5631);
  nand n14182(x14182, x1448, x5501);
  nand n14183(x14183, x14182, x14181);
  nand n14184(x14184, x71205, x14174);
  nand n14185(x14185, x1461, x14177);
  nand n14186(x14186, x14185, x14184);
  nand n14187(x14187, x71205, x14180);
  nand n14188(x14188, x1461, x14183);
  nand n14189(x14189, x14188, x14187);
  nand n14190(x14190, x71210, x14186);
  nand n14191(x14191, x1468, x14189);
  nand n14192(x14192, x14191, x14190);
  nand n14193(x14193, x71202, x6415);
  nand n14194(x14194, x1448, x6285);
  nand n14195(x14195, x14194, x14193);
  nand n14196(x14196, x71202, x6155);
  nand n14197(x14197, x1448, x6025);
  nand n14198(x14198, x14197, x14196);
  nand n14199(x14199, x71202, x5895);
  nand n14200(x14200, x1448, x5765);
  nand n14201(x14201, x14200, x14199);
  nand n14202(x14202, x71202, x5635);
  nand n14203(x14203, x1448, x5505);
  nand n14204(x14204, x14203, x14202);
  nand n14205(x14205, x71205, x14195);
  nand n14206(x14206, x1461, x14198);
  nand n14207(x14207, x14206, x14205);
  nand n14208(x14208, x71205, x14201);
  nand n14209(x14209, x1461, x14204);
  nand n14210(x14210, x14209, x14208);
  nand n14211(x14211, x71210, x14207);
  nand n14212(x14212, x1468, x14210);
  nand n14213(x14213, x14212, x14211);
  nand n14214(x14214, x71202, x6419);
  nand n14215(x14215, x1448, x6289);
  nand n14216(x14216, x14215, x14214);
  nand n14217(x14217, x71202, x6159);
  nand n14218(x14218, x1448, x6029);
  nand n14219(x14219, x14218, x14217);
  nand n14220(x14220, x71202, x5899);
  nand n14221(x14221, x1448, x5769);
  nand n14222(x14222, x14221, x14220);
  nand n14223(x14223, x71202, x5639);
  nand n14224(x14224, x1448, x5509);
  nand n14225(x14225, x14224, x14223);
  nand n14226(x14226, x71205, x14216);
  nand n14227(x14227, x1461, x14219);
  nand n14228(x14228, x14227, x14226);
  nand n14229(x14229, x71205, x14222);
  nand n14230(x14230, x1461, x14225);
  nand n14231(x14231, x14230, x14229);
  nand n14232(x14232, x71210, x14228);
  nand n14233(x14233, x1468, x14231);
  nand n14234(x14234, x14233, x14232);
  nand n14235(x14235, x71202, x6423);
  nand n14236(x14236, x1448, x6293);
  nand n14237(x14237, x14236, x14235);
  nand n14238(x14238, x71202, x6163);
  nand n14239(x14239, x1448, x6033);
  nand n14240(x14240, x14239, x14238);
  nand n14241(x14241, x71202, x5903);
  nand n14242(x14242, x1448, x5773);
  nand n14243(x14243, x14242, x14241);
  nand n14244(x14244, x71202, x5643);
  nand n14245(x14245, x1448, x5513);
  nand n14246(x14246, x14245, x14244);
  nand n14247(x14247, x71205, x14237);
  nand n14248(x14248, x1461, x14240);
  nand n14249(x14249, x14248, x14247);
  nand n14250(x14250, x71205, x14243);
  nand n14251(x14251, x1461, x14246);
  nand n14252(x14252, x14251, x14250);
  nand n14253(x14253, x71210, x14249);
  nand n14254(x14254, x1468, x14252);
  nand n14255(x14255, x14254, x14253);
  nand n14256(x14256, x71202, x6427);
  nand n14257(x14257, x1448, x6297);
  nand n14258(x14258, x14257, x14256);
  nand n14259(x14259, x71202, x6167);
  nand n14260(x14260, x1448, x6037);
  nand n14261(x14261, x14260, x14259);
  nand n14262(x14262, x71202, x5907);
  nand n14263(x14263, x1448, x5777);
  nand n14264(x14264, x14263, x14262);
  nand n14265(x14265, x71202, x5647);
  nand n14266(x14266, x1448, x5517);
  nand n14267(x14267, x14266, x14265);
  nand n14268(x14268, x71205, x14258);
  nand n14269(x14269, x1461, x14261);
  nand n14270(x14270, x14269, x14268);
  nand n14271(x14271, x71205, x14264);
  nand n14272(x14272, x1461, x14267);
  nand n14273(x14273, x14272, x14271);
  nand n14274(x14274, x71210, x14270);
  nand n14275(x14275, x1468, x14273);
  nand n14276(x14276, x14275, x14274);
  nand n14277(x14277, x71202, x6431);
  nand n14278(x14278, x1448, x6301);
  nand n14279(x14279, x14278, x14277);
  nand n14280(x14280, x71202, x6171);
  nand n14281(x14281, x1448, x6041);
  nand n14282(x14282, x14281, x14280);
  nand n14283(x14283, x71202, x5911);
  nand n14284(x14284, x1448, x5781);
  nand n14285(x14285, x14284, x14283);
  nand n14286(x14286, x71202, x5651);
  nand n14287(x14287, x1448, x5521);
  nand n14288(x14288, x14287, x14286);
  nand n14289(x14289, x71205, x14279);
  nand n14290(x14290, x1461, x14282);
  nand n14291(x14291, x14290, x14289);
  nand n14292(x14292, x71205, x14285);
  nand n14293(x14293, x1461, x14288);
  nand n14294(x14294, x14293, x14292);
  nand n14295(x14295, x71210, x14291);
  nand n14296(x14296, x1468, x14294);
  nand n14297(x14297, x14296, x14295);
  nand n14298(x14298, x71202, x6435);
  nand n14299(x14299, x1448, x6305);
  nand n14300(x14300, x14299, x14298);
  nand n14301(x14301, x71202, x6175);
  nand n14302(x14302, x1448, x6045);
  nand n14303(x14303, x14302, x14301);
  nand n14304(x14304, x71202, x5915);
  nand n14305(x14305, x1448, x5785);
  nand n14306(x14306, x14305, x14304);
  nand n14307(x14307, x71202, x5655);
  nand n14308(x14308, x1448, x5525);
  nand n14309(x14309, x14308, x14307);
  nand n14310(x14310, x71205, x14300);
  nand n14311(x14311, x1461, x14303);
  nand n14312(x14312, x14311, x14310);
  nand n14313(x14313, x71205, x14306);
  nand n14314(x14314, x1461, x14309);
  nand n14315(x14315, x14314, x14313);
  nand n14316(x14316, x71210, x14312);
  nand n14317(x14317, x1468, x14315);
  nand n14318(x14318, x14317, x14316);
  nand n14319(x14319, x71202, x6439);
  nand n14320(x14320, x1448, x6309);
  nand n14321(x14321, x14320, x14319);
  nand n14322(x14322, x71202, x6179);
  nand n14323(x14323, x1448, x6049);
  nand n14324(x14324, x14323, x14322);
  nand n14325(x14325, x71202, x5919);
  nand n14326(x14326, x1448, x5789);
  nand n14327(x14327, x14326, x14325);
  nand n14328(x14328, x71202, x5659);
  nand n14329(x14329, x1448, x5529);
  nand n14330(x14330, x14329, x14328);
  nand n14331(x14331, x71205, x14321);
  nand n14332(x14332, x1461, x14324);
  nand n14333(x14333, x14332, x14331);
  nand n14334(x14334, x71205, x14327);
  nand n14335(x14335, x1461, x14330);
  nand n14336(x14336, x14335, x14334);
  nand n14337(x14337, x71210, x14333);
  nand n14338(x14338, x1468, x14336);
  nand n14339(x14339, x14338, x14337);
  nand n14340(x14340, x71202, x6443);
  nand n14341(x14341, x1448, x6313);
  nand n14342(x14342, x14341, x14340);
  nand n14343(x14343, x71202, x6183);
  nand n14344(x14344, x1448, x6053);
  nand n14345(x14345, x14344, x14343);
  nand n14346(x14346, x71202, x5923);
  nand n14347(x14347, x1448, x5793);
  nand n14348(x14348, x14347, x14346);
  nand n14349(x14349, x71202, x5663);
  nand n14350(x14350, x1448, x5533);
  nand n14351(x14351, x14350, x14349);
  nand n14352(x14352, x71205, x14342);
  nand n14353(x14353, x1461, x14345);
  nand n14354(x14354, x14353, x14352);
  nand n14355(x14355, x71205, x14348);
  nand n14356(x14356, x1461, x14351);
  nand n14357(x14357, x14356, x14355);
  nand n14358(x14358, x71210, x14354);
  nand n14359(x14359, x1468, x14357);
  nand n14360(x14360, x14359, x14358);
  nand n14361(x14361, x71202, x6447);
  nand n14362(x14362, x1448, x6317);
  nand n14363(x14363, x14362, x14361);
  nand n14364(x14364, x71202, x6187);
  nand n14365(x14365, x1448, x6057);
  nand n14366(x14366, x14365, x14364);
  nand n14367(x14367, x71202, x5927);
  nand n14368(x14368, x1448, x5797);
  nand n14369(x14369, x14368, x14367);
  nand n14370(x14370, x71202, x5667);
  nand n14371(x14371, x1448, x5537);
  nand n14372(x14372, x14371, x14370);
  nand n14373(x14373, x71205, x14363);
  nand n14374(x14374, x1461, x14366);
  nand n14375(x14375, x14374, x14373);
  nand n14376(x14376, x71205, x14369);
  nand n14377(x14377, x1461, x14372);
  nand n14378(x14378, x14377, x14376);
  nand n14379(x14379, x71210, x14375);
  nand n14380(x14380, x1468, x14378);
  nand n14381(x14381, x14380, x14379);
  nand n14382(x14382, x71202, x6451);
  nand n14383(x14383, x1448, x6321);
  nand n14384(x14384, x14383, x14382);
  nand n14385(x14385, x71202, x6191);
  nand n14386(x14386, x1448, x6061);
  nand n14387(x14387, x14386, x14385);
  nand n14388(x14388, x71202, x5931);
  nand n14389(x14389, x1448, x5801);
  nand n14390(x14390, x14389, x14388);
  nand n14391(x14391, x71202, x5671);
  nand n14392(x14392, x1448, x5541);
  nand n14393(x14393, x14392, x14391);
  nand n14394(x14394, x71205, x14384);
  nand n14395(x14395, x1461, x14387);
  nand n14396(x14396, x14395, x14394);
  nand n14397(x14397, x71205, x14390);
  nand n14398(x14398, x1461, x14393);
  nand n14399(x14399, x14398, x14397);
  nand n14400(x14400, x71210, x14396);
  nand n14401(x14401, x1468, x14399);
  nand n14402(x14402, x14401, x14400);
  nand n14403(x14403, x71202, x6455);
  nand n14404(x14404, x1448, x6325);
  nand n14405(x14405, x14404, x14403);
  nand n14406(x14406, x71202, x6195);
  nand n14407(x14407, x1448, x6065);
  nand n14408(x14408, x14407, x14406);
  nand n14409(x14409, x71202, x5935);
  nand n14410(x14410, x1448, x5805);
  nand n14411(x14411, x14410, x14409);
  nand n14412(x14412, x71202, x5675);
  nand n14413(x14413, x1448, x5545);
  nand n14414(x14414, x14413, x14412);
  nand n14415(x14415, x71205, x14405);
  nand n14416(x14416, x1461, x14408);
  nand n14417(x14417, x14416, x14415);
  nand n14418(x14418, x71205, x14411);
  nand n14419(x14419, x1461, x14414);
  nand n14420(x14420, x14419, x14418);
  nand n14421(x14421, x71210, x14417);
  nand n14422(x14422, x1468, x14420);
  nand n14423(x14423, x14422, x14421);
  nand n14424(x14424, x71202, x6459);
  nand n14425(x14425, x1448, x6329);
  nand n14426(x14426, x14425, x14424);
  nand n14427(x14427, x71202, x6199);
  nand n14428(x14428, x1448, x6069);
  nand n14429(x14429, x14428, x14427);
  nand n14430(x14430, x71202, x5939);
  nand n14431(x14431, x1448, x5809);
  nand n14432(x14432, x14431, x14430);
  nand n14433(x14433, x71202, x5679);
  nand n14434(x14434, x1448, x5549);
  nand n14435(x14435, x14434, x14433);
  nand n14436(x14436, x71205, x14426);
  nand n14437(x14437, x1461, x14429);
  nand n14438(x14438, x14437, x14436);
  nand n14439(x14439, x71205, x14432);
  nand n14440(x14440, x1461, x14435);
  nand n14441(x14441, x14440, x14439);
  nand n14442(x14442, x71210, x14438);
  nand n14443(x14443, x1468, x14441);
  nand n14444(x14444, x14443, x14442);
  nand n14445(x14445, x71202, x6463);
  nand n14446(x14446, x1448, x6333);
  nand n14447(x14447, x14446, x14445);
  nand n14448(x14448, x71202, x6203);
  nand n14449(x14449, x1448, x6073);
  nand n14450(x14450, x14449, x14448);
  nand n14451(x14451, x71202, x5943);
  nand n14452(x14452, x1448, x5813);
  nand n14453(x14453, x14452, x14451);
  nand n14454(x14454, x71202, x5683);
  nand n14455(x14455, x1448, x5553);
  nand n14456(x14456, x14455, x14454);
  nand n14457(x14457, x71205, x14447);
  nand n14458(x14458, x1461, x14450);
  nand n14459(x14459, x14458, x14457);
  nand n14460(x14460, x71205, x14453);
  nand n14461(x14461, x1461, x14456);
  nand n14462(x14462, x14461, x14460);
  nand n14463(x14463, x71210, x14459);
  nand n14464(x14464, x1468, x14462);
  nand n14465(x14465, x14464, x14463);
  nand n14466(x14466, x71202, x6467);
  nand n14467(x14467, x1448, x6337);
  nand n14468(x14468, x14467, x14466);
  nand n14469(x14469, x71202, x6207);
  nand n14470(x14470, x1448, x6077);
  nand n14471(x14471, x14470, x14469);
  nand n14472(x14472, x71202, x5947);
  nand n14473(x14473, x1448, x5817);
  nand n14474(x14474, x14473, x14472);
  nand n14475(x14475, x71202, x5687);
  nand n14476(x14476, x1448, x5557);
  nand n14477(x14477, x14476, x14475);
  nand n14478(x14478, x71205, x14468);
  nand n14479(x14479, x1461, x14471);
  nand n14480(x14480, x14479, x14478);
  nand n14481(x14481, x71205, x14474);
  nand n14482(x14482, x1461, x14477);
  nand n14483(x14483, x14482, x14481);
  nand n14484(x14484, x71210, x14480);
  nand n14485(x14485, x1468, x14483);
  nand n14486(x14486, x14485, x14484);
  nand n14487(x14487, x71202, x6471);
  nand n14488(x14488, x1448, x6341);
  nand n14489(x14489, x14488, x14487);
  nand n14490(x14490, x71202, x6211);
  nand n14491(x14491, x1448, x6081);
  nand n14492(x14492, x14491, x14490);
  nand n14493(x14493, x71202, x5951);
  nand n14494(x14494, x1448, x5821);
  nand n14495(x14495, x14494, x14493);
  nand n14496(x14496, x71202, x5691);
  nand n14497(x14497, x1448, x5561);
  nand n14498(x14498, x14497, x14496);
  nand n14499(x14499, x71205, x14489);
  nand n14500(x14500, x1461, x14492);
  nand n14501(x14501, x14500, x14499);
  nand n14502(x14502, x71205, x14495);
  nand n14503(x14503, x1461, x14498);
  nand n14504(x14504, x14503, x14502);
  nand n14505(x14505, x71210, x14501);
  nand n14506(x14506, x1468, x14504);
  nand n14507(x14507, x14506, x14505);
  nand n14508(x14508, x71202, x6475);
  nand n14509(x14509, x1448, x6345);
  nand n14510(x14510, x14509, x14508);
  nand n14511(x14511, x71202, x6215);
  nand n14512(x14512, x1448, x6085);
  nand n14513(x14513, x14512, x14511);
  nand n14514(x14514, x71202, x5955);
  nand n14515(x14515, x1448, x5825);
  nand n14516(x14516, x14515, x14514);
  nand n14517(x14517, x71202, x5695);
  nand n14518(x14518, x1448, x5565);
  nand n14519(x14519, x14518, x14517);
  nand n14520(x14520, x71205, x14510);
  nand n14521(x14521, x1461, x14513);
  nand n14522(x14522, x14521, x14520);
  nand n14523(x14523, x71205, x14516);
  nand n14524(x14524, x1461, x14519);
  nand n14525(x14525, x14524, x14523);
  nand n14526(x14526, x71210, x14522);
  nand n14527(x14527, x1468, x14525);
  nand n14528(x14528, x14527, x14526);
  nand n14529(x14529, x71202, x6479);
  nand n14530(x14530, x1448, x6349);
  nand n14531(x14531, x14530, x14529);
  nand n14532(x14532, x71202, x6219);
  nand n14533(x14533, x1448, x6089);
  nand n14534(x14534, x14533, x14532);
  nand n14535(x14535, x71202, x5959);
  nand n14536(x14536, x1448, x5829);
  nand n14537(x14537, x14536, x14535);
  nand n14538(x14538, x71202, x5699);
  nand n14539(x14539, x1448, x5569);
  nand n14540(x14540, x14539, x14538);
  nand n14541(x14541, x71205, x14531);
  nand n14542(x14542, x1461, x14534);
  nand n14543(x14543, x14542, x14541);
  nand n14544(x14544, x71205, x14537);
  nand n14545(x14545, x1461, x14540);
  nand n14546(x14546, x14545, x14544);
  nand n14547(x14547, x71210, x14543);
  nand n14548(x14548, x1468, x14546);
  nand n14549(x14549, x14548, x14547);
  nand n14550(x14550, x1703, x2247);
  nand n14551(x14551, x1707, x2247);
  nand n14552(x14552, x1703, x2250);
  nand n14553(x14553, x1707, x2250);
  nand n14554(x14554, x14553, x14552);
  nand n14556(x14556, x14555, x14551);
  nand n14558(x14558, x14557, x14550);
  nand n14559(x14559, x14558, x1);
  nand n14561(x14561, x1693, x14560);
  nand n14562(x14562, x1695, x14560);
  nand n14563(x14563, x1697, x14560);
  nand n14564(x14564, x1699, x14560);
  nand n14565(x14565, x14563, x14564);
  nand n14566(x14566, x14561, x14562);
  nand n14569(x14569, x14568, x14567);
  nand n14570(x14570, x1727, x14569);
  nand n14572(x14572, x71240, x14569);
  nand n14574(x14574, x1732, x14571);
  nand n14576(x14576, x71235, x14571);
  nand n14578(x14578, x1732, x14573);
  nand n14580(x14580, x71235, x14573);
  nand n14582(x14582, x1741, x14575);
  nand n14583(x14583, x71230, x14575);
  nand n14584(x14584, x1741, x14577);
  nand n14585(x14585, x71230, x14577);
  nand n14586(x14586, x1741, x14579);
  nand n14587(x14587, x71230, x14579);
  nand n14588(x14588, x1741, x14581);
  nand n14589(x14589, x71230, x14581);
  nand n14590(x14590, x2297, x14582);
  nand n14592(x14592, x2296, x14582);
  nand n14593(x14593, x14592, x14591);
  nand n14595(x14595, x14594, x14599);
  nand n14596(x14596, x14595, x14593);
  nand n14600(x14600, x2299, x14583);
  nand n14602(x14602, x2298, x14583);
  nand n14603(x14603, x14602, x14601);
  nand n14605(x14605, x14604, x14609);
  nand n14606(x14606, x14605, x14603);
  nand n14610(x14610, x2301, x14584);
  nand n14612(x14612, x2300, x14584);
  nand n14613(x14613, x14612, x14611);
  nand n14615(x14615, x14614, x14619);
  nand n14616(x14616, x14615, x14613);
  nand n14620(x14620, x2303, x14585);
  nand n14622(x14622, x2302, x14585);
  nand n14623(x14623, x14622, x14621);
  nand n14625(x14625, x14624, x14629);
  nand n14626(x14626, x14625, x14623);
  nand n14630(x14630, x2305, x14586);
  nand n14632(x14632, x2304, x14586);
  nand n14633(x14633, x14632, x14631);
  nand n14635(x14635, x14634, x14639);
  nand n14636(x14636, x14635, x14633);
  nand n14640(x14640, x2307, x14587);
  nand n14642(x14642, x2306, x14587);
  nand n14643(x14643, x14642, x14641);
  nand n14645(x14645, x14644, x14649);
  nand n14646(x14646, x14645, x14643);
  nand n14650(x14650, x2309, x14588);
  nand n14652(x14652, x2308, x14588);
  nand n14653(x14653, x14652, x14651);
  nand n14655(x14655, x14654, x14659);
  nand n14656(x14656, x14655, x14653);
  nand n14660(x14660, x2311, x14589);
  nand n14662(x14662, x2310, x14589);
  nand n14663(x14663, x14662, x14661);
  nand n14665(x14665, x14664, x14669);
  nand n14666(x14666, x14665, x14663);
  nand n14670(x14670, x2258, x14669);
  nand n14671(x14671, x6481, x14659);
  nand n14672(x14672, x14671, x14670);
  nand n14673(x14673, x2258, x14649);
  nand n14674(x14674, x6481, x14639);
  nand n14675(x14675, x14674, x14673);
  nand n14676(x14676, x2258, x14629);
  nand n14677(x14677, x6481, x14619);
  nand n14678(x14678, x14677, x14676);
  nand n14679(x14679, x2258, x14609);
  nand n14680(x14680, x6481, x14599);
  nand n14681(x14681, x14680, x14679);
  nand n14682(x14682, x2261, x14672);
  nand n14683(x14683, x6494, x14675);
  nand n14684(x14684, x14683, x14682);
  nand n14685(x14685, x2261, x14678);
  nand n14686(x14686, x6494, x14681);
  nand n14687(x14687, x14686, x14685);
  nand n14688(x14688, x2264, x14684);
  nand n14689(x14689, x6501, x14687);
  nand n14690(x14690, x14689, x14688);
  nand n14691(x14691, x2269, x14669);
  nand n14692(x14692, x7156, x14659);
  nand n14693(x14693, x14692, x14691);
  nand n14694(x14694, x2269, x14649);
  nand n14695(x14695, x7156, x14639);
  nand n14696(x14696, x14695, x14694);
  nand n14697(x14697, x2269, x14629);
  nand n14698(x14698, x7156, x14619);
  nand n14699(x14699, x14698, x14697);
  nand n14700(x14700, x2269, x14609);
  nand n14701(x14701, x7156, x14599);
  nand n14702(x14702, x14701, x14700);
  nand n14703(x14703, x2272, x14693);
  nand n14704(x14704, x7169, x14696);
  nand n14705(x14705, x14704, x14703);
  nand n14706(x14706, x2272, x14699);
  nand n14707(x14707, x7169, x14702);
  nand n14708(x14708, x14707, x14706);
  nand n14709(x14709, x2275, x14705);
  nand n14710(x14710, x7176, x14708);
  nand n14711(x14711, x14710, x14709);
  nand n14712(x14712, x71202, x14669);
  nand n14713(x14713, x1448, x14659);
  nand n14714(x14714, x14713, x14712);
  nand n14715(x14715, x71202, x14649);
  nand n14716(x14716, x1448, x14639);
  nand n14717(x14717, x14716, x14715);
  nand n14718(x14718, x71202, x14629);
  nand n14719(x14719, x1448, x14619);
  nand n14720(x14720, x14719, x14718);
  nand n14721(x14721, x71202, x14609);
  nand n14722(x14722, x1448, x14599);
  nand n14723(x14723, x14722, x14721);
  nand n14724(x14724, x71205, x14714);
  nand n14725(x14725, x1461, x14717);
  nand n14726(x14726, x14725, x14724);
  nand n14727(x14727, x71205, x14720);
  nand n14728(x14728, x1461, x14723);
  nand n14729(x14729, x14728, x14727);
  nand n14730(x14730, x71210, x14726);
  nand n14731(x14731, x1468, x14729);
  nand n14732(x14732, x14731, x14730);
  nand n14734(x14734, x2251, x14553);
  nand n14736(x14736, x14735, x14552);
  nand n14738(x14738, x14737, x2248);
  nand n14740(x14740, x14739, x14550);
  nand n14742(x14742, x14741, x2245);
  nand n14744(x14744, x14743, x1712);
  nand n14745(x14745, x14744, x14733);
  nand n14747(x14747, x14552, x2248);
  nand n14749(x14749, x14748, x2245);
  nand n14750(x14750, x14749, x14746);
  nand n14753(x14753, x14752, x14751);
  nand n14762(x14762, x14754, x14569);
  nand n14764(x14764, x14763, x71454);
  nand n14765(x14765, x14762, x14767);
  nand n14766(x14766, x14765, x14764);
  nand n14768(x14768, x14763, x71459);
  nand n14769(x14769, x14762, x14771);
  nand n14770(x14770, x14769, x14768);
  nand n14772(x14772, x14763, x71464);
  nand n14773(x14773, x14762, x14775);
  nand n14774(x14774, x14773, x14772);
  nand n14776(x14776, x14763, x71469);
  nand n14777(x14777, x14762, x14779);
  nand n14778(x14778, x14777, x14776);
  nand n14780(x14780, x14763, x71474);
  nand n14781(x14781, x14762, x14783);
  nand n14782(x14782, x14781, x14780);
  nand n14784(x14784, x14763, x71479);
  nand n14785(x14785, x14762, x14787);
  nand n14786(x14786, x14785, x14784);
  nand n14788(x14788, x14755, x14569);
  nand n14790(x14790, x14789, x71454);
  nand n14791(x14791, x14788, x14793);
  nand n14792(x14792, x14791, x14790);
  nand n14794(x14794, x14789, x71459);
  nand n14795(x14795, x14788, x14797);
  nand n14796(x14796, x14795, x14794);
  nand n14798(x14798, x14789, x71464);
  nand n14799(x14799, x14788, x14801);
  nand n14800(x14800, x14799, x14798);
  nand n14802(x14802, x14789, x71469);
  nand n14803(x14803, x14788, x14805);
  nand n14804(x14804, x14803, x14802);
  nand n14806(x14806, x14789, x71474);
  nand n14807(x14807, x14788, x14809);
  nand n14808(x14808, x14807, x14806);
  nand n14810(x14810, x14789, x71479);
  nand n14811(x14811, x14788, x14813);
  nand n14812(x14812, x14811, x14810);
  nand n14814(x14814, x14756, x14569);
  nand n14816(x14816, x14815, x71454);
  nand n14817(x14817, x14814, x14819);
  nand n14818(x14818, x14817, x14816);
  nand n14820(x14820, x14815, x71459);
  nand n14821(x14821, x14814, x14823);
  nand n14822(x14822, x14821, x14820);
  nand n14824(x14824, x14815, x71464);
  nand n14825(x14825, x14814, x14827);
  nand n14826(x14826, x14825, x14824);
  nand n14828(x14828, x14815, x71469);
  nand n14829(x14829, x14814, x14831);
  nand n14830(x14830, x14829, x14828);
  nand n14832(x14832, x14815, x71474);
  nand n14833(x14833, x14814, x14835);
  nand n14834(x14834, x14833, x14832);
  nand n14836(x14836, x14815, x71479);
  nand n14837(x14837, x14814, x14839);
  nand n14838(x14838, x14837, x14836);
  nand n14840(x14840, x14757, x14569);
  nand n14842(x14842, x14841, x71454);
  nand n14843(x14843, x14840, x14845);
  nand n14844(x14844, x14843, x14842);
  nand n14846(x14846, x14841, x71459);
  nand n14847(x14847, x14840, x14849);
  nand n14848(x14848, x14847, x14846);
  nand n14850(x14850, x14841, x71464);
  nand n14851(x14851, x14840, x14853);
  nand n14852(x14852, x14851, x14850);
  nand n14854(x14854, x14841, x71469);
  nand n14855(x14855, x14840, x14857);
  nand n14856(x14856, x14855, x14854);
  nand n14858(x14858, x14841, x71474);
  nand n14859(x14859, x14840, x14861);
  nand n14860(x14860, x14859, x14858);
  nand n14862(x14862, x14841, x71479);
  nand n14863(x14863, x14840, x14865);
  nand n14864(x14864, x14863, x14862);
  nand n14866(x14866, x14758, x14569);
  nand n14868(x14868, x14867, x71454);
  nand n14869(x14869, x14866, x14871);
  nand n14870(x14870, x14869, x14868);
  nand n14872(x14872, x14867, x71459);
  nand n14873(x14873, x14866, x14875);
  nand n14874(x14874, x14873, x14872);
  nand n14876(x14876, x14867, x71464);
  nand n14877(x14877, x14866, x14879);
  nand n14878(x14878, x14877, x14876);
  nand n14880(x14880, x14867, x71469);
  nand n14881(x14881, x14866, x14883);
  nand n14882(x14882, x14881, x14880);
  nand n14884(x14884, x14867, x71474);
  nand n14885(x14885, x14866, x14887);
  nand n14886(x14886, x14885, x14884);
  nand n14888(x14888, x14867, x71479);
  nand n14889(x14889, x14866, x14891);
  nand n14890(x14890, x14889, x14888);
  nand n14892(x14892, x14759, x14569);
  nand n14894(x14894, x14893, x71454);
  nand n14895(x14895, x14892, x14897);
  nand n14896(x14896, x14895, x14894);
  nand n14898(x14898, x14893, x71459);
  nand n14899(x14899, x14892, x14901);
  nand n14900(x14900, x14899, x14898);
  nand n14902(x14902, x14893, x71464);
  nand n14903(x14903, x14892, x14905);
  nand n14904(x14904, x14903, x14902);
  nand n14906(x14906, x14893, x71469);
  nand n14907(x14907, x14892, x14909);
  nand n14908(x14908, x14907, x14906);
  nand n14910(x14910, x14893, x71474);
  nand n14911(x14911, x14892, x14913);
  nand n14912(x14912, x14911, x14910);
  nand n14914(x14914, x14893, x71479);
  nand n14915(x14915, x14892, x14917);
  nand n14916(x14916, x14915, x14914);
  nand n14918(x14918, x14760, x14569);
  nand n14920(x14920, x14919, x71454);
  nand n14921(x14921, x14918, x14923);
  nand n14922(x14922, x14921, x14920);
  nand n14924(x14924, x14919, x71459);
  nand n14925(x14925, x14918, x14927);
  nand n14926(x14926, x14925, x14924);
  nand n14928(x14928, x14919, x71464);
  nand n14929(x14929, x14918, x14931);
  nand n14930(x14930, x14929, x14928);
  nand n14932(x14932, x14919, x71469);
  nand n14933(x14933, x14918, x14935);
  nand n14934(x14934, x14933, x14932);
  nand n14936(x14936, x14919, x71474);
  nand n14937(x14937, x14918, x14939);
  nand n14938(x14938, x14937, x14936);
  nand n14940(x14940, x14919, x71479);
  nand n14941(x14941, x14918, x14943);
  nand n14942(x14942, x14941, x14940);
  nand n14944(x14944, x14761, x14569);
  nand n14946(x14946, x14945, x71454);
  nand n14947(x14947, x14944, x14949);
  nand n14948(x14948, x14947, x14946);
  nand n14950(x14950, x14945, x71459);
  nand n14951(x14951, x14944, x14953);
  nand n14952(x14952, x14951, x14950);
  nand n14954(x14954, x14945, x71464);
  nand n14955(x14955, x14944, x14957);
  nand n14956(x14956, x14955, x14954);
  nand n14958(x14958, x14945, x71469);
  nand n14959(x14959, x14944, x14961);
  nand n14960(x14960, x14959, x14958);
  nand n14962(x14962, x14945, x71474);
  nand n14963(x14963, x14944, x14965);
  nand n14964(x14964, x14963, x14962);
  nand n14966(x14966, x14945, x71479);
  nand n14967(x14967, x14944, x14969);
  nand n14968(x14968, x14967, x14966);
  nand n14970(x14970, x70689, x14949);
  nand n14971(x14971, x2295, x14923);
  nand n14972(x14972, x14971, x14970);
  nand n14973(x14973, x70689, x14897);
  nand n14974(x14974, x2295, x14871);
  nand n14975(x14975, x14974, x14973);
  nand n14976(x14976, x70689, x14845);
  nand n14977(x14977, x2295, x14819);
  nand n14978(x14978, x14977, x14976);
  nand n14979(x14979, x70689, x14793);
  nand n14980(x14980, x2295, x14767);
  nand n14981(x14981, x14980, x14979);
  nand n14982(x14982, x70705, x14972);
  nand n14983(x14983, x2286, x14975);
  nand n14984(x14984, x14983, x14982);
  nand n14985(x14985, x70705, x14978);
  nand n14986(x14986, x2286, x14981);
  nand n14987(x14987, x14986, x14985);
  nand n14988(x14988, x70721, x14984);
  nand n14989(x14989, x2281, x14987);
  nand n14990(x14990, x14989, x14988);
  nand n14991(x14991, x70689, x14953);
  nand n14992(x14992, x2295, x14927);
  nand n14993(x14993, x14992, x14991);
  nand n14994(x14994, x70689, x14901);
  nand n14995(x14995, x2295, x14875);
  nand n14996(x14996, x14995, x14994);
  nand n14997(x14997, x70689, x14849);
  nand n14998(x14998, x2295, x14823);
  nand n14999(x14999, x14998, x14997);
  nand n15000(x15000, x70689, x14797);
  nand n15001(x15001, x2295, x14771);
  nand n15002(x15002, x15001, x15000);
  nand n15003(x15003, x70705, x14993);
  nand n15004(x15004, x2286, x14996);
  nand n15005(x15005, x15004, x15003);
  nand n15006(x15006, x70705, x14999);
  nand n15007(x15007, x2286, x15002);
  nand n15008(x15008, x15007, x15006);
  nand n15009(x15009, x70721, x15005);
  nand n15010(x15010, x2281, x15008);
  nand n15011(x15011, x15010, x15009);
  nand n15012(x15012, x70689, x14957);
  nand n15013(x15013, x2295, x14931);
  nand n15014(x15014, x15013, x15012);
  nand n15015(x15015, x70689, x14905);
  nand n15016(x15016, x2295, x14879);
  nand n15017(x15017, x15016, x15015);
  nand n15018(x15018, x70689, x14853);
  nand n15019(x15019, x2295, x14827);
  nand n15020(x15020, x15019, x15018);
  nand n15021(x15021, x70689, x14801);
  nand n15022(x15022, x2295, x14775);
  nand n15023(x15023, x15022, x15021);
  nand n15024(x15024, x70705, x15014);
  nand n15025(x15025, x2286, x15017);
  nand n15026(x15026, x15025, x15024);
  nand n15027(x15027, x70705, x15020);
  nand n15028(x15028, x2286, x15023);
  nand n15029(x15029, x15028, x15027);
  nand n15030(x15030, x70721, x15026);
  nand n15031(x15031, x2281, x15029);
  nand n15032(x15032, x15031, x15030);
  nand n15033(x15033, x70689, x14961);
  nand n15034(x15034, x2295, x14935);
  nand n15035(x15035, x15034, x15033);
  nand n15036(x15036, x70689, x14909);
  nand n15037(x15037, x2295, x14883);
  nand n15038(x15038, x15037, x15036);
  nand n15039(x15039, x70689, x14857);
  nand n15040(x15040, x2295, x14831);
  nand n15041(x15041, x15040, x15039);
  nand n15042(x15042, x70689, x14805);
  nand n15043(x15043, x2295, x14779);
  nand n15044(x15044, x15043, x15042);
  nand n15045(x15045, x70705, x15035);
  nand n15046(x15046, x2286, x15038);
  nand n15047(x15047, x15046, x15045);
  nand n15048(x15048, x70705, x15041);
  nand n15049(x15049, x2286, x15044);
  nand n15050(x15050, x15049, x15048);
  nand n15051(x15051, x70721, x15047);
  nand n15052(x15052, x2281, x15050);
  nand n15053(x15053, x15052, x15051);
  nand n15054(x15054, x70689, x14965);
  nand n15055(x15055, x2295, x14939);
  nand n15056(x15056, x15055, x15054);
  nand n15057(x15057, x70689, x14913);
  nand n15058(x15058, x2295, x14887);
  nand n15059(x15059, x15058, x15057);
  nand n15060(x15060, x70689, x14861);
  nand n15061(x15061, x2295, x14835);
  nand n15062(x15062, x15061, x15060);
  nand n15063(x15063, x70689, x14809);
  nand n15064(x15064, x2295, x14783);
  nand n15065(x15065, x15064, x15063);
  nand n15066(x15066, x70705, x15056);
  nand n15067(x15067, x2286, x15059);
  nand n15068(x15068, x15067, x15066);
  nand n15069(x15069, x70705, x15062);
  nand n15070(x15070, x2286, x15065);
  nand n15071(x15071, x15070, x15069);
  nand n15072(x15072, x70721, x15068);
  nand n15073(x15073, x2281, x15071);
  nand n15074(x15074, x15073, x15072);
  nand n15075(x15075, x70689, x14969);
  nand n15076(x15076, x2295, x14943);
  nand n15077(x15077, x15076, x15075);
  nand n15078(x15078, x70689, x14917);
  nand n15079(x15079, x2295, x14891);
  nand n15080(x15080, x15079, x15078);
  nand n15081(x15081, x70689, x14865);
  nand n15082(x15082, x2295, x14839);
  nand n15083(x15083, x15082, x15081);
  nand n15084(x15084, x70689, x14813);
  nand n15085(x15085, x2295, x14787);
  nand n15086(x15086, x15085, x15084);
  nand n15087(x15087, x70705, x15077);
  nand n15088(x15088, x2286, x15080);
  nand n15089(x15089, x15088, x15087);
  nand n15090(x15090, x70705, x15083);
  nand n15091(x15091, x2286, x15086);
  nand n15092(x15092, x15091, x15090);
  nand n15093(x15093, x70721, x15089);
  nand n15094(x15094, x2281, x15092);
  nand n15095(x15095, x15094, x15093);
  nand n15097(x15097, x15096, x71147);
  nand n15098(x15098, x14551, x71147);
  nand n15099(x15099, x15098, x15097);
  nand n15100(x15100, x15096, x71152);
  nand n15101(x15101, x14551, x71152);
  nand n15102(x15102, x15101, x15100);
  nand n15103(x15103, x15096, x71157);
  nand n15104(x15104, x14551, x71157);
  nand n15105(x15105, x15104, x15103);
  nand n15106(x15106, x15096, x71162);
  nand n15107(x15107, x14551, x71162);
  nand n15108(x15108, x15107, x15106);
  nand n15109(x15109, x15096, x71167);
  nand n15110(x15110, x14551, x71167);
  nand n15111(x15111, x15110, x15109);
  nand n15112(x15112, x15096, x71172);
  nand n15113(x15113, x14551, x71172);
  nand n15114(x15114, x15113, x15112);
  nand n15115(x15115, x15096, x71177);
  nand n15116(x15116, x14551, x71177);
  nand n15117(x15117, x15116, x15115);
  nand n15118(x15118, x15096, x71182);
  nand n15119(x15119, x14551, x71182);
  nand n15120(x15120, x15119, x15118);
  nand n15121(x15121, x15096, x71185);
  nand n15122(x15122, x14551, x71185);
  nand n15123(x15123, x15122, x15121);
  nand n15124(x15124, x15096, x71188);
  nand n15125(x15125, x14551, x71188);
  nand n15126(x15126, x15125, x15124);
  nand n15127(x15127, x15096, x71191);
  nand n15128(x15128, x14551, x71191);
  nand n15129(x15129, x15128, x15127);
  nand n15130(x15130, x15096, x71194);
  nand n15131(x15131, x14551, x71194);
  nand n15132(x15132, x15131, x15130);
  nand n15133(x15133, x15096, x71197);
  nand n15134(x15134, x14551, x71197);
  nand n15135(x15135, x15134, x15133);
  nand n15136(x15136, x15096, x71202);
  nand n15137(x15137, x14551, x71202);
  nand n15138(x15138, x15137, x15136);
  nand n15139(x15139, x15096, x71205);
  nand n15140(x15140, x14551, x71205);
  nand n15141(x15141, x15140, x15139);
  nand n15142(x15142, x15096, x71210);
  nand n15143(x15143, x14551, x71210);
  nand n15144(x15144, x15143, x15142);
  nand n15145(x15145, x15096, x71215);
  nand n15146(x15146, x15143, x15145);
  nand n15147(x15147, x15096, x71220);
  nand n15148(x15148, x15143, x15147);
  nand n15149(x15149, x15096, x71225);
  nand n15150(x15150, x15143, x15149);
  nand n15151(x15151, x1711, x2247);
  nand n15153(x15153, x15152, x71147);
  nand n15154(x15154, x15151, x15099);
  nand n15155(x15155, x15154, x15153);
  nand n15156(x15156, x15152, x71152);
  nand n15157(x15157, x15151, x15102);
  nand n15158(x15158, x15157, x15156);
  nand n15159(x15159, x15152, x71157);
  nand n15160(x15160, x15151, x15105);
  nand n15161(x15161, x15160, x15159);
  nand n15162(x15162, x15152, x71162);
  nand n15163(x15163, x15151, x15108);
  nand n15164(x15164, x15163, x15162);
  nand n15165(x15165, x15152, x71167);
  nand n15166(x15166, x15151, x15111);
  nand n15167(x15167, x15166, x15165);
  nand n15168(x15168, x15152, x71172);
  nand n15169(x15169, x15151, x15114);
  nand n15170(x15170, x15169, x15168);
  nand n15171(x15171, x15152, x71177);
  nand n15172(x15172, x15151, x15117);
  nand n15173(x15173, x15172, x15171);
  nand n15174(x15174, x15152, x71182);
  nand n15175(x15175, x15151, x15120);
  nand n15176(x15176, x15175, x15174);
  nand n15177(x15177, x15152, x71185);
  nand n15178(x15178, x15151, x15123);
  nand n15179(x15179, x15178, x15177);
  nand n15180(x15180, x15152, x71188);
  nand n15181(x15181, x15151, x15126);
  nand n15182(x15182, x15181, x15180);
  nand n15183(x15183, x15152, x71191);
  nand n15184(x15184, x15151, x15129);
  nand n15185(x15185, x15184, x15183);
  nand n15186(x15186, x15152, x71194);
  nand n15187(x15187, x15151, x15132);
  nand n15188(x15188, x15187, x15186);
  nand n15189(x15189, x15152, x71197);
  nand n15190(x15190, x15151, x15135);
  nand n15191(x15191, x15190, x15189);
  nand n15192(x15192, x15152, x71202);
  nand n15193(x15193, x15151, x15138);
  nand n15194(x15194, x15193, x15192);
  nand n15195(x15195, x15152, x71205);
  nand n15196(x15196, x15151, x15141);
  nand n15197(x15197, x15196, x15195);
  nand n15198(x15198, x15152, x71210);
  nand n15199(x15199, x15151, x15144);
  nand n15200(x15200, x15199, x15198);
  nand n15201(x15201, x15152, x71215);
  nand n15202(x15202, x15151, x15146);
  nand n15203(x15203, x15202, x15201);
  nand n15204(x15204, x15152, x71220);
  nand n15205(x15205, x15151, x15148);
  nand n15206(x15206, x15205, x15204);
  nand n15207(x15207, x15152, x71225);
  nand n15208(x15208, x15151, x15150);
  nand n15209(x15209, x15208, x15207);
  nand n15210(x15210, x15152, x71230);
  nand n15211(x15211, x15208, x15210);
  nand n15212(x15212, x15152, x71235);
  nand n15213(x15213, x15208, x15212);
  nand n15214(x15214, x15152, x71240);
  nand n15215(x15215, x15208, x15214);
  nand n15216(x15216, x15151, x14551);
  nand n15218(x15218, x15217, x14550);
  nand n15220(x15220, x15219, x2245);
  nand n15221(x15221, x1107, x1037);
  nand n15223(x15223, x15222, x1099);
  nand n15225(x15225, x15224, x1010);
  nand n15226(x15226, x1, x1693);
  nand n15228(x15228, x15227, x15225);
  nand n15230(x15230, x71289, x15155);
  nand n15233(x15233, x15232, x15231);
  nand n15234(x15234, x15233, x15230);
  nand n15235(x15235, x71294, x15158);
  nand n15238(x15238, x15237, x15236);
  nand n15239(x15239, x15238, x15235);
  nand n15241(x15241, x71299, x15161);
  nand n15244(x15244, x15243, x15242);
  nand n15245(x15245, x15244, x15241);
  nand n15247(x15247, x71304, x15164);
  nand n15250(x15250, x15249, x15248);
  nand n15251(x15251, x15250, x15247);
  nand n15253(x15253, x71309, x15167);
  nand n15256(x15256, x15255, x15254);
  nand n15257(x15257, x15256, x15253);
  nand n15259(x15259, x71314, x15170);
  nand n15262(x15262, x15261, x15260);
  nand n15263(x15263, x15262, x15259);
  nand n15265(x15265, x71319, x15173);
  nand n15268(x15268, x15267, x15266);
  nand n15269(x15269, x15268, x15265);
  nand n15271(x15271, x71324, x15176);
  nand n15274(x15274, x15273, x15272);
  nand n15275(x15275, x15274, x15271);
  nand n15277(x15277, x71329, x15179);
  nand n15280(x15280, x15279, x15278);
  nand n15281(x15281, x15280, x15277);
  nand n15283(x15283, x71334, x15182);
  nand n15286(x15286, x15285, x15284);
  nand n15287(x15287, x15286, x15283);
  nand n15289(x15289, x71339, x15185);
  nand n15292(x15292, x15291, x15290);
  nand n15293(x15293, x15292, x15289);
  nand n15295(x15295, x71344, x15188);
  nand n15298(x15298, x15297, x15296);
  nand n15299(x15299, x15298, x15295);
  nand n15301(x15301, x71349, x15191);
  nand n15304(x15304, x15303, x15302);
  nand n15305(x15305, x15304, x15301);
  nand n15307(x15307, x71354, x15194);
  nand n15310(x15310, x15309, x15308);
  nand n15311(x15311, x15310, x15307);
  nand n15313(x15313, x71359, x15197);
  nand n15316(x15316, x15315, x15314);
  nand n15317(x15317, x15316, x15313);
  nand n15319(x15319, x71364, x15200);
  nand n15322(x15322, x15321, x15320);
  nand n15323(x15323, x15322, x15319);
  nand n15325(x15325, x71369, x15203);
  nand n15328(x15328, x15327, x15326);
  nand n15329(x15329, x15328, x15325);
  nand n15331(x15331, x71374, x15206);
  nand n15334(x15334, x15333, x15332);
  nand n15335(x15335, x15334, x15331);
  nand n15337(x15337, x71379, x15209);
  nand n15340(x15340, x15339, x15338);
  nand n15341(x15341, x15340, x15337);
  nand n15343(x15343, x71384, x15211);
  nand n15346(x15346, x15345, x15344);
  nand n15347(x15347, x15346, x15343);
  nand n15349(x15349, x71389, x15213);
  nand n15352(x15352, x15351, x15350);
  nand n15353(x15353, x15352, x15349);
  nand n15355(x15355, x71394, x15215);
  nand n15358(x15358, x15357, x15356);
  nand n15359(x15359, x15358, x15355);
  nand n15361(x15361, x71399, x15215);
  nand n15363(x15363, x15362, x15356);
  nand n15364(x15364, x15363, x15361);
  nand n15366(x15366, x71404, x15215);
  nand n15368(x15368, x15367, x15356);
  nand n15369(x15369, x15368, x15366);
  nand n15371(x15371, x71409, x15215);
  nand n15373(x15373, x15372, x15356);
  nand n15374(x15374, x15373, x15371);
  nand n15376(x15376, x71414, x15215);
  nand n15378(x15378, x15377, x15356);
  nand n15379(x15379, x15378, x15376);
  nand n15381(x15381, x71419, x15215);
  nand n15383(x15383, x15382, x15356);
  nand n15384(x15384, x15383, x15381);
  nand n15386(x15386, x71424, x15215);
  nand n15388(x15388, x15387, x15356);
  nand n15389(x15389, x15388, x15386);
  nand n15391(x15391, x71429, x15215);
  nand n15393(x15393, x15392, x15356);
  nand n15394(x15394, x15393, x15391);
  nand n15396(x15396, x71434, x15215);
  nand n15398(x15398, x15397, x15356);
  nand n15399(x15399, x15398, x15396);
  nand n15401(x15401, x71439, x15215);
  nand n15403(x15403, x15402, x15356);
  nand n15404(x15404, x15403, x15401);
  nand n15406(x15406, x71444, x15215);
  nand n15408(x15408, x15407, x15356);
  nand n15409(x15409, x15408, x15406);
  nand n15441(x15441, x15240, x15411);
  nand n15442(x15442, x15441, x15235);
  nand n15443(x15443, x15246, x15412);
  nand n15444(x15444, x15443, x15241);
  nand n15445(x15445, x15246, x15240);
  nand n15447(x15447, x15252, x15413);
  nand n15448(x15448, x15447, x15247);
  nand n15449(x15449, x15252, x15246);
  nand n15451(x15451, x15258, x15414);
  nand n15452(x15452, x15451, x15253);
  nand n15453(x15453, x15258, x15252);
  nand n15455(x15455, x15264, x15415);
  nand n15456(x15456, x15455, x15259);
  nand n15457(x15457, x15264, x15258);
  nand n15459(x15459, x15270, x15416);
  nand n15460(x15460, x15459, x15265);
  nand n15461(x15461, x15270, x15264);
  nand n15463(x15463, x15276, x15417);
  nand n15464(x15464, x15463, x15271);
  nand n15465(x15465, x15276, x15270);
  nand n15467(x15467, x15282, x15418);
  nand n15468(x15468, x15467, x15277);
  nand n15469(x15469, x15282, x15276);
  nand n15471(x15471, x15288, x15419);
  nand n15472(x15472, x15471, x15283);
  nand n15473(x15473, x15288, x15282);
  nand n15475(x15475, x15294, x15420);
  nand n15476(x15476, x15475, x15289);
  nand n15477(x15477, x15294, x15288);
  nand n15479(x15479, x15300, x15421);
  nand n15480(x15480, x15479, x15295);
  nand n15481(x15481, x15300, x15294);
  nand n15483(x15483, x15306, x15422);
  nand n15484(x15484, x15483, x15301);
  nand n15485(x15485, x15306, x15300);
  nand n15487(x15487, x15312, x15423);
  nand n15488(x15488, x15487, x15307);
  nand n15489(x15489, x15312, x15306);
  nand n15491(x15491, x15318, x15424);
  nand n15492(x15492, x15491, x15313);
  nand n15493(x15493, x15318, x15312);
  nand n15495(x15495, x15324, x15425);
  nand n15496(x15496, x15495, x15319);
  nand n15497(x15497, x15324, x15318);
  nand n15499(x15499, x15330, x15426);
  nand n15500(x15500, x15499, x15325);
  nand n15501(x15501, x15330, x15324);
  nand n15503(x15503, x15336, x15427);
  nand n15504(x15504, x15503, x15331);
  nand n15505(x15505, x15336, x15330);
  nand n15507(x15507, x15342, x15428);
  nand n15508(x15508, x15507, x15337);
  nand n15509(x15509, x15342, x15336);
  nand n15511(x15511, x15348, x15429);
  nand n15512(x15512, x15511, x15343);
  nand n15513(x15513, x15348, x15342);
  nand n15515(x15515, x15354, x15430);
  nand n15516(x15516, x15515, x15349);
  nand n15517(x15517, x15354, x15348);
  nand n15519(x15519, x15360, x15431);
  nand n15520(x15520, x15519, x15355);
  nand n15521(x15521, x15360, x15354);
  nand n15523(x15523, x15365, x15432);
  nand n15524(x15524, x15523, x15361);
  nand n15525(x15525, x15365, x15360);
  nand n15527(x15527, x15370, x15433);
  nand n15528(x15528, x15527, x15366);
  nand n15529(x15529, x15370, x15365);
  nand n15531(x15531, x15375, x15434);
  nand n15532(x15532, x15531, x15371);
  nand n15533(x15533, x15375, x15370);
  nand n15535(x15535, x15380, x15435);
  nand n15536(x15536, x15535, x15376);
  nand n15537(x15537, x15380, x15375);
  nand n15539(x15539, x15385, x15436);
  nand n15540(x15540, x15539, x15381);
  nand n15541(x15541, x15385, x15380);
  nand n15543(x15543, x15390, x15437);
  nand n15544(x15544, x15543, x15386);
  nand n15545(x15545, x15390, x15385);
  nand n15547(x15547, x15395, x15438);
  nand n15548(x15548, x15547, x15391);
  nand n15549(x15549, x15395, x15390);
  nand n15551(x15551, x15400, x15439);
  nand n15552(x15552, x15551, x15396);
  nand n15553(x15553, x15400, x15395);
  nand n15555(x15555, x15405, x15440);
  nand n15556(x15556, x15555, x15401);
  nand n15557(x15557, x15405, x15400);
  nand n15560(x15560, x15446, x15411);
  nand n15562(x15562, x15560, x15561);
  nand n15563(x15563, x15450, x15442);
  nand n15565(x15565, x15563, x15564);
  nand n15566(x15566, x15454, x15444);
  nand n15568(x15568, x15566, x15567);
  nand n15569(x15569, x15454, x15446);
  nand n15571(x15571, x15458, x15448);
  nand n15573(x15573, x15571, x15572);
  nand n15574(x15574, x15458, x15450);
  nand n15576(x15576, x15462, x15452);
  nand n15578(x15578, x15576, x15577);
  nand n15579(x15579, x15462, x15454);
  nand n15581(x15581, x15466, x15456);
  nand n15583(x15583, x15581, x15582);
  nand n15584(x15584, x15466, x15458);
  nand n15586(x15586, x15470, x15460);
  nand n15588(x15588, x15586, x15587);
  nand n15589(x15589, x15470, x15462);
  nand n15591(x15591, x15474, x15464);
  nand n15593(x15593, x15591, x15592);
  nand n15594(x15594, x15474, x15466);
  nand n15596(x15596, x15478, x15468);
  nand n15598(x15598, x15596, x15597);
  nand n15599(x15599, x15478, x15470);
  nand n15601(x15601, x15482, x15472);
  nand n15603(x15603, x15601, x15602);
  nand n15604(x15604, x15482, x15474);
  nand n15606(x15606, x15486, x15476);
  nand n15608(x15608, x15606, x15607);
  nand n15609(x15609, x15486, x15478);
  nand n15611(x15611, x15490, x15480);
  nand n15613(x15613, x15611, x15612);
  nand n15614(x15614, x15490, x15482);
  nand n15616(x15616, x15494, x15484);
  nand n15618(x15618, x15616, x15617);
  nand n15619(x15619, x15494, x15486);
  nand n15621(x15621, x15498, x15488);
  nand n15623(x15623, x15621, x15622);
  nand n15624(x15624, x15498, x15490);
  nand n15626(x15626, x15502, x15492);
  nand n15628(x15628, x15626, x15627);
  nand n15629(x15629, x15502, x15494);
  nand n15631(x15631, x15506, x15496);
  nand n15633(x15633, x15631, x15632);
  nand n15634(x15634, x15506, x15498);
  nand n15636(x15636, x15510, x15500);
  nand n15638(x15638, x15636, x15637);
  nand n15639(x15639, x15510, x15502);
  nand n15641(x15641, x15514, x15504);
  nand n15643(x15643, x15641, x15642);
  nand n15644(x15644, x15514, x15506);
  nand n15646(x15646, x15518, x15508);
  nand n15648(x15648, x15646, x15647);
  nand n15649(x15649, x15518, x15510);
  nand n15651(x15651, x15522, x15512);
  nand n15653(x15653, x15651, x15652);
  nand n15654(x15654, x15522, x15514);
  nand n15656(x15656, x15526, x15516);
  nand n15658(x15658, x15656, x15657);
  nand n15659(x15659, x15526, x15518);
  nand n15661(x15661, x15530, x15520);
  nand n15663(x15663, x15661, x15662);
  nand n15664(x15664, x15530, x15522);
  nand n15666(x15666, x15534, x15524);
  nand n15668(x15668, x15666, x15667);
  nand n15669(x15669, x15534, x15526);
  nand n15671(x15671, x15538, x15528);
  nand n15673(x15673, x15671, x15672);
  nand n15674(x15674, x15538, x15530);
  nand n15676(x15676, x15542, x15532);
  nand n15678(x15678, x15676, x15677);
  nand n15679(x15679, x15542, x15534);
  nand n15681(x15681, x15546, x15536);
  nand n15683(x15683, x15681, x15682);
  nand n15684(x15684, x15546, x15538);
  nand n15686(x15686, x15550, x15540);
  nand n15688(x15688, x15686, x15687);
  nand n15689(x15689, x15550, x15542);
  nand n15691(x15691, x15554, x15544);
  nand n15693(x15693, x15691, x15692);
  nand n15694(x15694, x15554, x15546);
  nand n15696(x15696, x15558, x15548);
  nand n15698(x15698, x15696, x15697);
  nand n15699(x15699, x15558, x15550);
  nand n15702(x15702, x15570, x15411);
  nand n15704(x15704, x15702, x15703);
  nand n15705(x15705, x15575, x15442);
  nand n15707(x15707, x15705, x15706);
  nand n15708(x15708, x15580, x15562);
  nand n15710(x15710, x15708, x15709);
  nand n15711(x15711, x15585, x15565);
  nand n15713(x15713, x15711, x15712);
  nand n15714(x15714, x15590, x15568);
  nand n15716(x15716, x15714, x15715);
  nand n15717(x15717, x15590, x15570);
  nand n15719(x15719, x15595, x15573);
  nand n15721(x15721, x15719, x15720);
  nand n15722(x15722, x15595, x15575);
  nand n15724(x15724, x15600, x15578);
  nand n15726(x15726, x15724, x15725);
  nand n15727(x15727, x15600, x15580);
  nand n15729(x15729, x15605, x15583);
  nand n15731(x15731, x15729, x15730);
  nand n15732(x15732, x15605, x15585);
  nand n15734(x15734, x15610, x15588);
  nand n15736(x15736, x15734, x15735);
  nand n15737(x15737, x15610, x15590);
  nand n15739(x15739, x15615, x15593);
  nand n15741(x15741, x15739, x15740);
  nand n15742(x15742, x15615, x15595);
  nand n15744(x15744, x15620, x15598);
  nand n15746(x15746, x15744, x15745);
  nand n15747(x15747, x15620, x15600);
  nand n15749(x15749, x15625, x15603);
  nand n15751(x15751, x15749, x15750);
  nand n15752(x15752, x15625, x15605);
  nand n15754(x15754, x15630, x15608);
  nand n15756(x15756, x15754, x15755);
  nand n15757(x15757, x15630, x15610);
  nand n15759(x15759, x15635, x15613);
  nand n15761(x15761, x15759, x15760);
  nand n15762(x15762, x15635, x15615);
  nand n15764(x15764, x15640, x15618);
  nand n15766(x15766, x15764, x15765);
  nand n15767(x15767, x15640, x15620);
  nand n15769(x15769, x15645, x15623);
  nand n15771(x15771, x15769, x15770);
  nand n15772(x15772, x15645, x15625);
  nand n15774(x15774, x15650, x15628);
  nand n15776(x15776, x15774, x15775);
  nand n15777(x15777, x15650, x15630);
  nand n15779(x15779, x15655, x15633);
  nand n15781(x15781, x15779, x15780);
  nand n15782(x15782, x15655, x15635);
  nand n15784(x15784, x15660, x15638);
  nand n15786(x15786, x15784, x15785);
  nand n15787(x15787, x15660, x15640);
  nand n15789(x15789, x15665, x15643);
  nand n15791(x15791, x15789, x15790);
  nand n15792(x15792, x15665, x15645);
  nand n15794(x15794, x15670, x15648);
  nand n15796(x15796, x15794, x15795);
  nand n15797(x15797, x15670, x15650);
  nand n15799(x15799, x15675, x15653);
  nand n15801(x15801, x15799, x15800);
  nand n15802(x15802, x15675, x15655);
  nand n15804(x15804, x15680, x15658);
  nand n15806(x15806, x15804, x15805);
  nand n15807(x15807, x15680, x15660);
  nand n15809(x15809, x15685, x15663);
  nand n15811(x15811, x15809, x15810);
  nand n15812(x15812, x15685, x15665);
  nand n15814(x15814, x15690, x15668);
  nand n15816(x15816, x15814, x15815);
  nand n15817(x15817, x15690, x15670);
  nand n15819(x15819, x15695, x15673);
  nand n15821(x15821, x15819, x15820);
  nand n15822(x15822, x15695, x15675);
  nand n15824(x15824, x15700, x15678);
  nand n15826(x15826, x15824, x15825);
  nand n15827(x15827, x15700, x15680);
  nand n15830(x15830, x15718, x15411);
  nand n15832(x15832, x15830, x15831);
  nand n15833(x15833, x15723, x15442);
  nand n15835(x15835, x15833, x15834);
  nand n15836(x15836, x15728, x15562);
  nand n15838(x15838, x15836, x15837);
  nand n15839(x15839, x15733, x15565);
  nand n15841(x15841, x15839, x15840);
  nand n15842(x15842, x15738, x15704);
  nand n15844(x15844, x15842, x15843);
  nand n15845(x15845, x15743, x15707);
  nand n15847(x15847, x15845, x15846);
  nand n15848(x15848, x15748, x15710);
  nand n15850(x15850, x15848, x15849);
  nand n15851(x15851, x15753, x15713);
  nand n15853(x15853, x15851, x15852);
  nand n15854(x15854, x15758, x15716);
  nand n15856(x15856, x15854, x15855);
  nand n15857(x15857, x15758, x15718);
  nand n15859(x15859, x15763, x15721);
  nand n15861(x15861, x15859, x15860);
  nand n15862(x15862, x15763, x15723);
  nand n15864(x15864, x15768, x15726);
  nand n15866(x15866, x15864, x15865);
  nand n15867(x15867, x15768, x15728);
  nand n15869(x15869, x15773, x15731);
  nand n15871(x15871, x15869, x15870);
  nand n15872(x15872, x15773, x15733);
  nand n15874(x15874, x15778, x15736);
  nand n15876(x15876, x15874, x15875);
  nand n15877(x15877, x15778, x15738);
  nand n15879(x15879, x15783, x15741);
  nand n15881(x15881, x15879, x15880);
  nand n15882(x15882, x15783, x15743);
  nand n15884(x15884, x15788, x15746);
  nand n15886(x15886, x15884, x15885);
  nand n15887(x15887, x15788, x15748);
  nand n15889(x15889, x15793, x15751);
  nand n15891(x15891, x15889, x15890);
  nand n15892(x15892, x15793, x15753);
  nand n15894(x15894, x15798, x15756);
  nand n15896(x15896, x15894, x15895);
  nand n15897(x15897, x15798, x15758);
  nand n15899(x15899, x15803, x15761);
  nand n15901(x15901, x15899, x15900);
  nand n15902(x15902, x15803, x15763);
  nand n15904(x15904, x15808, x15766);
  nand n15906(x15906, x15904, x15905);
  nand n15907(x15907, x15808, x15768);
  nand n15909(x15909, x15813, x15771);
  nand n15911(x15911, x15909, x15910);
  nand n15912(x15912, x15813, x15773);
  nand n15914(x15914, x15818, x15776);
  nand n15916(x15916, x15914, x15915);
  nand n15917(x15917, x15818, x15778);
  nand n15919(x15919, x15823, x15781);
  nand n15921(x15921, x15919, x15920);
  nand n15922(x15922, x15823, x15783);
  nand n15924(x15924, x15828, x15786);
  nand n15926(x15926, x15924, x15925);
  nand n15927(x15927, x15828, x15788);
  nand n15930(x15930, x15858, x15411);
  nand n15932(x15932, x15930, x15931);
  nand n15933(x15933, x15863, x15442);
  nand n15935(x15935, x15933, x15934);
  nand n15936(x15936, x15868, x15562);
  nand n15938(x15938, x15936, x15937);
  nand n15939(x15939, x15873, x15565);
  nand n15941(x15941, x15939, x15940);
  nand n15942(x15942, x15878, x15704);
  nand n15944(x15944, x15942, x15943);
  nand n15945(x15945, x15883, x15707);
  nand n15947(x15947, x15945, x15946);
  nand n15948(x15948, x15888, x15710);
  nand n15950(x15950, x15948, x15949);
  nand n15951(x15951, x15893, x15713);
  nand n15953(x15953, x15951, x15952);
  nand n15954(x15954, x15898, x15832);
  nand n15956(x15956, x15954, x15955);
  nand n15957(x15957, x15903, x15835);
  nand n15959(x15959, x15957, x15958);
  nand n15960(x15960, x15908, x15838);
  nand n15962(x15962, x15960, x15961);
  nand n15963(x15963, x15913, x15841);
  nand n15965(x15965, x15963, x15964);
  nand n15966(x15966, x15918, x15844);
  nand n15968(x15968, x15966, x15967);
  nand n15969(x15969, x15923, x15847);
  nand n15971(x15971, x15969, x15970);
  nand n15972(x15972, x15928, x15850);
  nand n15974(x15974, x15972, x15973);
  nand n15975(x15975, x15239, x15230);
  nand n15976(x15976, x15975, x15441);
  nand n15977(x15977, x15246, x15442);
  nand n15978(x15978, x15245, x15559);
  nand n15979(x15979, x15978, x15977);
  nand n15981(x15981, x15252, x15562);
  nand n15983(x15983, x15251, x15982);
  nand n15984(x15984, x15983, x15981);
  nand n15985(x15985, x15258, x15565);
  nand n15986(x15986, x15257, x15701);
  nand n15987(x15987, x15986, x15985);
  nand n15988(x15988, x15264, x15704);
  nand n15990(x15990, x15263, x15989);
  nand n15991(x15991, x15990, x15988);
  nand n15992(x15992, x15270, x15707);
  nand n15994(x15994, x15269, x15993);
  nand n15995(x15995, x15994, x15992);
  nand n15996(x15996, x15276, x15710);
  nand n15998(x15998, x15275, x15997);
  nand n15999(x15999, x15998, x15996);
  nand n16000(x16000, x15282, x15713);
  nand n16001(x16001, x15281, x15829);
  nand n16002(x16002, x16001, x16000);
  nand n16003(x16003, x15288, x15832);
  nand n16005(x16005, x15287, x16004);
  nand n16006(x16006, x16005, x16003);
  nand n16007(x16007, x15294, x15835);
  nand n16009(x16009, x15293, x16008);
  nand n16010(x16010, x16009, x16007);
  nand n16011(x16011, x15300, x15838);
  nand n16013(x16013, x15299, x16012);
  nand n16014(x16014, x16013, x16011);
  nand n16015(x16015, x15306, x15841);
  nand n16017(x16017, x15305, x16016);
  nand n16018(x16018, x16017, x16015);
  nand n16019(x16019, x15312, x15844);
  nand n16021(x16021, x15311, x16020);
  nand n16022(x16022, x16021, x16019);
  nand n16023(x16023, x15318, x15847);
  nand n16025(x16025, x15317, x16024);
  nand n16026(x16026, x16025, x16023);
  nand n16027(x16027, x15324, x15850);
  nand n16029(x16029, x15323, x16028);
  nand n16030(x16030, x16029, x16027);
  nand n16031(x16031, x15330, x15853);
  nand n16032(x16032, x15329, x15929);
  nand n16033(x16033, x16032, x16031);
  nand n16034(x16034, x15336, x15932);
  nand n16036(x16036, x15335, x16035);
  nand n16037(x16037, x16036, x16034);
  nand n16038(x16038, x15342, x15935);
  nand n16040(x16040, x15341, x16039);
  nand n16041(x16041, x16040, x16038);
  nand n16042(x16042, x15348, x15938);
  nand n16044(x16044, x15347, x16043);
  nand n16045(x16045, x16044, x16042);
  nand n16046(x16046, x15354, x15941);
  nand n16048(x16048, x15353, x16047);
  nand n16049(x16049, x16048, x16046);
  nand n16050(x16050, x15360, x15944);
  nand n16052(x16052, x15359, x16051);
  nand n16053(x16053, x16052, x16050);
  nand n16054(x16054, x15365, x15947);
  nand n16056(x16056, x15364, x16055);
  nand n16057(x16057, x16056, x16054);
  nand n16058(x16058, x15370, x15950);
  nand n16060(x16060, x15369, x16059);
  nand n16061(x16061, x16060, x16058);
  nand n16062(x16062, x15375, x15953);
  nand n16064(x16064, x15374, x16063);
  nand n16065(x16065, x16064, x16062);
  nand n16066(x16066, x15380, x15956);
  nand n16068(x16068, x15379, x16067);
  nand n16069(x16069, x16068, x16066);
  nand n16070(x16070, x15385, x15959);
  nand n16072(x16072, x15384, x16071);
  nand n16073(x16073, x16072, x16070);
  nand n16074(x16074, x15390, x15962);
  nand n16076(x16076, x15389, x16075);
  nand n16077(x16077, x16076, x16074);
  nand n16078(x16078, x15395, x15965);
  nand n16080(x16080, x15394, x16079);
  nand n16081(x16081, x16080, x16078);
  nand n16082(x16082, x15400, x15968);
  nand n16084(x16084, x15399, x16083);
  nand n16085(x16085, x16084, x16082);
  nand n16086(x16086, x15405, x15971);
  nand n16088(x16088, x15404, x16087);
  nand n16089(x16089, x16088, x16086);
  nand n16090(x16090, x15410, x15974);
  nand n16092(x16092, x15409, x16091);
  nand n16093(x16093, x16092, x16090);
  nand n16094(x16094, x83516, x15980);
  nand n16095(x16095, x83517, x83516);
  nand n16097(x16097, x83518, x83517);
  nand n16099(x16099, x83519, x83518);
  nand n16101(x16101, x83520, x83519);
  nand n16103(x16103, x83521, x83520);
  nand n16105(x16105, x83522, x83521);
  nand n16107(x16107, x83523, x83522);
  nand n16109(x16109, x83524, x83523);
  nand n16111(x16111, x83525, x83524);
  nand n16113(x16113, x83526, x83525);
  nand n16115(x16115, x83527, x83526);
  nand n16117(x16117, x83528, x83527);
  nand n16119(x16119, x83529, x83528);
  nand n16121(x16121, x83530, x83529);
  nand n16123(x16123, x83531, x83530);
  nand n16125(x16125, x83532, x83531);
  nand n16127(x16127, x83533, x83532);
  nand n16129(x16129, x83534, x83533);
  nand n16131(x16131, x83535, x83534);
  nand n16133(x16133, x83536, x83535);
  nand n16135(x16135, x83537, x83536);
  nand n16137(x16137, x83538, x83537);
  nand n16139(x16139, x83539, x83538);
  nand n16141(x16141, x83540, x83539);
  nand n16143(x16143, x83541, x83540);
  nand n16145(x16145, x83542, x83541);
  nand n16147(x16147, x83543, x83542);
  nand n16149(x16149, x16096, x15980);
  nand n16150(x16150, x16098, x83545);
  nand n16151(x16151, x16100, x16096);
  nand n16153(x16153, x16102, x16098);
  nand n16155(x16155, x16104, x16100);
  nand n16157(x16157, x16106, x16102);
  nand n16159(x16159, x16108, x16104);
  nand n16161(x16161, x16110, x16106);
  nand n16163(x16163, x16112, x16108);
  nand n16165(x16165, x16114, x16110);
  nand n16167(x16167, x16116, x16112);
  nand n16169(x16169, x16118, x16114);
  nand n16171(x16171, x16120, x16116);
  nand n16173(x16173, x16122, x16118);
  nand n16175(x16175, x16124, x16120);
  nand n16177(x16177, x16126, x16122);
  nand n16179(x16179, x16128, x16124);
  nand n16181(x16181, x16130, x16126);
  nand n16183(x16183, x16132, x16128);
  nand n16185(x16185, x16134, x16130);
  nand n16187(x16187, x16136, x16132);
  nand n16189(x16189, x16138, x16134);
  nand n16191(x16191, x16140, x16136);
  nand n16193(x16193, x16142, x16138);
  nand n16195(x16195, x16144, x16140);
  nand n16197(x16197, x16146, x16142);
  nand n16199(x16199, x16148, x16144);
  nand n16201(x16201, x16152, x15980);
  nand n16202(x16202, x16154, x83545);
  nand n16203(x16203, x16156, x83546);
  nand n16204(x16204, x16158, x83547);
  nand n16205(x16205, x16160, x16152);
  nand n16207(x16207, x16162, x16154);
  nand n16209(x16209, x16164, x16156);
  nand n16211(x16211, x16166, x16158);
  nand n16213(x16213, x16168, x16160);
  nand n16215(x16215, x16170, x16162);
  nand n16217(x16217, x16172, x16164);
  nand n16219(x16219, x16174, x16166);
  nand n16221(x16221, x16176, x16168);
  nand n16223(x16223, x16178, x16170);
  nand n16225(x16225, x16180, x16172);
  nand n16227(x16227, x16182, x16174);
  nand n16229(x16229, x16184, x16176);
  nand n16231(x16231, x16186, x16178);
  nand n16233(x16233, x16188, x16180);
  nand n16235(x16235, x16190, x16182);
  nand n16237(x16237, x16192, x16184);
  nand n16239(x16239, x16194, x16186);
  nand n16241(x16241, x16196, x16188);
  nand n16243(x16243, x16198, x16190);
  nand n16245(x16245, x16200, x16192);
  nand n16247(x16247, x16206, x15980);
  nand n16248(x16248, x16208, x83545);
  nand n16249(x16249, x16210, x83546);
  nand n16250(x16250, x16212, x83547);
  nand n16251(x16251, x16214, x83548);
  nand n16252(x16252, x16216, x83549);
  nand n16253(x16253, x16218, x83550);
  nand n16254(x16254, x16220, x83551);
  nand n16255(x16255, x16222, x16206);
  nand n16257(x16257, x16224, x16208);
  nand n16259(x16259, x16226, x16210);
  nand n16261(x16261, x16228, x16212);
  nand n16263(x16263, x16230, x16214);
  nand n16265(x16265, x16232, x16216);
  nand n16267(x16267, x16234, x16218);
  nand n16269(x16269, x16236, x16220);
  nand n16271(x16271, x16238, x16222);
  nand n16273(x16273, x16240, x16224);
  nand n16275(x16275, x16242, x16226);
  nand n16277(x16277, x16244, x16228);
  nand n16279(x16279, x16246, x16230);
  nand n16281(x16281, x16256, x15980);
  nand n16282(x16282, x16258, x83545);
  nand n16283(x16283, x16260, x83546);
  nand n16284(x16284, x16262, x83547);
  nand n16285(x16285, x16264, x83548);
  nand n16286(x16286, x16266, x83549);
  nand n16287(x16287, x16268, x83550);
  nand n16288(x16288, x16270, x83551);
  nand n16289(x16289, x16272, x83552);
  nand n16290(x16290, x16274, x83553);
  nand n16291(x16291, x16276, x83554);
  nand n16292(x16292, x16278, x83555);
  nand n16293(x16293, x16280, x83556);
  nand n16294(x16294, x15984, x15979);
  nand n16295(x16295, x16294, x16094);
  nand n16297(x16297, x83517, x83545);
  nand n16298(x16298, x15987, x16094);
  nand n16299(x16299, x16298, x16297);
  nand n16301(x16301, x83518, x83546);
  nand n16302(x16302, x15991, x16149);
  nand n16303(x16303, x16302, x16301);
  nand n16305(x16305, x83519, x83547);
  nand n16306(x16306, x15995, x16150);
  nand n16307(x16307, x16306, x16305);
  nand n16309(x16309, x83520, x83548);
  nand n16310(x16310, x15999, x16201);
  nand n16311(x16311, x16310, x16309);
  nand n16313(x16313, x83521, x83549);
  nand n16314(x16314, x16002, x16202);
  nand n16315(x16315, x16314, x16313);
  nand n16317(x16317, x83522, x83550);
  nand n16318(x16318, x16006, x16203);
  nand n16319(x16319, x16318, x16317);
  nand n16321(x16321, x83523, x83551);
  nand n16322(x16322, x16010, x16204);
  nand n16323(x16323, x16322, x16321);
  nand n16325(x16325, x83524, x83552);
  nand n16326(x16326, x16014, x16247);
  nand n16327(x16327, x16326, x16325);
  nand n16329(x16329, x83525, x83553);
  nand n16330(x16330, x16018, x16248);
  nand n16331(x16331, x16330, x16329);
  nand n16333(x16333, x83526, x83554);
  nand n16334(x16334, x16022, x16249);
  nand n16335(x16335, x16334, x16333);
  nand n16337(x16337, x83527, x83555);
  nand n16338(x16338, x16026, x16250);
  nand n16339(x16339, x16338, x16337);
  nand n16341(x16341, x83528, x83556);
  nand n16342(x16342, x16030, x16251);
  nand n16343(x16343, x16342, x16341);
  nand n16345(x16345, x83529, x83557);
  nand n16346(x16346, x16033, x16252);
  nand n16347(x16347, x16346, x16345);
  nand n16349(x16349, x83530, x83558);
  nand n16350(x16350, x16037, x16253);
  nand n16351(x16351, x16350, x16349);
  nand n16353(x16353, x83531, x83559);
  nand n16354(x16354, x16041, x16254);
  nand n16355(x16355, x16354, x16353);
  nand n16357(x16357, x83532, x83560);
  nand n16358(x16358, x16045, x16281);
  nand n16359(x16359, x16358, x16357);
  nand n16361(x16361, x83533, x83561);
  nand n16362(x16362, x16049, x16282);
  nand n16363(x16363, x16362, x16361);
  nand n16365(x16365, x83534, x83562);
  nand n16366(x16366, x16053, x16283);
  nand n16367(x16367, x16366, x16365);
  nand n16369(x16369, x83535, x83563);
  nand n16370(x16370, x16057, x16284);
  nand n16371(x16371, x16370, x16369);
  nand n16373(x16373, x83536, x83564);
  nand n16374(x16374, x16061, x16285);
  nand n16375(x16375, x16374, x16373);
  nand n16377(x16377, x83537, x83565);
  nand n16378(x16378, x16065, x16286);
  nand n16379(x16379, x16378, x16377);
  nand n16381(x16381, x83538, x83566);
  nand n16382(x16382, x16069, x16287);
  nand n16383(x16383, x16382, x16381);
  nand n16385(x16385, x83539, x83567);
  nand n16386(x16386, x16073, x16288);
  nand n16387(x16387, x16386, x16385);
  nand n16389(x16389, x83540, x83568);
  nand n16390(x16390, x16077, x16289);
  nand n16391(x16391, x16390, x16389);
  nand n16393(x16393, x83541, x83569);
  nand n16394(x16394, x16081, x16290);
  nand n16395(x16395, x16394, x16393);
  nand n16397(x16397, x83542, x83570);
  nand n16398(x16398, x16085, x16291);
  nand n16399(x16399, x16398, x16397);
  nand n16401(x16401, x83543, x83571);
  nand n16402(x16402, x16089, x16292);
  nand n16403(x16403, x16402, x16401);
  nand n16405(x16405, x83544, x83572);
  nand n16406(x16406, x16093, x16293);
  nand n16407(x16407, x16406, x16405);
  nand n16409(x16409, x15220, x83573);
  nand n16411(x16411, x16410, x6503);
  nand n16412(x16412, x16411, x16409);
  nand n16413(x16413, x15220, x83574);
  nand n16414(x16414, x16410, x6524);
  nand n16415(x16415, x16414, x16413);
  nand n16416(x16416, x15220, x15979);
  nand n16417(x16417, x16410, x6545);
  nand n16418(x16418, x16417, x16416);
  nand n16419(x16419, x15220, x16296);
  nand n16420(x16420, x16410, x6566);
  nand n16421(x16421, x16420, x16419);
  nand n16422(x16422, x15220, x16300);
  nand n16423(x16423, x16410, x6587);
  nand n16424(x16424, x16423, x16422);
  nand n16425(x16425, x15220, x16304);
  nand n16426(x16426, x16410, x6608);
  nand n16427(x16427, x16426, x16425);
  nand n16428(x16428, x15220, x16308);
  nand n16429(x16429, x16410, x6629);
  nand n16430(x16430, x16429, x16428);
  nand n16431(x16431, x15220, x16312);
  nand n16432(x16432, x16410, x6650);
  nand n16433(x16433, x16432, x16431);
  nand n16434(x16434, x15220, x16316);
  nand n16435(x16435, x16410, x6671);
  nand n16436(x16436, x16435, x16434);
  nand n16437(x16437, x15220, x16320);
  nand n16438(x16438, x16410, x6692);
  nand n16439(x16439, x16438, x16437);
  nand n16440(x16440, x15220, x16324);
  nand n16441(x16441, x16410, x6713);
  nand n16442(x16442, x16441, x16440);
  nand n16443(x16443, x15220, x16328);
  nand n16444(x16444, x16410, x6734);
  nand n16445(x16445, x16444, x16443);
  nand n16446(x16446, x15220, x16332);
  nand n16447(x16447, x16410, x6755);
  nand n16448(x16448, x16447, x16446);
  nand n16449(x16449, x15220, x16336);
  nand n16450(x16450, x16410, x6776);
  nand n16451(x16451, x16450, x16449);
  nand n16452(x16452, x15220, x16340);
  nand n16453(x16453, x16410, x6797);
  nand n16454(x16454, x16453, x16452);
  nand n16455(x16455, x15220, x16344);
  nand n16456(x16456, x16410, x6818);
  nand n16457(x16457, x16456, x16455);
  nand n16458(x16458, x15220, x16348);
  nand n16459(x16459, x16410, x6839);
  nand n16460(x16460, x16459, x16458);
  nand n16461(x16461, x15220, x16352);
  nand n16462(x16462, x16410, x6860);
  nand n16463(x16463, x16462, x16461);
  nand n16464(x16464, x15220, x16356);
  nand n16465(x16465, x16410, x6881);
  nand n16466(x16466, x16465, x16464);
  nand n16467(x16467, x15220, x16360);
  nand n16468(x16468, x16410, x6902);
  nand n16469(x16469, x16468, x16467);
  nand n16470(x16470, x15220, x16364);
  nand n16471(x16471, x16410, x6923);
  nand n16472(x16472, x16471, x16470);
  nand n16473(x16473, x15220, x16368);
  nand n16474(x16474, x16410, x6944);
  nand n16475(x16475, x16474, x16473);
  nand n16476(x16476, x15220, x16372);
  nand n16477(x16477, x16410, x6965);
  nand n16478(x16478, x16477, x16476);
  nand n16479(x16479, x15220, x16376);
  nand n16480(x16480, x16410, x6986);
  nand n16481(x16481, x16480, x16479);
  nand n16482(x16482, x15220, x16380);
  nand n16483(x16483, x16410, x7007);
  nand n16484(x16484, x16483, x16482);
  nand n16485(x16485, x15220, x16384);
  nand n16486(x16486, x16410, x7028);
  nand n16487(x16487, x16486, x16485);
  nand n16488(x16488, x15220, x16388);
  nand n16489(x16489, x16410, x7049);
  nand n16490(x16490, x16489, x16488);
  nand n16491(x16491, x15220, x16392);
  nand n16492(x16492, x16410, x7070);
  nand n16493(x16493, x16492, x16491);
  nand n16494(x16494, x15220, x16396);
  nand n16495(x16495, x16410, x7091);
  nand n16496(x16496, x16495, x16494);
  nand n16497(x16497, x15220, x16400);
  nand n16498(x16498, x16410, x7112);
  nand n16499(x16499, x16498, x16497);
  nand n16500(x16500, x15220, x16404);
  nand n16501(x16501, x16410, x7133);
  nand n16502(x16502, x16501, x16500);
  nand n16503(x16503, x15220, x16408);
  nand n16504(x16504, x16410, x7154);
  nand n16505(x16505, x16504, x16503);
  nand n16506(x16506, x1696, x1698);
  nand n16507(x16507, x1692, x1694);
  nand n16510(x16510, x16509, x16508);
  nand n16511(x16511, x1001, x16510);
  nand n16513(x16513, x71270, x16510);
  nand n16515(x16515, x1038, x16512);
  nand n16517(x16517, x71265, x16512);
  nand n16519(x16519, x1038, x16514);
  nand n16521(x16521, x71265, x16514);
  nand n16523(x16523, x1022, x16516);
  nand n16525(x16525, x71260, x16516);
  nand n16527(x16527, x1022, x16518);
  nand n16529(x16529, x71260, x16518);
  nand n16531(x16531, x1022, x16520);
  nand n16533(x16533, x71260, x16520);
  nand n16535(x16535, x1022, x16522);
  nand n16537(x16537, x71260, x16522);
  nand n16539(x16539, x71255, x16524);
  nand n16541(x16541, x1012, x16526);
  nand n16543(x16543, x71255, x16526);
  nand n16545(x16545, x1012, x16528);
  nand n16547(x16547, x71255, x16528);
  nand n16549(x16549, x1012, x16530);
  nand n16551(x16551, x71255, x16530);
  nand n16553(x16553, x1012, x16532);
  nand n16555(x16555, x71255, x16532);
  nand n16557(x16557, x1012, x16534);
  nand n16559(x16559, x71255, x16534);
  nand n16561(x16561, x1012, x16536);
  nand n16563(x16563, x71255, x16536);
  nand n16565(x16565, x1012, x16538);
  nand n16567(x16567, x1011, x16540);
  nand n16569(x16569, x71250, x16540);
  nand n16571(x16571, x1011, x16542);
  nand n16573(x16573, x71250, x16542);
  nand n16575(x16575, x1011, x16544);
  nand n16577(x16577, x71250, x16544);
  nand n16579(x16579, x1011, x16546);
  nand n16581(x16581, x71250, x16546);
  nand n16583(x16583, x1011, x16548);
  nand n16585(x16585, x71250, x16548);
  nand n16587(x16587, x1011, x16550);
  nand n16589(x16589, x71250, x16550);
  nand n16591(x16591, x1011, x16552);
  nand n16593(x16593, x71250, x16554);
  nand n16595(x16595, x1011, x16556);
  nand n16597(x16597, x71250, x16556);
  nand n16599(x16599, x1011, x16558);
  nand n16601(x16601, x71250, x16558);
  nand n16603(x16603, x1011, x16560);
  nand n16605(x16605, x71250, x16562);
  nand n16607(x16607, x1011, x16564);
  nand n16609(x16609, x71250, x16564);
  nand n16611(x16611, x1011, x16566);
  nand n16613(x16613, x71245, x16568);
  nand n16614(x16614, x1000, x16570);
  nand n16615(x16615, x71245, x16570);
  nand n16616(x16616, x1000, x16572);
  nand n16617(x16617, x71245, x16572);
  nand n16618(x16618, x1000, x16574);
  nand n16619(x16619, x71245, x16574);
  nand n16620(x16620, x1000, x16576);
  nand n16621(x16621, x71245, x16576);
  nand n16622(x16622, x1000, x16578);
  nand n16623(x16623, x71245, x16578);
  nand n16624(x16624, x1000, x16580);
  nand n16625(x16625, x71245, x16580);
  nand n16626(x16626, x1000, x16582);
  nand n16627(x16627, x71245, x16582);
  nand n16628(x16628, x1000, x16584);
  nand n16629(x16629, x71245, x16584);
  nand n16630(x16630, x1000, x16586);
  nand n16631(x16631, x71245, x16586);
  nand n16632(x16632, x1000, x16588);
  nand n16633(x16633, x71245, x16588);
  nand n16634(x16634, x1000, x16590);
  nand n16635(x16635, x71245, x16590);
  nand n16636(x16636, x1000, x16592);
  nand n16637(x16637, x71245, x16594);
  nand n16638(x16638, x1000, x16596);
  nand n16639(x16639, x71245, x16596);
  nand n16640(x16640, x1000, x16598);
  nand n16641(x16641, x71245, x16598);
  nand n16642(x16642, x1000, x16600);
  nand n16643(x16643, x71245, x16600);
  nand n16644(x16644, x1000, x16602);
  nand n16645(x16645, x71245, x16602);
  nand n16646(x16646, x1000, x16604);
  nand n16647(x16647, x71245, x16606);
  nand n16648(x16648, x1000, x16608);
  nand n16649(x16649, x71245, x16608);
  nand n16650(x16650, x1000, x16610);
  nand n16651(x16651, x71245, x16610);
  nand n16652(x16652, x1000, x16612);
  nand n16653(x16653, x71245, x16612);
  nand n16654(x16654, x14561, x1718);
  nand n16655(x16655, x14562, x1719);
  nand n16656(x16656, x14563, x1720);
  nand n16657(x16657, x14564, x1721);
  nand n16660(x16660, x16659, x16658);
  nand n16663(x16663, x16662, x16661);
  nand n16666(x16666, x16665, x16664);
  nand n16668(x16668, x16667, x1143);
  nand n16669(x16669, x16613, x16614);
  nand n16670(x16670, x16615, x16616);
  nand n16671(x16671, x16617, x16618);
  nand n16672(x16672, x16619, x16620);
  nand n16673(x16673, x16623, x16624);
  nand n16674(x16674, x16625, x16626);
  nand n16675(x16675, x16627, x16628);
  nand n16676(x16676, x16629, x16630);
  nand n16677(x16677, x16633, x16634);
  nand n16678(x16678, x16635, x16636);
  nand n16681(x16681, x16680, x16679);
  nand n16684(x16684, x16683, x16682);
  nand n16687(x16687, x16686, x16685);
  nand n16690(x16690, x16689, x16688);
  nand n16693(x16693, x16692, x16691);
  nand n16696(x16696, x16695, x16694);
  nand n16699(x16699, x16698, x16697);
  nand n16701(x16701, x16700, x16639);
  nand n16704(x16704, x16703, x16702);
  nand n16707(x16707, x16706, x16705);
  nand n16708(x16708, x16707, x16668);
  nand n16710(x16710, x16640, x16641);
  nand n16711(x16711, x16642, x16643);
  nand n16712(x16712, x16644, x16645);
  nand n16715(x16715, x16714, x16713);
  nand n16717(x16717, x16716, x16646);
  nand n16720(x16720, x16719, x16718);
  nand n16721(x16721, x16720, x16668);
  nand n16723(x16723, x16621, x16622);
  nand n16724(x16724, x16631, x16632);
  nand n16727(x16727, x16726, x16725);
  nand n16728(x16728, x16727, x16668);
  nand n16730(x16730, x16637, x16638);
  nand n16731(x16731, x16730, x16668);
  nand n16733(x16733, x16647, x16648);
  nand n16734(x16734, x16649, x16650);
  nand n16737(x16737, x16736, x16735);
  nand n16739(x16739, x16738, x16653);
  nand n16740(x16740, x16739, x16668);
  nand n16742(x16742, x16651, x16652);
  nand n16743(x16743, x16742, x16668);
  nand n16746(x16746, x71942, x71802);
  nand n16748(x16748, x16747, x72207);
  nand n16749(x16749, x16748, x16746);
  nand n16750(x16750, x71942, x71807);
  nand n16751(x16751, x16747, x72212);
  nand n16752(x16752, x16751, x16750);
  nand n16753(x16753, x71942, x71812);
  nand n16754(x16754, x16747, x72217);
  nand n16755(x16755, x16754, x16753);
  nand n16756(x16756, x71942, x71817);
  nand n16757(x16757, x16747, x72222);
  nand n16758(x16758, x16757, x16756);
  nand n16759(x16759, x71942, x71822);
  nand n16760(x16760, x16747, x72227);
  nand n16761(x16761, x16760, x16759);
  nand n16762(x16762, x71942, x71827);
  nand n16763(x16763, x16747, x72232);
  nand n16764(x16764, x16763, x16762);
  nand n16765(x16765, x71942, x71832);
  nand n16766(x16766, x16747, x72237);
  nand n16767(x16767, x16766, x16765);
  nand n16768(x16768, x71942, x71837);
  nand n16769(x16769, x16747, x72242);
  nand n16770(x16770, x16769, x16768);
  nand n16771(x16771, x71942, x71842);
  nand n16772(x16772, x16747, x72247);
  nand n16773(x16773, x16772, x16771);
  nand n16774(x16774, x71942, x71847);
  nand n16775(x16775, x16747, x72252);
  nand n16776(x16776, x16775, x16774);
  nand n16777(x16777, x71942, x71852);
  nand n16778(x16778, x16747, x72257);
  nand n16779(x16779, x16778, x16777);
  nand n16780(x16780, x71942, x71857);
  nand n16781(x16781, x16747, x72262);
  nand n16782(x16782, x16781, x16780);
  nand n16783(x16783, x71942, x71862);
  nand n16784(x16784, x16747, x72267);
  nand n16785(x16785, x16784, x16783);
  nand n16786(x16786, x71942, x71867);
  nand n16787(x16787, x16747, x72272);
  nand n16788(x16788, x16787, x16786);
  nand n16789(x16789, x71942, x71872);
  nand n16790(x16790, x16747, x72277);
  nand n16791(x16791, x16790, x16789);
  nand n16792(x16792, x71942, x71877);
  nand n16793(x16793, x16747, x72282);
  nand n16794(x16794, x16793, x16792);
  nand n16795(x16795, x71942, x71882);
  nand n16796(x16796, x16747, x72287);
  nand n16797(x16797, x16796, x16795);
  nand n16798(x16798, x71942, x71887);
  nand n16799(x16799, x16747, x72292);
  nand n16800(x16800, x16799, x16798);
  nand n16801(x16801, x71942, x71892);
  nand n16802(x16802, x16747, x72297);
  nand n16803(x16803, x16802, x16801);
  nand n16804(x16804, x71942, x71897);
  nand n16805(x16805, x16747, x72302);
  nand n16806(x16806, x16805, x16804);
  nand n16807(x16807, x71942, x71902);
  nand n16808(x16808, x16747, x72307);
  nand n16809(x16809, x16808, x16807);
  nand n16810(x16810, x71942, x71907);
  nand n16811(x16811, x16747, x72312);
  nand n16812(x16812, x16811, x16810);
  nand n16813(x16813, x71942, x71910);
  nand n16814(x16814, x16747, x72317);
  nand n16815(x16815, x16814, x16813);
  nand n16816(x16816, x71942, x71913);
  nand n16817(x16817, x16747, x72322);
  nand n16818(x16818, x16817, x16816);
  nand n16819(x16819, x71942, x71916);
  nand n16820(x16820, x16747, x72327);
  nand n16821(x16821, x16820, x16819);
  nand n16822(x16822, x71942, x71919);
  nand n16823(x16823, x16747, x72332);
  nand n16824(x16824, x16823, x16822);
  nand n16825(x16825, x71942, x71922);
  nand n16826(x16826, x16747, x72337);
  nand n16827(x16827, x16826, x16825);
  nand n16828(x16828, x71942, x71925);
  nand n16829(x16829, x16747, x72342);
  nand n16830(x16830, x16829, x16828);
  nand n16831(x16831, x71942, x71928);
  nand n16832(x16832, x16747, x72347);
  nand n16833(x16833, x16832, x16831);
  nand n16834(x16834, x71942, x71931);
  nand n16835(x16835, x16747, x72352);
  nand n16836(x16836, x16835, x16834);
  nand n16837(x16837, x71942, x71934);
  nand n16838(x16838, x16747, x72357);
  nand n16839(x16839, x16838, x16837);
  nand n16840(x16840, x71942, x71937);
  nand n16841(x16841, x16747, x72362);
  nand n16842(x16842, x16841, x16840);
  nand n16875(x16875, x71977, x16843);
  nand n16877(x16877, x16876, x16749);
  nand n16878(x16878, x16877, x16875);
  nand n16879(x16879, x71977, x16844);
  nand n16880(x16880, x16876, x16752);
  nand n16881(x16881, x16880, x16879);
  nand n16882(x16882, x71977, x16845);
  nand n16883(x16883, x16876, x16755);
  nand n16884(x16884, x16883, x16882);
  nand n16885(x16885, x71977, x16846);
  nand n16886(x16886, x16876, x16758);
  nand n16887(x16887, x16886, x16885);
  nand n16888(x16888, x71977, x16847);
  nand n16889(x16889, x16876, x16761);
  nand n16890(x16890, x16889, x16888);
  nand n16891(x16891, x71977, x16848);
  nand n16892(x16892, x16876, x16764);
  nand n16893(x16893, x16892, x16891);
  nand n16894(x16894, x71977, x16849);
  nand n16895(x16895, x16876, x16767);
  nand n16896(x16896, x16895, x16894);
  nand n16897(x16897, x71977, x16850);
  nand n16898(x16898, x16876, x16770);
  nand n16899(x16899, x16898, x16897);
  nand n16900(x16900, x71977, x16851);
  nand n16901(x16901, x16876, x16773);
  nand n16902(x16902, x16901, x16900);
  nand n16903(x16903, x71977, x16852);
  nand n16904(x16904, x16876, x16776);
  nand n16905(x16905, x16904, x16903);
  nand n16906(x16906, x71977, x16853);
  nand n16907(x16907, x16876, x16779);
  nand n16908(x16908, x16907, x16906);
  nand n16909(x16909, x71977, x16854);
  nand n16910(x16910, x16876, x16782);
  nand n16911(x16911, x16910, x16909);
  nand n16912(x16912, x71977, x16855);
  nand n16913(x16913, x16876, x16785);
  nand n16914(x16914, x16913, x16912);
  nand n16915(x16915, x71977, x16856);
  nand n16916(x16916, x16876, x16788);
  nand n16917(x16917, x16916, x16915);
  nand n16918(x16918, x71977, x16857);
  nand n16919(x16919, x16876, x16791);
  nand n16920(x16920, x16919, x16918);
  nand n16921(x16921, x71977, x16858);
  nand n16922(x16922, x16876, x16794);
  nand n16923(x16923, x16922, x16921);
  nand n16924(x16924, x71977, x16859);
  nand n16925(x16925, x16876, x16797);
  nand n16926(x16926, x16925, x16924);
  nand n16927(x16927, x71977, x16860);
  nand n16928(x16928, x16876, x16800);
  nand n16929(x16929, x16928, x16927);
  nand n16930(x16930, x71977, x16861);
  nand n16931(x16931, x16876, x16803);
  nand n16932(x16932, x16931, x16930);
  nand n16933(x16933, x71977, x16862);
  nand n16934(x16934, x16876, x16806);
  nand n16935(x16935, x16934, x16933);
  nand n16936(x16936, x71977, x16863);
  nand n16937(x16937, x16876, x16809);
  nand n16938(x16938, x16937, x16936);
  nand n16939(x16939, x71977, x16864);
  nand n16940(x16940, x16876, x16812);
  nand n16941(x16941, x16940, x16939);
  nand n16942(x16942, x71977, x16865);
  nand n16943(x16943, x16876, x16815);
  nand n16944(x16944, x16943, x16942);
  nand n16945(x16945, x71977, x16866);
  nand n16946(x16946, x16876, x16818);
  nand n16947(x16947, x16946, x16945);
  nand n16948(x16948, x71977, x16867);
  nand n16949(x16949, x16876, x16821);
  nand n16950(x16950, x16949, x16948);
  nand n16951(x16951, x71977, x16868);
  nand n16952(x16952, x16876, x16824);
  nand n16953(x16953, x16952, x16951);
  nand n16954(x16954, x71977, x16869);
  nand n16955(x16955, x16876, x16827);
  nand n16956(x16956, x16955, x16954);
  nand n16957(x16957, x71977, x16870);
  nand n16958(x16958, x16876, x16830);
  nand n16959(x16959, x16958, x16957);
  nand n16960(x16960, x71977, x16871);
  nand n16961(x16961, x16876, x16833);
  nand n16962(x16962, x16961, x16960);
  nand n16963(x16963, x71977, x16872);
  nand n16964(x16964, x16876, x16836);
  nand n16965(x16965, x16964, x16963);
  nand n16966(x16966, x71977, x16873);
  nand n16967(x16967, x16876, x16839);
  nand n16968(x16968, x16967, x16966);
  nand n16969(x16969, x71977, x16874);
  nand n16970(x16970, x16876, x16842);
  nand n16971(x16971, x16970, x16969);
  nand n16972(x16972, x72047, x16878);
  nand n16975(x16975, x16974, x16973);
  nand n16976(x16976, x16975, x16972);
  nand n16978(x16978, x72052, x16881);
  nand n16981(x16981, x16980, x16979);
  nand n16982(x16982, x16981, x16978);
  nand n16984(x16984, x72057, x16884);
  nand n16987(x16987, x16986, x16985);
  nand n16988(x16988, x16987, x16984);
  nand n16990(x16990, x72062, x16887);
  nand n16993(x16993, x16992, x16991);
  nand n16994(x16994, x16993, x16990);
  nand n16996(x16996, x72067, x16890);
  nand n16999(x16999, x16998, x16997);
  nand n17000(x17000, x16999, x16996);
  nand n17002(x17002, x72072, x16893);
  nand n17005(x17005, x17004, x17003);
  nand n17006(x17006, x17005, x17002);
  nand n17008(x17008, x72077, x16896);
  nand n17011(x17011, x17010, x17009);
  nand n17012(x17012, x17011, x17008);
  nand n17014(x17014, x72082, x16899);
  nand n17017(x17017, x17016, x17015);
  nand n17018(x17018, x17017, x17014);
  nand n17020(x17020, x72087, x16902);
  nand n17023(x17023, x17022, x17021);
  nand n17024(x17024, x17023, x17020);
  nand n17026(x17026, x72092, x16905);
  nand n17029(x17029, x17028, x17027);
  nand n17030(x17030, x17029, x17026);
  nand n17032(x17032, x72097, x16908);
  nand n17035(x17035, x17034, x17033);
  nand n17036(x17036, x17035, x17032);
  nand n17038(x17038, x72102, x16911);
  nand n17041(x17041, x17040, x17039);
  nand n17042(x17042, x17041, x17038);
  nand n17044(x17044, x72107, x16914);
  nand n17047(x17047, x17046, x17045);
  nand n17048(x17048, x17047, x17044);
  nand n17050(x17050, x72112, x16917);
  nand n17053(x17053, x17052, x17051);
  nand n17054(x17054, x17053, x17050);
  nand n17056(x17056, x72117, x16920);
  nand n17059(x17059, x17058, x17057);
  nand n17060(x17060, x17059, x17056);
  nand n17062(x17062, x72122, x16923);
  nand n17065(x17065, x17064, x17063);
  nand n17066(x17066, x17065, x17062);
  nand n17068(x17068, x72127, x16926);
  nand n17071(x17071, x17070, x17069);
  nand n17072(x17072, x17071, x17068);
  nand n17074(x17074, x72132, x16929);
  nand n17077(x17077, x17076, x17075);
  nand n17078(x17078, x17077, x17074);
  nand n17080(x17080, x72137, x16932);
  nand n17083(x17083, x17082, x17081);
  nand n17084(x17084, x17083, x17080);
  nand n17086(x17086, x72142, x16935);
  nand n17089(x17089, x17088, x17087);
  nand n17090(x17090, x17089, x17086);
  nand n17092(x17092, x72147, x16938);
  nand n17095(x17095, x17094, x17093);
  nand n17096(x17096, x17095, x17092);
  nand n17098(x17098, x72152, x16941);
  nand n17101(x17101, x17100, x17099);
  nand n17102(x17102, x17101, x17098);
  nand n17104(x17104, x72157, x16944);
  nand n17107(x17107, x17106, x17105);
  nand n17108(x17108, x17107, x17104);
  nand n17110(x17110, x72162, x16947);
  nand n17113(x17113, x17112, x17111);
  nand n17114(x17114, x17113, x17110);
  nand n17116(x17116, x72167, x16950);
  nand n17119(x17119, x17118, x17117);
  nand n17120(x17120, x17119, x17116);
  nand n17122(x17122, x72172, x16953);
  nand n17125(x17125, x17124, x17123);
  nand n17126(x17126, x17125, x17122);
  nand n17128(x17128, x72177, x16956);
  nand n17131(x17131, x17130, x17129);
  nand n17132(x17132, x17131, x17128);
  nand n17134(x17134, x72182, x16959);
  nand n17137(x17137, x17136, x17135);
  nand n17138(x17138, x17137, x17134);
  nand n17140(x17140, x72187, x16962);
  nand n17143(x17143, x17142, x17141);
  nand n17144(x17144, x17143, x17140);
  nand n17146(x17146, x72192, x16965);
  nand n17149(x17149, x17148, x17147);
  nand n17150(x17150, x17149, x17146);
  nand n17152(x17152, x72197, x16968);
  nand n17155(x17155, x17154, x17153);
  nand n17156(x17156, x17155, x17152);
  nand n17158(x17158, x72202, x16971);
  nand n17161(x17161, x17160, x17159);
  nand n17162(x17162, x17161, x17158);
  nand n17194(x17194, x16977, x71977);
  nand n17195(x17195, x17194, x16972);
  nand n17196(x17196, x16983, x17164);
  nand n17197(x17197, x17196, x16978);
  nand n17198(x17198, x16983, x16977);
  nand n17200(x17200, x16989, x17165);
  nand n17201(x17201, x17200, x16984);
  nand n17202(x17202, x16989, x16983);
  nand n17204(x17204, x16995, x17166);
  nand n17205(x17205, x17204, x16990);
  nand n17206(x17206, x16995, x16989);
  nand n17208(x17208, x17001, x17167);
  nand n17209(x17209, x17208, x16996);
  nand n17210(x17210, x17001, x16995);
  nand n17212(x17212, x17007, x17168);
  nand n17213(x17213, x17212, x17002);
  nand n17214(x17214, x17007, x17001);
  nand n17216(x17216, x17013, x17169);
  nand n17217(x17217, x17216, x17008);
  nand n17218(x17218, x17013, x17007);
  nand n17220(x17220, x17019, x17170);
  nand n17221(x17221, x17220, x17014);
  nand n17222(x17222, x17019, x17013);
  nand n17224(x17224, x17025, x17171);
  nand n17225(x17225, x17224, x17020);
  nand n17226(x17226, x17025, x17019);
  nand n17228(x17228, x17031, x17172);
  nand n17229(x17229, x17228, x17026);
  nand n17230(x17230, x17031, x17025);
  nand n17232(x17232, x17037, x17173);
  nand n17233(x17233, x17232, x17032);
  nand n17234(x17234, x17037, x17031);
  nand n17236(x17236, x17043, x17174);
  nand n17237(x17237, x17236, x17038);
  nand n17238(x17238, x17043, x17037);
  nand n17240(x17240, x17049, x17175);
  nand n17241(x17241, x17240, x17044);
  nand n17242(x17242, x17049, x17043);
  nand n17244(x17244, x17055, x17176);
  nand n17245(x17245, x17244, x17050);
  nand n17246(x17246, x17055, x17049);
  nand n17248(x17248, x17061, x17177);
  nand n17249(x17249, x17248, x17056);
  nand n17250(x17250, x17061, x17055);
  nand n17252(x17252, x17067, x17178);
  nand n17253(x17253, x17252, x17062);
  nand n17254(x17254, x17067, x17061);
  nand n17256(x17256, x17073, x17179);
  nand n17257(x17257, x17256, x17068);
  nand n17258(x17258, x17073, x17067);
  nand n17260(x17260, x17079, x17180);
  nand n17261(x17261, x17260, x17074);
  nand n17262(x17262, x17079, x17073);
  nand n17264(x17264, x17085, x17181);
  nand n17265(x17265, x17264, x17080);
  nand n17266(x17266, x17085, x17079);
  nand n17268(x17268, x17091, x17182);
  nand n17269(x17269, x17268, x17086);
  nand n17270(x17270, x17091, x17085);
  nand n17272(x17272, x17097, x17183);
  nand n17273(x17273, x17272, x17092);
  nand n17274(x17274, x17097, x17091);
  nand n17276(x17276, x17103, x17184);
  nand n17277(x17277, x17276, x17098);
  nand n17278(x17278, x17103, x17097);
  nand n17280(x17280, x17109, x17185);
  nand n17281(x17281, x17280, x17104);
  nand n17282(x17282, x17109, x17103);
  nand n17284(x17284, x17115, x17186);
  nand n17285(x17285, x17284, x17110);
  nand n17286(x17286, x17115, x17109);
  nand n17288(x17288, x17121, x17187);
  nand n17289(x17289, x17288, x17116);
  nand n17290(x17290, x17121, x17115);
  nand n17292(x17292, x17127, x17188);
  nand n17293(x17293, x17292, x17122);
  nand n17294(x17294, x17127, x17121);
  nand n17296(x17296, x17133, x17189);
  nand n17297(x17297, x17296, x17128);
  nand n17298(x17298, x17133, x17127);
  nand n17300(x17300, x17139, x17190);
  nand n17301(x17301, x17300, x17134);
  nand n17302(x17302, x17139, x17133);
  nand n17304(x17304, x17145, x17191);
  nand n17305(x17305, x17304, x17140);
  nand n17306(x17306, x17145, x17139);
  nand n17308(x17308, x17151, x17192);
  nand n17309(x17309, x17308, x17146);
  nand n17310(x17310, x17151, x17145);
  nand n17312(x17312, x17157, x17193);
  nand n17313(x17313, x17312, x17152);
  nand n17314(x17314, x17157, x17151);
  nand n17316(x17316, x17199, x71977);
  nand n17318(x17318, x17316, x17317);
  nand n17319(x17319, x17203, x17195);
  nand n17321(x17321, x17319, x17320);
  nand n17322(x17322, x17207, x17197);
  nand n17324(x17324, x17322, x17323);
  nand n17325(x17325, x17207, x17199);
  nand n17327(x17327, x17211, x17201);
  nand n17329(x17329, x17327, x17328);
  nand n17330(x17330, x17211, x17203);
  nand n17332(x17332, x17215, x17205);
  nand n17334(x17334, x17332, x17333);
  nand n17335(x17335, x17215, x17207);
  nand n17337(x17337, x17219, x17209);
  nand n17339(x17339, x17337, x17338);
  nand n17340(x17340, x17219, x17211);
  nand n17342(x17342, x17223, x17213);
  nand n17344(x17344, x17342, x17343);
  nand n17345(x17345, x17223, x17215);
  nand n17347(x17347, x17227, x17217);
  nand n17349(x17349, x17347, x17348);
  nand n17350(x17350, x17227, x17219);
  nand n17352(x17352, x17231, x17221);
  nand n17354(x17354, x17352, x17353);
  nand n17355(x17355, x17231, x17223);
  nand n17357(x17357, x17235, x17225);
  nand n17359(x17359, x17357, x17358);
  nand n17360(x17360, x17235, x17227);
  nand n17362(x17362, x17239, x17229);
  nand n17364(x17364, x17362, x17363);
  nand n17365(x17365, x17239, x17231);
  nand n17367(x17367, x17243, x17233);
  nand n17369(x17369, x17367, x17368);
  nand n17370(x17370, x17243, x17235);
  nand n17372(x17372, x17247, x17237);
  nand n17374(x17374, x17372, x17373);
  nand n17375(x17375, x17247, x17239);
  nand n17377(x17377, x17251, x17241);
  nand n17379(x17379, x17377, x17378);
  nand n17380(x17380, x17251, x17243);
  nand n17382(x17382, x17255, x17245);
  nand n17384(x17384, x17382, x17383);
  nand n17385(x17385, x17255, x17247);
  nand n17387(x17387, x17259, x17249);
  nand n17389(x17389, x17387, x17388);
  nand n17390(x17390, x17259, x17251);
  nand n17392(x17392, x17263, x17253);
  nand n17394(x17394, x17392, x17393);
  nand n17395(x17395, x17263, x17255);
  nand n17397(x17397, x17267, x17257);
  nand n17399(x17399, x17397, x17398);
  nand n17400(x17400, x17267, x17259);
  nand n17402(x17402, x17271, x17261);
  nand n17404(x17404, x17402, x17403);
  nand n17405(x17405, x17271, x17263);
  nand n17407(x17407, x17275, x17265);
  nand n17409(x17409, x17407, x17408);
  nand n17410(x17410, x17275, x17267);
  nand n17412(x17412, x17279, x17269);
  nand n17414(x17414, x17412, x17413);
  nand n17415(x17415, x17279, x17271);
  nand n17417(x17417, x17283, x17273);
  nand n17419(x17419, x17417, x17418);
  nand n17420(x17420, x17283, x17275);
  nand n17422(x17422, x17287, x17277);
  nand n17424(x17424, x17422, x17423);
  nand n17425(x17425, x17287, x17279);
  nand n17427(x17427, x17291, x17281);
  nand n17429(x17429, x17427, x17428);
  nand n17430(x17430, x17291, x17283);
  nand n17432(x17432, x17295, x17285);
  nand n17434(x17434, x17432, x17433);
  nand n17435(x17435, x17295, x17287);
  nand n17437(x17437, x17299, x17289);
  nand n17439(x17439, x17437, x17438);
  nand n17440(x17440, x17299, x17291);
  nand n17442(x17442, x17303, x17293);
  nand n17444(x17444, x17442, x17443);
  nand n17445(x17445, x17303, x17295);
  nand n17447(x17447, x17307, x17297);
  nand n17449(x17449, x17447, x17448);
  nand n17450(x17450, x17307, x17299);
  nand n17452(x17452, x17311, x17301);
  nand n17454(x17454, x17452, x17453);
  nand n17455(x17455, x17311, x17303);
  nand n17457(x17457, x17315, x17305);
  nand n17459(x17459, x17457, x17458);
  nand n17460(x17460, x17315, x17307);
  nand n17462(x17462, x17326, x71977);
  nand n17464(x17464, x17462, x17463);
  nand n17465(x17465, x17331, x17195);
  nand n17467(x17467, x17465, x17466);
  nand n17468(x17468, x17336, x17318);
  nand n17470(x17470, x17468, x17469);
  nand n17471(x17471, x17341, x17321);
  nand n17473(x17473, x17471, x17472);
  nand n17474(x17474, x17346, x17324);
  nand n17476(x17476, x17474, x17475);
  nand n17477(x17477, x17346, x17326);
  nand n17479(x17479, x17351, x17329);
  nand n17481(x17481, x17479, x17480);
  nand n17482(x17482, x17351, x17331);
  nand n17484(x17484, x17356, x17334);
  nand n17486(x17486, x17484, x17485);
  nand n17487(x17487, x17356, x17336);
  nand n17489(x17489, x17361, x17339);
  nand n17491(x17491, x17489, x17490);
  nand n17492(x17492, x17361, x17341);
  nand n17494(x17494, x17366, x17344);
  nand n17496(x17496, x17494, x17495);
  nand n17497(x17497, x17366, x17346);
  nand n17499(x17499, x17371, x17349);
  nand n17501(x17501, x17499, x17500);
  nand n17502(x17502, x17371, x17351);
  nand n17504(x17504, x17376, x17354);
  nand n17506(x17506, x17504, x17505);
  nand n17507(x17507, x17376, x17356);
  nand n17509(x17509, x17381, x17359);
  nand n17511(x17511, x17509, x17510);
  nand n17512(x17512, x17381, x17361);
  nand n17514(x17514, x17386, x17364);
  nand n17516(x17516, x17514, x17515);
  nand n17517(x17517, x17386, x17366);
  nand n17519(x17519, x17391, x17369);
  nand n17521(x17521, x17519, x17520);
  nand n17522(x17522, x17391, x17371);
  nand n17524(x17524, x17396, x17374);
  nand n17526(x17526, x17524, x17525);
  nand n17527(x17527, x17396, x17376);
  nand n17529(x17529, x17401, x17379);
  nand n17531(x17531, x17529, x17530);
  nand n17532(x17532, x17401, x17381);
  nand n17534(x17534, x17406, x17384);
  nand n17536(x17536, x17534, x17535);
  nand n17537(x17537, x17406, x17386);
  nand n17539(x17539, x17411, x17389);
  nand n17541(x17541, x17539, x17540);
  nand n17542(x17542, x17411, x17391);
  nand n17544(x17544, x17416, x17394);
  nand n17546(x17546, x17544, x17545);
  nand n17547(x17547, x17416, x17396);
  nand n17549(x17549, x17421, x17399);
  nand n17551(x17551, x17549, x17550);
  nand n17552(x17552, x17421, x17401);
  nand n17554(x17554, x17426, x17404);
  nand n17556(x17556, x17554, x17555);
  nand n17557(x17557, x17426, x17406);
  nand n17559(x17559, x17431, x17409);
  nand n17561(x17561, x17559, x17560);
  nand n17562(x17562, x17431, x17411);
  nand n17564(x17564, x17436, x17414);
  nand n17566(x17566, x17564, x17565);
  nand n17567(x17567, x17436, x17416);
  nand n17569(x17569, x17441, x17419);
  nand n17571(x17571, x17569, x17570);
  nand n17572(x17572, x17441, x17421);
  nand n17574(x17574, x17446, x17424);
  nand n17576(x17576, x17574, x17575);
  nand n17577(x17577, x17446, x17426);
  nand n17579(x17579, x17451, x17429);
  nand n17581(x17581, x17579, x17580);
  nand n17582(x17582, x17451, x17431);
  nand n17584(x17584, x17456, x17434);
  nand n17586(x17586, x17584, x17585);
  nand n17587(x17587, x17456, x17436);
  nand n17589(x17589, x17461, x17439);
  nand n17591(x17591, x17589, x17590);
  nand n17592(x17592, x17461, x17441);
  nand n17594(x17594, x17478, x71977);
  nand n17596(x17596, x17594, x17595);
  nand n17597(x17597, x17483, x17195);
  nand n17599(x17599, x17597, x17598);
  nand n17600(x17600, x17488, x17318);
  nand n17602(x17602, x17600, x17601);
  nand n17603(x17603, x17493, x17321);
  nand n17605(x17605, x17603, x17604);
  nand n17606(x17606, x17498, x17464);
  nand n17608(x17608, x17606, x17607);
  nand n17609(x17609, x17503, x17467);
  nand n17611(x17611, x17609, x17610);
  nand n17612(x17612, x17508, x17470);
  nand n17614(x17614, x17612, x17613);
  nand n17615(x17615, x17513, x17473);
  nand n17617(x17617, x17615, x17616);
  nand n17618(x17618, x17518, x17476);
  nand n17620(x17620, x17618, x17619);
  nand n17621(x17621, x17518, x17478);
  nand n17623(x17623, x17523, x17481);
  nand n17625(x17625, x17623, x17624);
  nand n17626(x17626, x17523, x17483);
  nand n17628(x17628, x17528, x17486);
  nand n17630(x17630, x17628, x17629);
  nand n17631(x17631, x17528, x17488);
  nand n17633(x17633, x17533, x17491);
  nand n17635(x17635, x17633, x17634);
  nand n17636(x17636, x17533, x17493);
  nand n17638(x17638, x17538, x17496);
  nand n17640(x17640, x17638, x17639);
  nand n17641(x17641, x17538, x17498);
  nand n17643(x17643, x17543, x17501);
  nand n17645(x17645, x17643, x17644);
  nand n17646(x17646, x17543, x17503);
  nand n17648(x17648, x17548, x17506);
  nand n17650(x17650, x17648, x17649);
  nand n17651(x17651, x17548, x17508);
  nand n17653(x17653, x17553, x17511);
  nand n17655(x17655, x17653, x17654);
  nand n17656(x17656, x17553, x17513);
  nand n17658(x17658, x17558, x17516);
  nand n17660(x17660, x17658, x17659);
  nand n17661(x17661, x17558, x17518);
  nand n17663(x17663, x17563, x17521);
  nand n17665(x17665, x17663, x17664);
  nand n17666(x17666, x17563, x17523);
  nand n17668(x17668, x17568, x17526);
  nand n17670(x17670, x17668, x17669);
  nand n17671(x17671, x17568, x17528);
  nand n17673(x17673, x17573, x17531);
  nand n17675(x17675, x17673, x17674);
  nand n17676(x17676, x17573, x17533);
  nand n17678(x17678, x17578, x17536);
  nand n17680(x17680, x17678, x17679);
  nand n17681(x17681, x17578, x17538);
  nand n17683(x17683, x17583, x17541);
  nand n17685(x17685, x17683, x17684);
  nand n17686(x17686, x17583, x17543);
  nand n17688(x17688, x17588, x17546);
  nand n17690(x17690, x17688, x17689);
  nand n17691(x17691, x17588, x17548);
  nand n17693(x17693, x17593, x17551);
  nand n17695(x17695, x17693, x17694);
  nand n17696(x17696, x17593, x17553);
  nand n17698(x17698, x17622, x71977);
  nand n17700(x17700, x17698, x17699);
  nand n17701(x17701, x17627, x17195);
  nand n17703(x17703, x17701, x17702);
  nand n17704(x17704, x17632, x17318);
  nand n17706(x17706, x17704, x17705);
  nand n17707(x17707, x17637, x17321);
  nand n17709(x17709, x17707, x17708);
  nand n17710(x17710, x17642, x17464);
  nand n17712(x17712, x17710, x17711);
  nand n17713(x17713, x17647, x17467);
  nand n17715(x17715, x17713, x17714);
  nand n17716(x17716, x17652, x17470);
  nand n17718(x17718, x17716, x17717);
  nand n17719(x17719, x17657, x17473);
  nand n17721(x17721, x17719, x17720);
  nand n17722(x17722, x17662, x17596);
  nand n17724(x17724, x17722, x17723);
  nand n17725(x17725, x17667, x17599);
  nand n17727(x17727, x17725, x17726);
  nand n17728(x17728, x17672, x17602);
  nand n17730(x17730, x17728, x17729);
  nand n17731(x17731, x17677, x17605);
  nand n17733(x17733, x17731, x17732);
  nand n17734(x17734, x17682, x17608);
  nand n17736(x17736, x17734, x17735);
  nand n17737(x17737, x17687, x17611);
  nand n17739(x17739, x17737, x17738);
  nand n17740(x17740, x17692, x17614);
  nand n17742(x17742, x17740, x17741);
  nand n17743(x17743, x17697, x17617);
  nand n17745(x17745, x17743, x17744);
  nand n17746(x17746, x16976, x16876);
  nand n17747(x17747, x17746, x17194);
  nand n17749(x17749, x16983, x17195);
  nand n17751(x17751, x16982, x17750);
  nand n17752(x17752, x17751, x17749);
  nand n17754(x17754, x16989, x17318);
  nand n17756(x17756, x16988, x17755);
  nand n17757(x17757, x17756, x17754);
  nand n17759(x17759, x16995, x17321);
  nand n17761(x17761, x16994, x17760);
  nand n17762(x17762, x17761, x17759);
  nand n17764(x17764, x17001, x17464);
  nand n17766(x17766, x17000, x17765);
  nand n17767(x17767, x17766, x17764);
  nand n17769(x17769, x17007, x17467);
  nand n17771(x17771, x17006, x17770);
  nand n17772(x17772, x17771, x17769);
  nand n17774(x17774, x17013, x17470);
  nand n17776(x17776, x17012, x17775);
  nand n17777(x17777, x17776, x17774);
  nand n17779(x17779, x17019, x17473);
  nand n17781(x17781, x17018, x17780);
  nand n17782(x17782, x17781, x17779);
  nand n17784(x17784, x17025, x17596);
  nand n17786(x17786, x17024, x17785);
  nand n17787(x17787, x17786, x17784);
  nand n17789(x17789, x17031, x17599);
  nand n17791(x17791, x17030, x17790);
  nand n17792(x17792, x17791, x17789);
  nand n17794(x17794, x17037, x17602);
  nand n17796(x17796, x17036, x17795);
  nand n17797(x17797, x17796, x17794);
  nand n17799(x17799, x17043, x17605);
  nand n17801(x17801, x17042, x17800);
  nand n17802(x17802, x17801, x17799);
  nand n17804(x17804, x17049, x17608);
  nand n17806(x17806, x17048, x17805);
  nand n17807(x17807, x17806, x17804);
  nand n17809(x17809, x17055, x17611);
  nand n17811(x17811, x17054, x17810);
  nand n17812(x17812, x17811, x17809);
  nand n17814(x17814, x17061, x17614);
  nand n17816(x17816, x17060, x17815);
  nand n17817(x17817, x17816, x17814);
  nand n17819(x17819, x17067, x17617);
  nand n17821(x17821, x17066, x17820);
  nand n17822(x17822, x17821, x17819);
  nand n17824(x17824, x17073, x17700);
  nand n17826(x17826, x17072, x17825);
  nand n17827(x17827, x17826, x17824);
  nand n17829(x17829, x17079, x17703);
  nand n17831(x17831, x17078, x17830);
  nand n17832(x17832, x17831, x17829);
  nand n17834(x17834, x17085, x17706);
  nand n17836(x17836, x17084, x17835);
  nand n17837(x17837, x17836, x17834);
  nand n17839(x17839, x17091, x17709);
  nand n17841(x17841, x17090, x17840);
  nand n17842(x17842, x17841, x17839);
  nand n17844(x17844, x17097, x17712);
  nand n17846(x17846, x17096, x17845);
  nand n17847(x17847, x17846, x17844);
  nand n17849(x17849, x17103, x17715);
  nand n17851(x17851, x17102, x17850);
  nand n17852(x17852, x17851, x17849);
  nand n17854(x17854, x17109, x17718);
  nand n17856(x17856, x17108, x17855);
  nand n17857(x17857, x17856, x17854);
  nand n17859(x17859, x17115, x17721);
  nand n17861(x17861, x17114, x17860);
  nand n17862(x17862, x17861, x17859);
  nand n17864(x17864, x17121, x17724);
  nand n17866(x17866, x17120, x17865);
  nand n17867(x17867, x17866, x17864);
  nand n17869(x17869, x17127, x17727);
  nand n17871(x17871, x17126, x17870);
  nand n17872(x17872, x17871, x17869);
  nand n17874(x17874, x17133, x17730);
  nand n17876(x17876, x17132, x17875);
  nand n17877(x17877, x17876, x17874);
  nand n17879(x17879, x17139, x17733);
  nand n17881(x17881, x17138, x17880);
  nand n17882(x17882, x17881, x17879);
  nand n17884(x17884, x17145, x17736);
  nand n17886(x17886, x17144, x17885);
  nand n17887(x17887, x17886, x17884);
  nand n17889(x17889, x17151, x17739);
  nand n17891(x17891, x17150, x17890);
  nand n17892(x17892, x17891, x17889);
  nand n17894(x17894, x17157, x17742);
  nand n17896(x17896, x17156, x17895);
  nand n17897(x17897, x17896, x17894);
  nand n17899(x17899, x17163, x17745);
  nand n17901(x17901, x17162, x17900);
  nand n17902(x17902, x17901, x17899);
  nand n17904(x17904, x72047, x16749);
  nand n17905(x17905, x72052, x16749);
  nand n17907(x17907, x72047, x16752);
  nand n17909(x17909, x72057, x16749);
  nand n17911(x17911, x72052, x16752);
  nand n17913(x17913, x72047, x16755);
  nand n17915(x17915, x72062, x16749);
  nand n17917(x17917, x72057, x16752);
  nand n17919(x17919, x72052, x16755);
  nand n17921(x17921, x72047, x16758);
  nand n17922(x17922, x72067, x16749);
  nand n17924(x17924, x72062, x16752);
  nand n17926(x17926, x72057, x16755);
  nand n17928(x17928, x72052, x16758);
  nand n17930(x17930, x72047, x16761);
  nand n17932(x17932, x72072, x16749);
  nand n17934(x17934, x72067, x16752);
  nand n17936(x17936, x72062, x16755);
  nand n17938(x17938, x72057, x16758);
  nand n17940(x17940, x72052, x16761);
  nand n17942(x17942, x72047, x16764);
  nand n17944(x17944, x72077, x16749);
  nand n17946(x17946, x72072, x16752);
  nand n17948(x17948, x72067, x16755);
  nand n17950(x17950, x72062, x16758);
  nand n17952(x17952, x72057, x16761);
  nand n17954(x17954, x72052, x16764);
  nand n17956(x17956, x72047, x16767);
  nand n17957(x17957, x72082, x16749);
  nand n17959(x17959, x72077, x16752);
  nand n17961(x17961, x72072, x16755);
  nand n17963(x17963, x72067, x16758);
  nand n17965(x17965, x72062, x16761);
  nand n17967(x17967, x72057, x16764);
  nand n17969(x17969, x72052, x16767);
  nand n17971(x17971, x72047, x16770);
  nand n17973(x17973, x72087, x16749);
  nand n17975(x17975, x72082, x16752);
  nand n17977(x17977, x72077, x16755);
  nand n17979(x17979, x72072, x16758);
  nand n17981(x17981, x72067, x16761);
  nand n17983(x17983, x72062, x16764);
  nand n17985(x17985, x72057, x16767);
  nand n17987(x17987, x72052, x16770);
  nand n17989(x17989, x72047, x16773);
  nand n17991(x17991, x72092, x16749);
  nand n17993(x17993, x72087, x16752);
  nand n17995(x17995, x72082, x16755);
  nand n17997(x17997, x72077, x16758);
  nand n17999(x17999, x72072, x16761);
  nand n18001(x18001, x72067, x16764);
  nand n18003(x18003, x72062, x16767);
  nand n18005(x18005, x72057, x16770);
  nand n18007(x18007, x72052, x16773);
  nand n18009(x18009, x72047, x16776);
  nand n18010(x18010, x72097, x16749);
  nand n18012(x18012, x72092, x16752);
  nand n18014(x18014, x72087, x16755);
  nand n18016(x18016, x72082, x16758);
  nand n18018(x18018, x72077, x16761);
  nand n18020(x18020, x72072, x16764);
  nand n18022(x18022, x72067, x16767);
  nand n18024(x18024, x72062, x16770);
  nand n18026(x18026, x72057, x16773);
  nand n18028(x18028, x72052, x16776);
  nand n18030(x18030, x72047, x16779);
  nand n18032(x18032, x72102, x16749);
  nand n18034(x18034, x72097, x16752);
  nand n18036(x18036, x72092, x16755);
  nand n18038(x18038, x72087, x16758);
  nand n18040(x18040, x72082, x16761);
  nand n18042(x18042, x72077, x16764);
  nand n18044(x18044, x72072, x16767);
  nand n18046(x18046, x72067, x16770);
  nand n18048(x18048, x72062, x16773);
  nand n18050(x18050, x72057, x16776);
  nand n18052(x18052, x72052, x16779);
  nand n18054(x18054, x72047, x16782);
  nand n18056(x18056, x72107, x16749);
  nand n18058(x18058, x72102, x16752);
  nand n18060(x18060, x72097, x16755);
  nand n18062(x18062, x72092, x16758);
  nand n18064(x18064, x72087, x16761);
  nand n18066(x18066, x72082, x16764);
  nand n18068(x18068, x72077, x16767);
  nand n18070(x18070, x72072, x16770);
  nand n18072(x18072, x72067, x16773);
  nand n18074(x18074, x72062, x16776);
  nand n18076(x18076, x72057, x16779);
  nand n18078(x18078, x72052, x16782);
  nand n18080(x18080, x72047, x16785);
  nand n18081(x18081, x72112, x16749);
  nand n18083(x18083, x72107, x16752);
  nand n18085(x18085, x72102, x16755);
  nand n18087(x18087, x72097, x16758);
  nand n18089(x18089, x72092, x16761);
  nand n18091(x18091, x72087, x16764);
  nand n18093(x18093, x72082, x16767);
  nand n18095(x18095, x72077, x16770);
  nand n18097(x18097, x72072, x16773);
  nand n18099(x18099, x72067, x16776);
  nand n18101(x18101, x72062, x16779);
  nand n18103(x18103, x72057, x16782);
  nand n18105(x18105, x72052, x16785);
  nand n18107(x18107, x72047, x16788);
  nand n18109(x18109, x72117, x16749);
  nand n18111(x18111, x72112, x16752);
  nand n18113(x18113, x72107, x16755);
  nand n18115(x18115, x72102, x16758);
  nand n18117(x18117, x72097, x16761);
  nand n18119(x18119, x72092, x16764);
  nand n18121(x18121, x72087, x16767);
  nand n18123(x18123, x72082, x16770);
  nand n18125(x18125, x72077, x16773);
  nand n18127(x18127, x72072, x16776);
  nand n18129(x18129, x72067, x16779);
  nand n18131(x18131, x72062, x16782);
  nand n18133(x18133, x72057, x16785);
  nand n18135(x18135, x72052, x16788);
  nand n18137(x18137, x72047, x16791);
  nand n18139(x18139, x72122, x16749);
  nand n18141(x18141, x72117, x16752);
  nand n18143(x18143, x72112, x16755);
  nand n18145(x18145, x72107, x16758);
  nand n18147(x18147, x72102, x16761);
  nand n18149(x18149, x72097, x16764);
  nand n18151(x18151, x72092, x16767);
  nand n18153(x18153, x72087, x16770);
  nand n18155(x18155, x72082, x16773);
  nand n18157(x18157, x72077, x16776);
  nand n18159(x18159, x72072, x16779);
  nand n18161(x18161, x72067, x16782);
  nand n18163(x18163, x72062, x16785);
  nand n18165(x18165, x72057, x16788);
  nand n18167(x18167, x72052, x16791);
  nand n18169(x18169, x72047, x16794);
  nand n18170(x18170, x72127, x16749);
  nand n18172(x18172, x72122, x16752);
  nand n18174(x18174, x72117, x16755);
  nand n18176(x18176, x72112, x16758);
  nand n18178(x18178, x72107, x16761);
  nand n18180(x18180, x72102, x16764);
  nand n18182(x18182, x72097, x16767);
  nand n18184(x18184, x72092, x16770);
  nand n18186(x18186, x72087, x16773);
  nand n18188(x18188, x72082, x16776);
  nand n18190(x18190, x72077, x16779);
  nand n18192(x18192, x72072, x16782);
  nand n18194(x18194, x72067, x16785);
  nand n18196(x18196, x72062, x16788);
  nand n18198(x18198, x72057, x16791);
  nand n18200(x18200, x72052, x16794);
  nand n18202(x18202, x72047, x16797);
  nand n18204(x18204, x72132, x16749);
  nand n18206(x18206, x72127, x16752);
  nand n18208(x18208, x72122, x16755);
  nand n18210(x18210, x72117, x16758);
  nand n18212(x18212, x72112, x16761);
  nand n18214(x18214, x72107, x16764);
  nand n18216(x18216, x72102, x16767);
  nand n18218(x18218, x72097, x16770);
  nand n18220(x18220, x72092, x16773);
  nand n18222(x18222, x72087, x16776);
  nand n18224(x18224, x72082, x16779);
  nand n18226(x18226, x72077, x16782);
  nand n18228(x18228, x72072, x16785);
  nand n18230(x18230, x72067, x16788);
  nand n18232(x18232, x72062, x16791);
  nand n18234(x18234, x72057, x16794);
  nand n18236(x18236, x72052, x16797);
  nand n18238(x18238, x72047, x16800);
  nand n18240(x18240, x72137, x16749);
  nand n18242(x18242, x72132, x16752);
  nand n18244(x18244, x72127, x16755);
  nand n18246(x18246, x72122, x16758);
  nand n18248(x18248, x72117, x16761);
  nand n18250(x18250, x72112, x16764);
  nand n18252(x18252, x72107, x16767);
  nand n18254(x18254, x72102, x16770);
  nand n18256(x18256, x72097, x16773);
  nand n18258(x18258, x72092, x16776);
  nand n18260(x18260, x72087, x16779);
  nand n18262(x18262, x72082, x16782);
  nand n18264(x18264, x72077, x16785);
  nand n18266(x18266, x72072, x16788);
  nand n18268(x18268, x72067, x16791);
  nand n18270(x18270, x72062, x16794);
  nand n18272(x18272, x72057, x16797);
  nand n18274(x18274, x72052, x16800);
  nand n18276(x18276, x72047, x16803);
  nand n18277(x18277, x72142, x16749);
  nand n18279(x18279, x72137, x16752);
  nand n18281(x18281, x72132, x16755);
  nand n18283(x18283, x72127, x16758);
  nand n18285(x18285, x72122, x16761);
  nand n18287(x18287, x72117, x16764);
  nand n18289(x18289, x72112, x16767);
  nand n18291(x18291, x72107, x16770);
  nand n18293(x18293, x72102, x16773);
  nand n18295(x18295, x72097, x16776);
  nand n18297(x18297, x72092, x16779);
  nand n18299(x18299, x72087, x16782);
  nand n18301(x18301, x72082, x16785);
  nand n18303(x18303, x72077, x16788);
  nand n18305(x18305, x72072, x16791);
  nand n18307(x18307, x72067, x16794);
  nand n18309(x18309, x72062, x16797);
  nand n18311(x18311, x72057, x16800);
  nand n18313(x18313, x72052, x16803);
  nand n18315(x18315, x72047, x16806);
  nand n18317(x18317, x72147, x16749);
  nand n18319(x18319, x72142, x16752);
  nand n18321(x18321, x72137, x16755);
  nand n18323(x18323, x72132, x16758);
  nand n18325(x18325, x72127, x16761);
  nand n18327(x18327, x72122, x16764);
  nand n18329(x18329, x72117, x16767);
  nand n18331(x18331, x72112, x16770);
  nand n18333(x18333, x72107, x16773);
  nand n18335(x18335, x72102, x16776);
  nand n18337(x18337, x72097, x16779);
  nand n18339(x18339, x72092, x16782);
  nand n18341(x18341, x72087, x16785);
  nand n18343(x18343, x72082, x16788);
  nand n18345(x18345, x72077, x16791);
  nand n18347(x18347, x72072, x16794);
  nand n18349(x18349, x72067, x16797);
  nand n18351(x18351, x72062, x16800);
  nand n18353(x18353, x72057, x16803);
  nand n18355(x18355, x72052, x16806);
  nand n18357(x18357, x72047, x16809);
  nand n18359(x18359, x72152, x16749);
  nand n18361(x18361, x72147, x16752);
  nand n18363(x18363, x72142, x16755);
  nand n18365(x18365, x72137, x16758);
  nand n18367(x18367, x72132, x16761);
  nand n18369(x18369, x72127, x16764);
  nand n18371(x18371, x72122, x16767);
  nand n18373(x18373, x72117, x16770);
  nand n18375(x18375, x72112, x16773);
  nand n18377(x18377, x72107, x16776);
  nand n18379(x18379, x72102, x16779);
  nand n18381(x18381, x72097, x16782);
  nand n18383(x18383, x72092, x16785);
  nand n18385(x18385, x72087, x16788);
  nand n18387(x18387, x72082, x16791);
  nand n18389(x18389, x72077, x16794);
  nand n18391(x18391, x72072, x16797);
  nand n18393(x18393, x72067, x16800);
  nand n18395(x18395, x72062, x16803);
  nand n18397(x18397, x72057, x16806);
  nand n18399(x18399, x72052, x16809);
  nand n18401(x18401, x72047, x16812);
  nand n18402(x18402, x72157, x16749);
  nand n18404(x18404, x72152, x16752);
  nand n18406(x18406, x72147, x16755);
  nand n18408(x18408, x72142, x16758);
  nand n18410(x18410, x72137, x16761);
  nand n18412(x18412, x72132, x16764);
  nand n18414(x18414, x72127, x16767);
  nand n18416(x18416, x72122, x16770);
  nand n18418(x18418, x72117, x16773);
  nand n18420(x18420, x72112, x16776);
  nand n18422(x18422, x72107, x16779);
  nand n18424(x18424, x72102, x16782);
  nand n18426(x18426, x72097, x16785);
  nand n18428(x18428, x72092, x16788);
  nand n18430(x18430, x72087, x16791);
  nand n18432(x18432, x72082, x16794);
  nand n18434(x18434, x72077, x16797);
  nand n18436(x18436, x72072, x16800);
  nand n18438(x18438, x72067, x16803);
  nand n18440(x18440, x72062, x16806);
  nand n18442(x18442, x72057, x16809);
  nand n18444(x18444, x72052, x16812);
  nand n18446(x18446, x72047, x16815);
  nand n18448(x18448, x72162, x16749);
  nand n18450(x18450, x72157, x16752);
  nand n18452(x18452, x72152, x16755);
  nand n18454(x18454, x72147, x16758);
  nand n18456(x18456, x72142, x16761);
  nand n18458(x18458, x72137, x16764);
  nand n18460(x18460, x72132, x16767);
  nand n18462(x18462, x72127, x16770);
  nand n18464(x18464, x72122, x16773);
  nand n18466(x18466, x72117, x16776);
  nand n18468(x18468, x72112, x16779);
  nand n18470(x18470, x72107, x16782);
  nand n18472(x18472, x72102, x16785);
  nand n18474(x18474, x72097, x16788);
  nand n18476(x18476, x72092, x16791);
  nand n18478(x18478, x72087, x16794);
  nand n18480(x18480, x72082, x16797);
  nand n18482(x18482, x72077, x16800);
  nand n18484(x18484, x72072, x16803);
  nand n18486(x18486, x72067, x16806);
  nand n18488(x18488, x72062, x16809);
  nand n18490(x18490, x72057, x16812);
  nand n18492(x18492, x72052, x16815);
  nand n18494(x18494, x72047, x16818);
  nand n18496(x18496, x72167, x16749);
  nand n18498(x18498, x72162, x16752);
  nand n18500(x18500, x72157, x16755);
  nand n18502(x18502, x72152, x16758);
  nand n18504(x18504, x72147, x16761);
  nand n18506(x18506, x72142, x16764);
  nand n18508(x18508, x72137, x16767);
  nand n18510(x18510, x72132, x16770);
  nand n18512(x18512, x72127, x16773);
  nand n18514(x18514, x72122, x16776);
  nand n18516(x18516, x72117, x16779);
  nand n18518(x18518, x72112, x16782);
  nand n18520(x18520, x72107, x16785);
  nand n18522(x18522, x72102, x16788);
  nand n18524(x18524, x72097, x16791);
  nand n18526(x18526, x72092, x16794);
  nand n18528(x18528, x72087, x16797);
  nand n18530(x18530, x72082, x16800);
  nand n18532(x18532, x72077, x16803);
  nand n18534(x18534, x72072, x16806);
  nand n18536(x18536, x72067, x16809);
  nand n18538(x18538, x72062, x16812);
  nand n18540(x18540, x72057, x16815);
  nand n18542(x18542, x72052, x16818);
  nand n18544(x18544, x72047, x16821);
  nand n18545(x18545, x72172, x16749);
  nand n18547(x18547, x72167, x16752);
  nand n18549(x18549, x72162, x16755);
  nand n18551(x18551, x72157, x16758);
  nand n18553(x18553, x72152, x16761);
  nand n18555(x18555, x72147, x16764);
  nand n18557(x18557, x72142, x16767);
  nand n18559(x18559, x72137, x16770);
  nand n18561(x18561, x72132, x16773);
  nand n18563(x18563, x72127, x16776);
  nand n18565(x18565, x72122, x16779);
  nand n18567(x18567, x72117, x16782);
  nand n18569(x18569, x72112, x16785);
  nand n18571(x18571, x72107, x16788);
  nand n18573(x18573, x72102, x16791);
  nand n18575(x18575, x72097, x16794);
  nand n18577(x18577, x72092, x16797);
  nand n18579(x18579, x72087, x16800);
  nand n18581(x18581, x72082, x16803);
  nand n18583(x18583, x72077, x16806);
  nand n18585(x18585, x72072, x16809);
  nand n18587(x18587, x72067, x16812);
  nand n18589(x18589, x72062, x16815);
  nand n18591(x18591, x72057, x16818);
  nand n18593(x18593, x72052, x16821);
  nand n18595(x18595, x72047, x16824);
  nand n18597(x18597, x72177, x16749);
  nand n18599(x18599, x72172, x16752);
  nand n18601(x18601, x72167, x16755);
  nand n18603(x18603, x72162, x16758);
  nand n18605(x18605, x72157, x16761);
  nand n18607(x18607, x72152, x16764);
  nand n18609(x18609, x72147, x16767);
  nand n18611(x18611, x72142, x16770);
  nand n18613(x18613, x72137, x16773);
  nand n18615(x18615, x72132, x16776);
  nand n18617(x18617, x72127, x16779);
  nand n18619(x18619, x72122, x16782);
  nand n18621(x18621, x72117, x16785);
  nand n18623(x18623, x72112, x16788);
  nand n18625(x18625, x72107, x16791);
  nand n18627(x18627, x72102, x16794);
  nand n18629(x18629, x72097, x16797);
  nand n18631(x18631, x72092, x16800);
  nand n18633(x18633, x72087, x16803);
  nand n18635(x18635, x72082, x16806);
  nand n18637(x18637, x72077, x16809);
  nand n18639(x18639, x72072, x16812);
  nand n18641(x18641, x72067, x16815);
  nand n18643(x18643, x72062, x16818);
  nand n18645(x18645, x72057, x16821);
  nand n18647(x18647, x72052, x16824);
  nand n18649(x18649, x72047, x16827);
  nand n18651(x18651, x72182, x16749);
  nand n18653(x18653, x72177, x16752);
  nand n18655(x18655, x72172, x16755);
  nand n18657(x18657, x72167, x16758);
  nand n18659(x18659, x72162, x16761);
  nand n18661(x18661, x72157, x16764);
  nand n18663(x18663, x72152, x16767);
  nand n18665(x18665, x72147, x16770);
  nand n18667(x18667, x72142, x16773);
  nand n18669(x18669, x72137, x16776);
  nand n18671(x18671, x72132, x16779);
  nand n18673(x18673, x72127, x16782);
  nand n18675(x18675, x72122, x16785);
  nand n18677(x18677, x72117, x16788);
  nand n18679(x18679, x72112, x16791);
  nand n18681(x18681, x72107, x16794);
  nand n18683(x18683, x72102, x16797);
  nand n18685(x18685, x72097, x16800);
  nand n18687(x18687, x72092, x16803);
  nand n18689(x18689, x72087, x16806);
  nand n18691(x18691, x72082, x16809);
  nand n18693(x18693, x72077, x16812);
  nand n18695(x18695, x72072, x16815);
  nand n18697(x18697, x72067, x16818);
  nand n18699(x18699, x72062, x16821);
  nand n18701(x18701, x72057, x16824);
  nand n18703(x18703, x72052, x16827);
  nand n18705(x18705, x72047, x16830);
  nand n18706(x18706, x72187, x16749);
  nand n18708(x18708, x72182, x16752);
  nand n18710(x18710, x72177, x16755);
  nand n18712(x18712, x72172, x16758);
  nand n18714(x18714, x72167, x16761);
  nand n18716(x18716, x72162, x16764);
  nand n18718(x18718, x72157, x16767);
  nand n18720(x18720, x72152, x16770);
  nand n18722(x18722, x72147, x16773);
  nand n18724(x18724, x72142, x16776);
  nand n18726(x18726, x72137, x16779);
  nand n18728(x18728, x72132, x16782);
  nand n18730(x18730, x72127, x16785);
  nand n18732(x18732, x72122, x16788);
  nand n18734(x18734, x72117, x16791);
  nand n18736(x18736, x72112, x16794);
  nand n18738(x18738, x72107, x16797);
  nand n18740(x18740, x72102, x16800);
  nand n18742(x18742, x72097, x16803);
  nand n18744(x18744, x72092, x16806);
  nand n18746(x18746, x72087, x16809);
  nand n18748(x18748, x72082, x16812);
  nand n18750(x18750, x72077, x16815);
  nand n18752(x18752, x72072, x16818);
  nand n18754(x18754, x72067, x16821);
  nand n18756(x18756, x72062, x16824);
  nand n18758(x18758, x72057, x16827);
  nand n18760(x18760, x72052, x16830);
  nand n18762(x18762, x72047, x16833);
  nand n18764(x18764, x72192, x16749);
  nand n18766(x18766, x72187, x16752);
  nand n18768(x18768, x72182, x16755);
  nand n18770(x18770, x72177, x16758);
  nand n18772(x18772, x72172, x16761);
  nand n18774(x18774, x72167, x16764);
  nand n18776(x18776, x72162, x16767);
  nand n18778(x18778, x72157, x16770);
  nand n18780(x18780, x72152, x16773);
  nand n18782(x18782, x72147, x16776);
  nand n18784(x18784, x72142, x16779);
  nand n18786(x18786, x72137, x16782);
  nand n18788(x18788, x72132, x16785);
  nand n18790(x18790, x72127, x16788);
  nand n18792(x18792, x72122, x16791);
  nand n18794(x18794, x72117, x16794);
  nand n18796(x18796, x72112, x16797);
  nand n18798(x18798, x72107, x16800);
  nand n18800(x18800, x72102, x16803);
  nand n18802(x18802, x72097, x16806);
  nand n18804(x18804, x72092, x16809);
  nand n18806(x18806, x72087, x16812);
  nand n18808(x18808, x72082, x16815);
  nand n18810(x18810, x72077, x16818);
  nand n18812(x18812, x72072, x16821);
  nand n18814(x18814, x72067, x16824);
  nand n18816(x18816, x72062, x16827);
  nand n18818(x18818, x72057, x16830);
  nand n18820(x18820, x72052, x16833);
  nand n18822(x18822, x72047, x16836);
  nand n18824(x18824, x72197, x16749);
  nand n18826(x18826, x72192, x16752);
  nand n18828(x18828, x72187, x16755);
  nand n18830(x18830, x72182, x16758);
  nand n18832(x18832, x72177, x16761);
  nand n18834(x18834, x72172, x16764);
  nand n18836(x18836, x72167, x16767);
  nand n18838(x18838, x72162, x16770);
  nand n18840(x18840, x72157, x16773);
  nand n18842(x18842, x72152, x16776);
  nand n18844(x18844, x72147, x16779);
  nand n18846(x18846, x72142, x16782);
  nand n18848(x18848, x72137, x16785);
  nand n18850(x18850, x72132, x16788);
  nand n18852(x18852, x72127, x16791);
  nand n18854(x18854, x72122, x16794);
  nand n18856(x18856, x72117, x16797);
  nand n18858(x18858, x72112, x16800);
  nand n18860(x18860, x72107, x16803);
  nand n18862(x18862, x72102, x16806);
  nand n18864(x18864, x72097, x16809);
  nand n18866(x18866, x72092, x16812);
  nand n18868(x18868, x72087, x16815);
  nand n18870(x18870, x72082, x16818);
  nand n18872(x18872, x72077, x16821);
  nand n18874(x18874, x72072, x16824);
  nand n18876(x18876, x72067, x16827);
  nand n18878(x18878, x72062, x16830);
  nand n18880(x18880, x72057, x16833);
  nand n18882(x18882, x72052, x16836);
  nand n18884(x18884, x72047, x16839);
  nand n18885(x18885, x72202, x16749);
  nand n18887(x18887, x72197, x16752);
  nand n18889(x18889, x72192, x16755);
  nand n18891(x18891, x72187, x16758);
  nand n18893(x18893, x72182, x16761);
  nand n18895(x18895, x72177, x16764);
  nand n18897(x18897, x72172, x16767);
  nand n18899(x18899, x72167, x16770);
  nand n18901(x18901, x72162, x16773);
  nand n18903(x18903, x72157, x16776);
  nand n18905(x18905, x72152, x16779);
  nand n18907(x18907, x72147, x16782);
  nand n18909(x18909, x72142, x16785);
  nand n18911(x18911, x72137, x16788);
  nand n18913(x18913, x72132, x16791);
  nand n18915(x18915, x72127, x16794);
  nand n18917(x18917, x72122, x16797);
  nand n18919(x18919, x72117, x16800);
  nand n18921(x18921, x72112, x16803);
  nand n18923(x18923, x72107, x16806);
  nand n18925(x18925, x72102, x16809);
  nand n18927(x18927, x72097, x16812);
  nand n18929(x18929, x72092, x16815);
  nand n18931(x18931, x72087, x16818);
  nand n18933(x18933, x72082, x16821);
  nand n18935(x18935, x72077, x16824);
  nand n18937(x18937, x72072, x16827);
  nand n18939(x18939, x72067, x16830);
  nand n18941(x18941, x72062, x16833);
  nand n18943(x18943, x72057, x16836);
  nand n18945(x18945, x72052, x16839);
  nand n18947(x18947, x72047, x16842);
  nand n18949(x18949, x17906, x17908);
  nand n18950(x18950, x17905, x17907);
  nand n18951(x18951, x18950, x18949);
  nand n18952(x18952, x17910, x17912);
  nand n18953(x18953, x17909, x17911);
  nand n18954(x18954, x18953, x18952);
  nand n18956(x18956, x17914, x18955);
  nand n18957(x18957, x17913, x18954);
  nand n18958(x18958, x18957, x18956);
  nand n18959(x18959, x18952, x18956);
  nand n18960(x18960, x17916, x17918);
  nand n18961(x18961, x17915, x17917);
  nand n18962(x18962, x18961, x18960);
  nand n18964(x18964, x17920, x18963);
  nand n18965(x18965, x17919, x18962);
  nand n18966(x18966, x18965, x18964);
  nand n18967(x18967, x18960, x18964);
  nand n18968(x18968, x17923, x17925);
  nand n18969(x18969, x17922, x17924);
  nand n18970(x18970, x18969, x18968);
  nand n18972(x18972, x17927, x18971);
  nand n18973(x18973, x17926, x18970);
  nand n18974(x18974, x18973, x18972);
  nand n18975(x18975, x18968, x18972);
  nand n18976(x18976, x17929, x17931);
  nand n18977(x18977, x17928, x17930);
  nand n18978(x18978, x18977, x18976);
  nand n18979(x18979, x17933, x17935);
  nand n18980(x18980, x17932, x17934);
  nand n18981(x18981, x18980, x18979);
  nand n18983(x18983, x17937, x18982);
  nand n18984(x18984, x17936, x18981);
  nand n18985(x18985, x18984, x18983);
  nand n18986(x18986, x18979, x18983);
  nand n18987(x18987, x17939, x17941);
  nand n18988(x18988, x17938, x17940);
  nand n18989(x18989, x18988, x18987);
  nand n18991(x18991, x17943, x18990);
  nand n18992(x18992, x17942, x18989);
  nand n18993(x18993, x18992, x18991);
  nand n18994(x18994, x18987, x18991);
  nand n18995(x18995, x17945, x17947);
  nand n18996(x18996, x17944, x17946);
  nand n18997(x18997, x18996, x18995);
  nand n18999(x18999, x17949, x18998);
  nand n19000(x19000, x17948, x18997);
  nand n19001(x19001, x19000, x18999);
  nand n19002(x19002, x18995, x18999);
  nand n19003(x19003, x17951, x17953);
  nand n19004(x19004, x17950, x17952);
  nand n19005(x19005, x19004, x19003);
  nand n19007(x19007, x17955, x19006);
  nand n19008(x19008, x17954, x19005);
  nand n19009(x19009, x19008, x19007);
  nand n19011(x19011, x19003, x19007);
  nand n19012(x19012, x17958, x17960);
  nand n19013(x19013, x17957, x17959);
  nand n19014(x19014, x19013, x19012);
  nand n19016(x19016, x17962, x19015);
  nand n19017(x19017, x17961, x19014);
  nand n19018(x19018, x19017, x19016);
  nand n19019(x19019, x19012, x19016);
  nand n19020(x19020, x17964, x17966);
  nand n19021(x19021, x17963, x17965);
  nand n19022(x19022, x19021, x19020);
  nand n19024(x19024, x17968, x19023);
  nand n19025(x19025, x17967, x19022);
  nand n19026(x19026, x19025, x19024);
  nand n19028(x19028, x19020, x19024);
  nand n19029(x19029, x17970, x17972);
  nand n19030(x19030, x17969, x17971);
  nand n19031(x19031, x19030, x19029);
  nand n19032(x19032, x17974, x17976);
  nand n19033(x19033, x17973, x17975);
  nand n19034(x19034, x19033, x19032);
  nand n19036(x19036, x17978, x19035);
  nand n19037(x19037, x17977, x19034);
  nand n19038(x19038, x19037, x19036);
  nand n19039(x19039, x19032, x19036);
  nand n19040(x19040, x17980, x17982);
  nand n19041(x19041, x17979, x17981);
  nand n19042(x19042, x19041, x19040);
  nand n19044(x19044, x17984, x19043);
  nand n19045(x19045, x17983, x19042);
  nand n19046(x19046, x19045, x19044);
  nand n19048(x19048, x19040, x19044);
  nand n19049(x19049, x17986, x17988);
  nand n19050(x19050, x17985, x17987);
  nand n19051(x19051, x19050, x19049);
  nand n19053(x19053, x17990, x19052);
  nand n19054(x19054, x17989, x19051);
  nand n19055(x19055, x19054, x19053);
  nand n19057(x19057, x19049, x19053);
  nand n19058(x19058, x17992, x17994);
  nand n19059(x19059, x17991, x17993);
  nand n19060(x19060, x19059, x19058);
  nand n19062(x19062, x17996, x19061);
  nand n19063(x19063, x17995, x19060);
  nand n19064(x19064, x19063, x19062);
  nand n19065(x19065, x19058, x19062);
  nand n19066(x19066, x17998, x18000);
  nand n19067(x19067, x17997, x17999);
  nand n19068(x19068, x19067, x19066);
  nand n19070(x19070, x18002, x19069);
  nand n19071(x19071, x18001, x19068);
  nand n19072(x19072, x19071, x19070);
  nand n19074(x19074, x19066, x19070);
  nand n19075(x19075, x18004, x18006);
  nand n19076(x19076, x18003, x18005);
  nand n19077(x19077, x19076, x19075);
  nand n19079(x19079, x18008, x19078);
  nand n19080(x19080, x18007, x19077);
  nand n19081(x19081, x19080, x19079);
  nand n19083(x19083, x19075, x19079);
  nand n19084(x19084, x18011, x18013);
  nand n19085(x19085, x18010, x18012);
  nand n19086(x19086, x19085, x19084);
  nand n19088(x19088, x18015, x19087);
  nand n19089(x19089, x18014, x19086);
  nand n19090(x19090, x19089, x19088);
  nand n19091(x19091, x19084, x19088);
  nand n19092(x19092, x18017, x18019);
  nand n19093(x19093, x18016, x18018);
  nand n19094(x19094, x19093, x19092);
  nand n19096(x19096, x18021, x19095);
  nand n19097(x19097, x18020, x19094);
  nand n19098(x19098, x19097, x19096);
  nand n19100(x19100, x19092, x19096);
  nand n19101(x19101, x18023, x18025);
  nand n19102(x19102, x18022, x18024);
  nand n19103(x19103, x19102, x19101);
  nand n19105(x19105, x18027, x19104);
  nand n19106(x19106, x18026, x19103);
  nand n19107(x19107, x19106, x19105);
  nand n19109(x19109, x19101, x19105);
  nand n19110(x19110, x18029, x18031);
  nand n19111(x19111, x18028, x18030);
  nand n19112(x19112, x19111, x19110);
  nand n19113(x19113, x18033, x18035);
  nand n19114(x19114, x18032, x18034);
  nand n19115(x19115, x19114, x19113);
  nand n19117(x19117, x18037, x19116);
  nand n19118(x19118, x18036, x19115);
  nand n19119(x19119, x19118, x19117);
  nand n19120(x19120, x19113, x19117);
  nand n19121(x19121, x18039, x18041);
  nand n19122(x19122, x18038, x18040);
  nand n19123(x19123, x19122, x19121);
  nand n19125(x19125, x18043, x19124);
  nand n19126(x19126, x18042, x19123);
  nand n19127(x19127, x19126, x19125);
  nand n19129(x19129, x19121, x19125);
  nand n19130(x19130, x18045, x18047);
  nand n19131(x19131, x18044, x18046);
  nand n19132(x19132, x19131, x19130);
  nand n19134(x19134, x18049, x19133);
  nand n19135(x19135, x18048, x19132);
  nand n19136(x19136, x19135, x19134);
  nand n19138(x19138, x19130, x19134);
  nand n19139(x19139, x18051, x18053);
  nand n19140(x19140, x18050, x18052);
  nand n19141(x19141, x19140, x19139);
  nand n19143(x19143, x18055, x19142);
  nand n19144(x19144, x18054, x19141);
  nand n19145(x19145, x19144, x19143);
  nand n19147(x19147, x19139, x19143);
  nand n19148(x19148, x18057, x18059);
  nand n19149(x19149, x18056, x18058);
  nand n19150(x19150, x19149, x19148);
  nand n19152(x19152, x18061, x19151);
  nand n19153(x19153, x18060, x19150);
  nand n19154(x19154, x19153, x19152);
  nand n19155(x19155, x19148, x19152);
  nand n19156(x19156, x18063, x18065);
  nand n19157(x19157, x18062, x18064);
  nand n19158(x19158, x19157, x19156);
  nand n19160(x19160, x18067, x19159);
  nand n19161(x19161, x18066, x19158);
  nand n19162(x19162, x19161, x19160);
  nand n19164(x19164, x19156, x19160);
  nand n19165(x19165, x18069, x18071);
  nand n19166(x19166, x18068, x18070);
  nand n19167(x19167, x19166, x19165);
  nand n19169(x19169, x18073, x19168);
  nand n19170(x19170, x18072, x19167);
  nand n19171(x19171, x19170, x19169);
  nand n19173(x19173, x19165, x19169);
  nand n19174(x19174, x18075, x18077);
  nand n19175(x19175, x18074, x18076);
  nand n19176(x19176, x19175, x19174);
  nand n19178(x19178, x18079, x19177);
  nand n19179(x19179, x18078, x19176);
  nand n19180(x19180, x19179, x19178);
  nand n19182(x19182, x19174, x19178);
  nand n19183(x19183, x18082, x18084);
  nand n19184(x19184, x18081, x18083);
  nand n19185(x19185, x19184, x19183);
  nand n19187(x19187, x18086, x19186);
  nand n19188(x19188, x18085, x19185);
  nand n19189(x19189, x19188, x19187);
  nand n19190(x19190, x19183, x19187);
  nand n19191(x19191, x18088, x18090);
  nand n19192(x19192, x18087, x18089);
  nand n19193(x19193, x19192, x19191);
  nand n19195(x19195, x18092, x19194);
  nand n19196(x19196, x18091, x19193);
  nand n19197(x19197, x19196, x19195);
  nand n19199(x19199, x19191, x19195);
  nand n19200(x19200, x18094, x18096);
  nand n19201(x19201, x18093, x18095);
  nand n19202(x19202, x19201, x19200);
  nand n19204(x19204, x18098, x19203);
  nand n19205(x19205, x18097, x19202);
  nand n19206(x19206, x19205, x19204);
  nand n19208(x19208, x19200, x19204);
  nand n19209(x19209, x18100, x18102);
  nand n19210(x19210, x18099, x18101);
  nand n19211(x19211, x19210, x19209);
  nand n19213(x19213, x18104, x19212);
  nand n19214(x19214, x18103, x19211);
  nand n19215(x19215, x19214, x19213);
  nand n19217(x19217, x19209, x19213);
  nand n19218(x19218, x18106, x18108);
  nand n19219(x19219, x18105, x18107);
  nand n19220(x19220, x19219, x19218);
  nand n19221(x19221, x18110, x18112);
  nand n19222(x19222, x18109, x18111);
  nand n19223(x19223, x19222, x19221);
  nand n19225(x19225, x18114, x19224);
  nand n19226(x19226, x18113, x19223);
  nand n19227(x19227, x19226, x19225);
  nand n19228(x19228, x19221, x19225);
  nand n19229(x19229, x18116, x18118);
  nand n19230(x19230, x18115, x18117);
  nand n19231(x19231, x19230, x19229);
  nand n19233(x19233, x18120, x19232);
  nand n19234(x19234, x18119, x19231);
  nand n19235(x19235, x19234, x19233);
  nand n19237(x19237, x19229, x19233);
  nand n19238(x19238, x18122, x18124);
  nand n19239(x19239, x18121, x18123);
  nand n19240(x19240, x19239, x19238);
  nand n19242(x19242, x18126, x19241);
  nand n19243(x19243, x18125, x19240);
  nand n19244(x19244, x19243, x19242);
  nand n19246(x19246, x19238, x19242);
  nand n19247(x19247, x18128, x18130);
  nand n19248(x19248, x18127, x18129);
  nand n19249(x19249, x19248, x19247);
  nand n19251(x19251, x18132, x19250);
  nand n19252(x19252, x18131, x19249);
  nand n19253(x19253, x19252, x19251);
  nand n19255(x19255, x19247, x19251);
  nand n19256(x19256, x18134, x18136);
  nand n19257(x19257, x18133, x18135);
  nand n19258(x19258, x19257, x19256);
  nand n19260(x19260, x18138, x19259);
  nand n19261(x19261, x18137, x19258);
  nand n19262(x19262, x19261, x19260);
  nand n19263(x19263, x19256, x19260);
  nand n19264(x19264, x18140, x18142);
  nand n19265(x19265, x18139, x18141);
  nand n19266(x19266, x19265, x19264);
  nand n19268(x19268, x18144, x19267);
  nand n19269(x19269, x18143, x19266);
  nand n19270(x19270, x19269, x19268);
  nand n19271(x19271, x19264, x19268);
  nand n19272(x19272, x18146, x18148);
  nand n19273(x19273, x18145, x18147);
  nand n19274(x19274, x19273, x19272);
  nand n19276(x19276, x18150, x19275);
  nand n19277(x19277, x18149, x19274);
  nand n19278(x19278, x19277, x19276);
  nand n19280(x19280, x19272, x19276);
  nand n19281(x19281, x18152, x18154);
  nand n19282(x19282, x18151, x18153);
  nand n19283(x19283, x19282, x19281);
  nand n19285(x19285, x18156, x19284);
  nand n19286(x19286, x18155, x19283);
  nand n19287(x19287, x19286, x19285);
  nand n19289(x19289, x19281, x19285);
  nand n19290(x19290, x18158, x18160);
  nand n19291(x19291, x18157, x18159);
  nand n19292(x19292, x19291, x19290);
  nand n19294(x19294, x18162, x19293);
  nand n19295(x19295, x18161, x19292);
  nand n19296(x19296, x19295, x19294);
  nand n19298(x19298, x19290, x19294);
  nand n19299(x19299, x18164, x18166);
  nand n19300(x19300, x18163, x18165);
  nand n19301(x19301, x19300, x19299);
  nand n19303(x19303, x18168, x19302);
  nand n19304(x19304, x18167, x19301);
  nand n19305(x19305, x19304, x19303);
  nand n19307(x19307, x19299, x19303);
  nand n19308(x19308, x18171, x18173);
  nand n19309(x19309, x18170, x18172);
  nand n19310(x19310, x19309, x19308);
  nand n19312(x19312, x18175, x19311);
  nand n19313(x19313, x18174, x19310);
  nand n19314(x19314, x19313, x19312);
  nand n19315(x19315, x19308, x19312);
  nand n19316(x19316, x18177, x18179);
  nand n19317(x19317, x18176, x18178);
  nand n19318(x19318, x19317, x19316);
  nand n19320(x19320, x18181, x19319);
  nand n19321(x19321, x18180, x19318);
  nand n19322(x19322, x19321, x19320);
  nand n19324(x19324, x19316, x19320);
  nand n19325(x19325, x18183, x18185);
  nand n19326(x19326, x18182, x18184);
  nand n19327(x19327, x19326, x19325);
  nand n19329(x19329, x18187, x19328);
  nand n19330(x19330, x18186, x19327);
  nand n19331(x19331, x19330, x19329);
  nand n19333(x19333, x19325, x19329);
  nand n19334(x19334, x18189, x18191);
  nand n19335(x19335, x18188, x18190);
  nand n19336(x19336, x19335, x19334);
  nand n19338(x19338, x18193, x19337);
  nand n19339(x19339, x18192, x19336);
  nand n19340(x19340, x19339, x19338);
  nand n19342(x19342, x19334, x19338);
  nand n19343(x19343, x18195, x18197);
  nand n19344(x19344, x18194, x18196);
  nand n19345(x19345, x19344, x19343);
  nand n19347(x19347, x18199, x19346);
  nand n19348(x19348, x18198, x19345);
  nand n19349(x19349, x19348, x19347);
  nand n19351(x19351, x19343, x19347);
  nand n19352(x19352, x18201, x18203);
  nand n19353(x19353, x18200, x18202);
  nand n19354(x19354, x19353, x19352);
  nand n19355(x19355, x18205, x18207);
  nand n19356(x19356, x18204, x18206);
  nand n19357(x19357, x19356, x19355);
  nand n19359(x19359, x18209, x19358);
  nand n19360(x19360, x18208, x19357);
  nand n19361(x19361, x19360, x19359);
  nand n19362(x19362, x19355, x19359);
  nand n19363(x19363, x18211, x18213);
  nand n19364(x19364, x18210, x18212);
  nand n19365(x19365, x19364, x19363);
  nand n19367(x19367, x18215, x19366);
  nand n19368(x19368, x18214, x19365);
  nand n19369(x19369, x19368, x19367);
  nand n19371(x19371, x19363, x19367);
  nand n19372(x19372, x18217, x18219);
  nand n19373(x19373, x18216, x18218);
  nand n19374(x19374, x19373, x19372);
  nand n19376(x19376, x18221, x19375);
  nand n19377(x19377, x18220, x19374);
  nand n19378(x19378, x19377, x19376);
  nand n19380(x19380, x19372, x19376);
  nand n19381(x19381, x18223, x18225);
  nand n19382(x19382, x18222, x18224);
  nand n19383(x19383, x19382, x19381);
  nand n19385(x19385, x18227, x19384);
  nand n19386(x19386, x18226, x19383);
  nand n19387(x19387, x19386, x19385);
  nand n19389(x19389, x19381, x19385);
  nand n19390(x19390, x18229, x18231);
  nand n19391(x19391, x18228, x18230);
  nand n19392(x19392, x19391, x19390);
  nand n19394(x19394, x18233, x19393);
  nand n19395(x19395, x18232, x19392);
  nand n19396(x19396, x19395, x19394);
  nand n19398(x19398, x19390, x19394);
  nand n19399(x19399, x18235, x18237);
  nand n19400(x19400, x18234, x18236);
  nand n19401(x19401, x19400, x19399);
  nand n19403(x19403, x18239, x19402);
  nand n19404(x19404, x18238, x19401);
  nand n19405(x19405, x19404, x19403);
  nand n19407(x19407, x19399, x19403);
  nand n19408(x19408, x18241, x18243);
  nand n19409(x19409, x18240, x18242);
  nand n19410(x19410, x19409, x19408);
  nand n19412(x19412, x18245, x19411);
  nand n19413(x19413, x18244, x19410);
  nand n19414(x19414, x19413, x19412);
  nand n19415(x19415, x19408, x19412);
  nand n19416(x19416, x18247, x18249);
  nand n19417(x19417, x18246, x18248);
  nand n19418(x19418, x19417, x19416);
  nand n19420(x19420, x18251, x19419);
  nand n19421(x19421, x18250, x19418);
  nand n19422(x19422, x19421, x19420);
  nand n19424(x19424, x19416, x19420);
  nand n19425(x19425, x18253, x18255);
  nand n19426(x19426, x18252, x18254);
  nand n19427(x19427, x19426, x19425);
  nand n19429(x19429, x18257, x19428);
  nand n19430(x19430, x18256, x19427);
  nand n19431(x19431, x19430, x19429);
  nand n19433(x19433, x19425, x19429);
  nand n19434(x19434, x18259, x18261);
  nand n19435(x19435, x18258, x18260);
  nand n19436(x19436, x19435, x19434);
  nand n19438(x19438, x18263, x19437);
  nand n19439(x19439, x18262, x19436);
  nand n19440(x19440, x19439, x19438);
  nand n19442(x19442, x19434, x19438);
  nand n19443(x19443, x18265, x18267);
  nand n19444(x19444, x18264, x18266);
  nand n19445(x19445, x19444, x19443);
  nand n19447(x19447, x18269, x19446);
  nand n19448(x19448, x18268, x19445);
  nand n19449(x19449, x19448, x19447);
  nand n19451(x19451, x19443, x19447);
  nand n19452(x19452, x18271, x18273);
  nand n19453(x19453, x18270, x18272);
  nand n19454(x19454, x19453, x19452);
  nand n19456(x19456, x18275, x19455);
  nand n19457(x19457, x18274, x19454);
  nand n19458(x19458, x19457, x19456);
  nand n19460(x19460, x19452, x19456);
  nand n19461(x19461, x18278, x18280);
  nand n19462(x19462, x18277, x18279);
  nand n19463(x19463, x19462, x19461);
  nand n19465(x19465, x18282, x19464);
  nand n19466(x19466, x18281, x19463);
  nand n19467(x19467, x19466, x19465);
  nand n19468(x19468, x19461, x19465);
  nand n19469(x19469, x18284, x18286);
  nand n19470(x19470, x18283, x18285);
  nand n19471(x19471, x19470, x19469);
  nand n19473(x19473, x18288, x19472);
  nand n19474(x19474, x18287, x19471);
  nand n19475(x19475, x19474, x19473);
  nand n19477(x19477, x19469, x19473);
  nand n19478(x19478, x18290, x18292);
  nand n19479(x19479, x18289, x18291);
  nand n19480(x19480, x19479, x19478);
  nand n19482(x19482, x18294, x19481);
  nand n19483(x19483, x18293, x19480);
  nand n19484(x19484, x19483, x19482);
  nand n19486(x19486, x19478, x19482);
  nand n19487(x19487, x18296, x18298);
  nand n19488(x19488, x18295, x18297);
  nand n19489(x19489, x19488, x19487);
  nand n19491(x19491, x18300, x19490);
  nand n19492(x19492, x18299, x19489);
  nand n19493(x19493, x19492, x19491);
  nand n19495(x19495, x19487, x19491);
  nand n19496(x19496, x18302, x18304);
  nand n19497(x19497, x18301, x18303);
  nand n19498(x19498, x19497, x19496);
  nand n19500(x19500, x18306, x19499);
  nand n19501(x19501, x18305, x19498);
  nand n19502(x19502, x19501, x19500);
  nand n19504(x19504, x19496, x19500);
  nand n19505(x19505, x18308, x18310);
  nand n19506(x19506, x18307, x18309);
  nand n19507(x19507, x19506, x19505);
  nand n19509(x19509, x18312, x19508);
  nand n19510(x19510, x18311, x19507);
  nand n19511(x19511, x19510, x19509);
  nand n19513(x19513, x19505, x19509);
  nand n19514(x19514, x18314, x18316);
  nand n19515(x19515, x18313, x18315);
  nand n19516(x19516, x19515, x19514);
  nand n19517(x19517, x18318, x18320);
  nand n19518(x19518, x18317, x18319);
  nand n19519(x19519, x19518, x19517);
  nand n19521(x19521, x18322, x19520);
  nand n19522(x19522, x18321, x19519);
  nand n19523(x19523, x19522, x19521);
  nand n19524(x19524, x19517, x19521);
  nand n19525(x19525, x18324, x18326);
  nand n19526(x19526, x18323, x18325);
  nand n19527(x19527, x19526, x19525);
  nand n19529(x19529, x18328, x19528);
  nand n19530(x19530, x18327, x19527);
  nand n19531(x19531, x19530, x19529);
  nand n19533(x19533, x19525, x19529);
  nand n19534(x19534, x18330, x18332);
  nand n19535(x19535, x18329, x18331);
  nand n19536(x19536, x19535, x19534);
  nand n19538(x19538, x18334, x19537);
  nand n19539(x19539, x18333, x19536);
  nand n19540(x19540, x19539, x19538);
  nand n19542(x19542, x19534, x19538);
  nand n19543(x19543, x18336, x18338);
  nand n19544(x19544, x18335, x18337);
  nand n19545(x19545, x19544, x19543);
  nand n19547(x19547, x18340, x19546);
  nand n19548(x19548, x18339, x19545);
  nand n19549(x19549, x19548, x19547);
  nand n19551(x19551, x19543, x19547);
  nand n19552(x19552, x18342, x18344);
  nand n19553(x19553, x18341, x18343);
  nand n19554(x19554, x19553, x19552);
  nand n19556(x19556, x18346, x19555);
  nand n19557(x19557, x18345, x19554);
  nand n19558(x19558, x19557, x19556);
  nand n19560(x19560, x19552, x19556);
  nand n19561(x19561, x18348, x18350);
  nand n19562(x19562, x18347, x18349);
  nand n19563(x19563, x19562, x19561);
  nand n19565(x19565, x18352, x19564);
  nand n19566(x19566, x18351, x19563);
  nand n19567(x19567, x19566, x19565);
  nand n19569(x19569, x19561, x19565);
  nand n19570(x19570, x18354, x18356);
  nand n19571(x19571, x18353, x18355);
  nand n19572(x19572, x19571, x19570);
  nand n19574(x19574, x18358, x19573);
  nand n19575(x19575, x18357, x19572);
  nand n19576(x19576, x19575, x19574);
  nand n19578(x19578, x19570, x19574);
  nand n19579(x19579, x18360, x18362);
  nand n19580(x19580, x18359, x18361);
  nand n19581(x19581, x19580, x19579);
  nand n19583(x19583, x18364, x19582);
  nand n19584(x19584, x18363, x19581);
  nand n19585(x19585, x19584, x19583);
  nand n19586(x19586, x19579, x19583);
  nand n19587(x19587, x18366, x18368);
  nand n19588(x19588, x18365, x18367);
  nand n19589(x19589, x19588, x19587);
  nand n19591(x19591, x18370, x19590);
  nand n19592(x19592, x18369, x19589);
  nand n19593(x19593, x19592, x19591);
  nand n19595(x19595, x19587, x19591);
  nand n19596(x19596, x18372, x18374);
  nand n19597(x19597, x18371, x18373);
  nand n19598(x19598, x19597, x19596);
  nand n19600(x19600, x18376, x19599);
  nand n19601(x19601, x18375, x19598);
  nand n19602(x19602, x19601, x19600);
  nand n19604(x19604, x19596, x19600);
  nand n19605(x19605, x18378, x18380);
  nand n19606(x19606, x18377, x18379);
  nand n19607(x19607, x19606, x19605);
  nand n19609(x19609, x18382, x19608);
  nand n19610(x19610, x18381, x19607);
  nand n19611(x19611, x19610, x19609);
  nand n19613(x19613, x19605, x19609);
  nand n19614(x19614, x18384, x18386);
  nand n19615(x19615, x18383, x18385);
  nand n19616(x19616, x19615, x19614);
  nand n19618(x19618, x18388, x19617);
  nand n19619(x19619, x18387, x19616);
  nand n19620(x19620, x19619, x19618);
  nand n19622(x19622, x19614, x19618);
  nand n19623(x19623, x18390, x18392);
  nand n19624(x19624, x18389, x18391);
  nand n19625(x19625, x19624, x19623);
  nand n19627(x19627, x18394, x19626);
  nand n19628(x19628, x18393, x19625);
  nand n19629(x19629, x19628, x19627);
  nand n19631(x19631, x19623, x19627);
  nand n19632(x19632, x18396, x18398);
  nand n19633(x19633, x18395, x18397);
  nand n19634(x19634, x19633, x19632);
  nand n19636(x19636, x18400, x19635);
  nand n19637(x19637, x18399, x19634);
  nand n19638(x19638, x19637, x19636);
  nand n19640(x19640, x19632, x19636);
  nand n19641(x19641, x18403, x18405);
  nand n19642(x19642, x18402, x18404);
  nand n19643(x19643, x19642, x19641);
  nand n19645(x19645, x18407, x19644);
  nand n19646(x19646, x18406, x19643);
  nand n19647(x19647, x19646, x19645);
  nand n19648(x19648, x19641, x19645);
  nand n19649(x19649, x18409, x18411);
  nand n19650(x19650, x18408, x18410);
  nand n19651(x19651, x19650, x19649);
  nand n19653(x19653, x18413, x19652);
  nand n19654(x19654, x18412, x19651);
  nand n19655(x19655, x19654, x19653);
  nand n19657(x19657, x19649, x19653);
  nand n19658(x19658, x18415, x18417);
  nand n19659(x19659, x18414, x18416);
  nand n19660(x19660, x19659, x19658);
  nand n19662(x19662, x18419, x19661);
  nand n19663(x19663, x18418, x19660);
  nand n19664(x19664, x19663, x19662);
  nand n19666(x19666, x19658, x19662);
  nand n19667(x19667, x18421, x18423);
  nand n19668(x19668, x18420, x18422);
  nand n19669(x19669, x19668, x19667);
  nand n19671(x19671, x18425, x19670);
  nand n19672(x19672, x18424, x19669);
  nand n19673(x19673, x19672, x19671);
  nand n19675(x19675, x19667, x19671);
  nand n19676(x19676, x18427, x18429);
  nand n19677(x19677, x18426, x18428);
  nand n19678(x19678, x19677, x19676);
  nand n19680(x19680, x18431, x19679);
  nand n19681(x19681, x18430, x19678);
  nand n19682(x19682, x19681, x19680);
  nand n19684(x19684, x19676, x19680);
  nand n19685(x19685, x18433, x18435);
  nand n19686(x19686, x18432, x18434);
  nand n19687(x19687, x19686, x19685);
  nand n19689(x19689, x18437, x19688);
  nand n19690(x19690, x18436, x19687);
  nand n19691(x19691, x19690, x19689);
  nand n19693(x19693, x19685, x19689);
  nand n19694(x19694, x18439, x18441);
  nand n19695(x19695, x18438, x18440);
  nand n19696(x19696, x19695, x19694);
  nand n19698(x19698, x18443, x19697);
  nand n19699(x19699, x18442, x19696);
  nand n19700(x19700, x19699, x19698);
  nand n19702(x19702, x19694, x19698);
  nand n19703(x19703, x18445, x18447);
  nand n19704(x19704, x18444, x18446);
  nand n19705(x19705, x19704, x19703);
  nand n19706(x19706, x18449, x18451);
  nand n19707(x19707, x18448, x18450);
  nand n19708(x19708, x19707, x19706);
  nand n19710(x19710, x18453, x19709);
  nand n19711(x19711, x18452, x19708);
  nand n19712(x19712, x19711, x19710);
  nand n19713(x19713, x19706, x19710);
  nand n19714(x19714, x18455, x18457);
  nand n19715(x19715, x18454, x18456);
  nand n19716(x19716, x19715, x19714);
  nand n19718(x19718, x18459, x19717);
  nand n19719(x19719, x18458, x19716);
  nand n19720(x19720, x19719, x19718);
  nand n19722(x19722, x19714, x19718);
  nand n19723(x19723, x18461, x18463);
  nand n19724(x19724, x18460, x18462);
  nand n19725(x19725, x19724, x19723);
  nand n19727(x19727, x18465, x19726);
  nand n19728(x19728, x18464, x19725);
  nand n19729(x19729, x19728, x19727);
  nand n19731(x19731, x19723, x19727);
  nand n19732(x19732, x18467, x18469);
  nand n19733(x19733, x18466, x18468);
  nand n19734(x19734, x19733, x19732);
  nand n19736(x19736, x18471, x19735);
  nand n19737(x19737, x18470, x19734);
  nand n19738(x19738, x19737, x19736);
  nand n19740(x19740, x19732, x19736);
  nand n19741(x19741, x18473, x18475);
  nand n19742(x19742, x18472, x18474);
  nand n19743(x19743, x19742, x19741);
  nand n19745(x19745, x18477, x19744);
  nand n19746(x19746, x18476, x19743);
  nand n19747(x19747, x19746, x19745);
  nand n19749(x19749, x19741, x19745);
  nand n19750(x19750, x18479, x18481);
  nand n19751(x19751, x18478, x18480);
  nand n19752(x19752, x19751, x19750);
  nand n19754(x19754, x18483, x19753);
  nand n19755(x19755, x18482, x19752);
  nand n19756(x19756, x19755, x19754);
  nand n19758(x19758, x19750, x19754);
  nand n19759(x19759, x18485, x18487);
  nand n19760(x19760, x18484, x18486);
  nand n19761(x19761, x19760, x19759);
  nand n19763(x19763, x18489, x19762);
  nand n19764(x19764, x18488, x19761);
  nand n19765(x19765, x19764, x19763);
  nand n19767(x19767, x19759, x19763);
  nand n19768(x19768, x18491, x18493);
  nand n19769(x19769, x18490, x18492);
  nand n19770(x19770, x19769, x19768);
  nand n19772(x19772, x18495, x19771);
  nand n19773(x19773, x18494, x19770);
  nand n19774(x19774, x19773, x19772);
  nand n19775(x19775, x19768, x19772);
  nand n19776(x19776, x18497, x18499);
  nand n19777(x19777, x18496, x18498);
  nand n19778(x19778, x19777, x19776);
  nand n19780(x19780, x18501, x19779);
  nand n19781(x19781, x18500, x19778);
  nand n19782(x19782, x19781, x19780);
  nand n19783(x19783, x19776, x19780);
  nand n19784(x19784, x18503, x18505);
  nand n19785(x19785, x18502, x18504);
  nand n19786(x19786, x19785, x19784);
  nand n19788(x19788, x18507, x19787);
  nand n19789(x19789, x18506, x19786);
  nand n19790(x19790, x19789, x19788);
  nand n19792(x19792, x19784, x19788);
  nand n19793(x19793, x18509, x18511);
  nand n19794(x19794, x18508, x18510);
  nand n19795(x19795, x19794, x19793);
  nand n19797(x19797, x18513, x19796);
  nand n19798(x19798, x18512, x19795);
  nand n19799(x19799, x19798, x19797);
  nand n19801(x19801, x19793, x19797);
  nand n19802(x19802, x18515, x18517);
  nand n19803(x19803, x18514, x18516);
  nand n19804(x19804, x19803, x19802);
  nand n19806(x19806, x18519, x19805);
  nand n19807(x19807, x18518, x19804);
  nand n19808(x19808, x19807, x19806);
  nand n19810(x19810, x19802, x19806);
  nand n19811(x19811, x18521, x18523);
  nand n19812(x19812, x18520, x18522);
  nand n19813(x19813, x19812, x19811);
  nand n19815(x19815, x18525, x19814);
  nand n19816(x19816, x18524, x19813);
  nand n19817(x19817, x19816, x19815);
  nand n19819(x19819, x19811, x19815);
  nand n19820(x19820, x18527, x18529);
  nand n19821(x19821, x18526, x18528);
  nand n19822(x19822, x19821, x19820);
  nand n19824(x19824, x18531, x19823);
  nand n19825(x19825, x18530, x19822);
  nand n19826(x19826, x19825, x19824);
  nand n19828(x19828, x19820, x19824);
  nand n19829(x19829, x18533, x18535);
  nand n19830(x19830, x18532, x18534);
  nand n19831(x19831, x19830, x19829);
  nand n19833(x19833, x18537, x19832);
  nand n19834(x19834, x18536, x19831);
  nand n19835(x19835, x19834, x19833);
  nand n19837(x19837, x19829, x19833);
  nand n19838(x19838, x18539, x18541);
  nand n19839(x19839, x18538, x18540);
  nand n19840(x19840, x19839, x19838);
  nand n19842(x19842, x18543, x19841);
  nand n19843(x19843, x18542, x19840);
  nand n19844(x19844, x19843, x19842);
  nand n19846(x19846, x19838, x19842);
  nand n19847(x19847, x18546, x18548);
  nand n19848(x19848, x18545, x18547);
  nand n19849(x19849, x19848, x19847);
  nand n19851(x19851, x18550, x19850);
  nand n19852(x19852, x18549, x19849);
  nand n19853(x19853, x19852, x19851);
  nand n19854(x19854, x19847, x19851);
  nand n19855(x19855, x18552, x18554);
  nand n19856(x19856, x18551, x18553);
  nand n19857(x19857, x19856, x19855);
  nand n19859(x19859, x18556, x19858);
  nand n19860(x19860, x18555, x19857);
  nand n19861(x19861, x19860, x19859);
  nand n19863(x19863, x19855, x19859);
  nand n19864(x19864, x18558, x18560);
  nand n19865(x19865, x18557, x18559);
  nand n19866(x19866, x19865, x19864);
  nand n19868(x19868, x18562, x19867);
  nand n19869(x19869, x18561, x19866);
  nand n19870(x19870, x19869, x19868);
  nand n19872(x19872, x19864, x19868);
  nand n19873(x19873, x18564, x18566);
  nand n19874(x19874, x18563, x18565);
  nand n19875(x19875, x19874, x19873);
  nand n19877(x19877, x18568, x19876);
  nand n19878(x19878, x18567, x19875);
  nand n19879(x19879, x19878, x19877);
  nand n19881(x19881, x19873, x19877);
  nand n19882(x19882, x18570, x18572);
  nand n19883(x19883, x18569, x18571);
  nand n19884(x19884, x19883, x19882);
  nand n19886(x19886, x18574, x19885);
  nand n19887(x19887, x18573, x19884);
  nand n19888(x19888, x19887, x19886);
  nand n19890(x19890, x19882, x19886);
  nand n19891(x19891, x18576, x18578);
  nand n19892(x19892, x18575, x18577);
  nand n19893(x19893, x19892, x19891);
  nand n19895(x19895, x18580, x19894);
  nand n19896(x19896, x18579, x19893);
  nand n19897(x19897, x19896, x19895);
  nand n19899(x19899, x19891, x19895);
  nand n19900(x19900, x18582, x18584);
  nand n19901(x19901, x18581, x18583);
  nand n19902(x19902, x19901, x19900);
  nand n19904(x19904, x18586, x19903);
  nand n19905(x19905, x18585, x19902);
  nand n19906(x19906, x19905, x19904);
  nand n19908(x19908, x19900, x19904);
  nand n19909(x19909, x18588, x18590);
  nand n19910(x19910, x18587, x18589);
  nand n19911(x19911, x19910, x19909);
  nand n19913(x19913, x18592, x19912);
  nand n19914(x19914, x18591, x19911);
  nand n19915(x19915, x19914, x19913);
  nand n19917(x19917, x19909, x19913);
  nand n19918(x19918, x18594, x18596);
  nand n19919(x19919, x18593, x18595);
  nand n19920(x19920, x19919, x19918);
  nand n19921(x19921, x18598, x18600);
  nand n19922(x19922, x18597, x18599);
  nand n19923(x19923, x19922, x19921);
  nand n19925(x19925, x18602, x19924);
  nand n19926(x19926, x18601, x19923);
  nand n19927(x19927, x19926, x19925);
  nand n19928(x19928, x19921, x19925);
  nand n19929(x19929, x18604, x18606);
  nand n19930(x19930, x18603, x18605);
  nand n19931(x19931, x19930, x19929);
  nand n19933(x19933, x18608, x19932);
  nand n19934(x19934, x18607, x19931);
  nand n19935(x19935, x19934, x19933);
  nand n19937(x19937, x19929, x19933);
  nand n19938(x19938, x18610, x18612);
  nand n19939(x19939, x18609, x18611);
  nand n19940(x19940, x19939, x19938);
  nand n19942(x19942, x18614, x19941);
  nand n19943(x19943, x18613, x19940);
  nand n19944(x19944, x19943, x19942);
  nand n19946(x19946, x19938, x19942);
  nand n19947(x19947, x18616, x18618);
  nand n19948(x19948, x18615, x18617);
  nand n19949(x19949, x19948, x19947);
  nand n19951(x19951, x18620, x19950);
  nand n19952(x19952, x18619, x19949);
  nand n19953(x19953, x19952, x19951);
  nand n19955(x19955, x19947, x19951);
  nand n19956(x19956, x18622, x18624);
  nand n19957(x19957, x18621, x18623);
  nand n19958(x19958, x19957, x19956);
  nand n19960(x19960, x18626, x19959);
  nand n19961(x19961, x18625, x19958);
  nand n19962(x19962, x19961, x19960);
  nand n19964(x19964, x19956, x19960);
  nand n19965(x19965, x18628, x18630);
  nand n19966(x19966, x18627, x18629);
  nand n19967(x19967, x19966, x19965);
  nand n19969(x19969, x18632, x19968);
  nand n19970(x19970, x18631, x19967);
  nand n19971(x19971, x19970, x19969);
  nand n19973(x19973, x19965, x19969);
  nand n19974(x19974, x18634, x18636);
  nand n19975(x19975, x18633, x18635);
  nand n19976(x19976, x19975, x19974);
  nand n19978(x19978, x18638, x19977);
  nand n19979(x19979, x18637, x19976);
  nand n19980(x19980, x19979, x19978);
  nand n19982(x19982, x19974, x19978);
  nand n19983(x19983, x18640, x18642);
  nand n19984(x19984, x18639, x18641);
  nand n19985(x19985, x19984, x19983);
  nand n19987(x19987, x18644, x19986);
  nand n19988(x19988, x18643, x19985);
  nand n19989(x19989, x19988, x19987);
  nand n19991(x19991, x19983, x19987);
  nand n19992(x19992, x18646, x18648);
  nand n19993(x19993, x18645, x18647);
  nand n19994(x19994, x19993, x19992);
  nand n19996(x19996, x18650, x19995);
  nand n19997(x19997, x18649, x19994);
  nand n19998(x19998, x19997, x19996);
  nand n20000(x20000, x19992, x19996);
  nand n20001(x20001, x18652, x18654);
  nand n20002(x20002, x18651, x18653);
  nand n20003(x20003, x20002, x20001);
  nand n20005(x20005, x18656, x20004);
  nand n20006(x20006, x18655, x20003);
  nand n20007(x20007, x20006, x20005);
  nand n20008(x20008, x20001, x20005);
  nand n20009(x20009, x18658, x18660);
  nand n20010(x20010, x18657, x18659);
  nand n20011(x20011, x20010, x20009);
  nand n20013(x20013, x18662, x20012);
  nand n20014(x20014, x18661, x20011);
  nand n20015(x20015, x20014, x20013);
  nand n20017(x20017, x20009, x20013);
  nand n20018(x20018, x18664, x18666);
  nand n20019(x20019, x18663, x18665);
  nand n20020(x20020, x20019, x20018);
  nand n20022(x20022, x18668, x20021);
  nand n20023(x20023, x18667, x20020);
  nand n20024(x20024, x20023, x20022);
  nand n20026(x20026, x20018, x20022);
  nand n20027(x20027, x18670, x18672);
  nand n20028(x20028, x18669, x18671);
  nand n20029(x20029, x20028, x20027);
  nand n20031(x20031, x18674, x20030);
  nand n20032(x20032, x18673, x20029);
  nand n20033(x20033, x20032, x20031);
  nand n20035(x20035, x20027, x20031);
  nand n20036(x20036, x18676, x18678);
  nand n20037(x20037, x18675, x18677);
  nand n20038(x20038, x20037, x20036);
  nand n20040(x20040, x18680, x20039);
  nand n20041(x20041, x18679, x20038);
  nand n20042(x20042, x20041, x20040);
  nand n20044(x20044, x20036, x20040);
  nand n20045(x20045, x18682, x18684);
  nand n20046(x20046, x18681, x18683);
  nand n20047(x20047, x20046, x20045);
  nand n20049(x20049, x18686, x20048);
  nand n20050(x20050, x18685, x20047);
  nand n20051(x20051, x20050, x20049);
  nand n20053(x20053, x20045, x20049);
  nand n20054(x20054, x18688, x18690);
  nand n20055(x20055, x18687, x18689);
  nand n20056(x20056, x20055, x20054);
  nand n20058(x20058, x18692, x20057);
  nand n20059(x20059, x18691, x20056);
  nand n20060(x20060, x20059, x20058);
  nand n20062(x20062, x20054, x20058);
  nand n20063(x20063, x18694, x18696);
  nand n20064(x20064, x18693, x18695);
  nand n20065(x20065, x20064, x20063);
  nand n20067(x20067, x18698, x20066);
  nand n20068(x20068, x18697, x20065);
  nand n20069(x20069, x20068, x20067);
  nand n20071(x20071, x20063, x20067);
  nand n20072(x20072, x18700, x18702);
  nand n20073(x20073, x18699, x18701);
  nand n20074(x20074, x20073, x20072);
  nand n20076(x20076, x18704, x20075);
  nand n20077(x20077, x18703, x20074);
  nand n20078(x20078, x20077, x20076);
  nand n20080(x20080, x20072, x20076);
  nand n20081(x20081, x18707, x18709);
  nand n20082(x20082, x18706, x18708);
  nand n20083(x20083, x20082, x20081);
  nand n20085(x20085, x18711, x20084);
  nand n20086(x20086, x18710, x20083);
  nand n20087(x20087, x20086, x20085);
  nand n20088(x20088, x20081, x20085);
  nand n20089(x20089, x18713, x18715);
  nand n20090(x20090, x18712, x18714);
  nand n20091(x20091, x20090, x20089);
  nand n20093(x20093, x18717, x20092);
  nand n20094(x20094, x18716, x20091);
  nand n20095(x20095, x20094, x20093);
  nand n20097(x20097, x20089, x20093);
  nand n20098(x20098, x18719, x18721);
  nand n20099(x20099, x18718, x18720);
  nand n20100(x20100, x20099, x20098);
  nand n20102(x20102, x18723, x20101);
  nand n20103(x20103, x18722, x20100);
  nand n20104(x20104, x20103, x20102);
  nand n20106(x20106, x20098, x20102);
  nand n20107(x20107, x18725, x18727);
  nand n20108(x20108, x18724, x18726);
  nand n20109(x20109, x20108, x20107);
  nand n20111(x20111, x18729, x20110);
  nand n20112(x20112, x18728, x20109);
  nand n20113(x20113, x20112, x20111);
  nand n20115(x20115, x20107, x20111);
  nand n20116(x20116, x18731, x18733);
  nand n20117(x20117, x18730, x18732);
  nand n20118(x20118, x20117, x20116);
  nand n20120(x20120, x18735, x20119);
  nand n20121(x20121, x18734, x20118);
  nand n20122(x20122, x20121, x20120);
  nand n20124(x20124, x20116, x20120);
  nand n20125(x20125, x18737, x18739);
  nand n20126(x20126, x18736, x18738);
  nand n20127(x20127, x20126, x20125);
  nand n20129(x20129, x18741, x20128);
  nand n20130(x20130, x18740, x20127);
  nand n20131(x20131, x20130, x20129);
  nand n20133(x20133, x20125, x20129);
  nand n20134(x20134, x18743, x18745);
  nand n20135(x20135, x18742, x18744);
  nand n20136(x20136, x20135, x20134);
  nand n20138(x20138, x18747, x20137);
  nand n20139(x20139, x18746, x20136);
  nand n20140(x20140, x20139, x20138);
  nand n20142(x20142, x20134, x20138);
  nand n20143(x20143, x18749, x18751);
  nand n20144(x20144, x18748, x18750);
  nand n20145(x20145, x20144, x20143);
  nand n20147(x20147, x18753, x20146);
  nand n20148(x20148, x18752, x20145);
  nand n20149(x20149, x20148, x20147);
  nand n20151(x20151, x20143, x20147);
  nand n20152(x20152, x18755, x18757);
  nand n20153(x20153, x18754, x18756);
  nand n20154(x20154, x20153, x20152);
  nand n20156(x20156, x18759, x20155);
  nand n20157(x20157, x18758, x20154);
  nand n20158(x20158, x20157, x20156);
  nand n20160(x20160, x20152, x20156);
  nand n20161(x20161, x18761, x18763);
  nand n20162(x20162, x18760, x18762);
  nand n20163(x20163, x20162, x20161);
  nand n20164(x20164, x18765, x18767);
  nand n20165(x20165, x18764, x18766);
  nand n20166(x20166, x20165, x20164);
  nand n20168(x20168, x18769, x20167);
  nand n20169(x20169, x18768, x20166);
  nand n20170(x20170, x20169, x20168);
  nand n20172(x20172, x20164, x20168);
  nand n20173(x20173, x18771, x18773);
  nand n20174(x20174, x18770, x18772);
  nand n20175(x20175, x20174, x20173);
  nand n20177(x20177, x18775, x20176);
  nand n20178(x20178, x18774, x20175);
  nand n20179(x20179, x20178, x20177);
  nand n20181(x20181, x20173, x20177);
  nand n20182(x20182, x18777, x18779);
  nand n20183(x20183, x18776, x18778);
  nand n20184(x20184, x20183, x20182);
  nand n20186(x20186, x18781, x20185);
  nand n20187(x20187, x18780, x20184);
  nand n20188(x20188, x20187, x20186);
  nand n20190(x20190, x20182, x20186);
  nand n20191(x20191, x18783, x18785);
  nand n20192(x20192, x18782, x18784);
  nand n20193(x20193, x20192, x20191);
  nand n20195(x20195, x18787, x20194);
  nand n20196(x20196, x18786, x20193);
  nand n20197(x20197, x20196, x20195);
  nand n20199(x20199, x20191, x20195);
  nand n20200(x20200, x18789, x18791);
  nand n20201(x20201, x18788, x18790);
  nand n20202(x20202, x20201, x20200);
  nand n20204(x20204, x18793, x20203);
  nand n20205(x20205, x18792, x20202);
  nand n20206(x20206, x20205, x20204);
  nand n20208(x20208, x20200, x20204);
  nand n20209(x20209, x18795, x18797);
  nand n20210(x20210, x18794, x18796);
  nand n20211(x20211, x20210, x20209);
  nand n20213(x20213, x18799, x20212);
  nand n20214(x20214, x18798, x20211);
  nand n20215(x20215, x20214, x20213);
  nand n20217(x20217, x20209, x20213);
  nand n20218(x20218, x18801, x18803);
  nand n20219(x20219, x18800, x18802);
  nand n20220(x20220, x20219, x20218);
  nand n20222(x20222, x18805, x20221);
  nand n20223(x20223, x18804, x20220);
  nand n20224(x20224, x20223, x20222);
  nand n20226(x20226, x20218, x20222);
  nand n20227(x20227, x18807, x18809);
  nand n20228(x20228, x18806, x18808);
  nand n20229(x20229, x20228, x20227);
  nand n20231(x20231, x18811, x20230);
  nand n20232(x20232, x18810, x20229);
  nand n20233(x20233, x20232, x20231);
  nand n20235(x20235, x20227, x20231);
  nand n20236(x20236, x18813, x18815);
  nand n20237(x20237, x18812, x18814);
  nand n20238(x20238, x20237, x20236);
  nand n20240(x20240, x18817, x20239);
  nand n20241(x20241, x18816, x20238);
  nand n20242(x20242, x20241, x20240);
  nand n20244(x20244, x20236, x20240);
  nand n20245(x20245, x18819, x18821);
  nand n20246(x20246, x18818, x18820);
  nand n20247(x20247, x20246, x20245);
  nand n20249(x20249, x18823, x20248);
  nand n20250(x20250, x18822, x20247);
  nand n20251(x20251, x20250, x20249);
  nand n20253(x20253, x20245, x20249);
  nand n20254(x20254, x18825, x18827);
  nand n20255(x20255, x18824, x18826);
  nand n20256(x20256, x20255, x20254);
  nand n20258(x20258, x18829, x20257);
  nand n20259(x20259, x18828, x20256);
  nand n20260(x20260, x20259, x20258);
  nand n20262(x20262, x20254, x20258);
  nand n20263(x20263, x18831, x18833);
  nand n20264(x20264, x18830, x18832);
  nand n20265(x20265, x20264, x20263);
  nand n20267(x20267, x18835, x20266);
  nand n20268(x20268, x18834, x20265);
  nand n20269(x20269, x20268, x20267);
  nand n20271(x20271, x20263, x20267);
  nand n20272(x20272, x18837, x18839);
  nand n20273(x20273, x18836, x18838);
  nand n20274(x20274, x20273, x20272);
  nand n20276(x20276, x18841, x20275);
  nand n20277(x20277, x18840, x20274);
  nand n20278(x20278, x20277, x20276);
  nand n20280(x20280, x20272, x20276);
  nand n20281(x20281, x18843, x18845);
  nand n20282(x20282, x18842, x18844);
  nand n20283(x20283, x20282, x20281);
  nand n20285(x20285, x18847, x20284);
  nand n20286(x20286, x18846, x20283);
  nand n20287(x20287, x20286, x20285);
  nand n20289(x20289, x20281, x20285);
  nand n20290(x20290, x18849, x18851);
  nand n20291(x20291, x18848, x18850);
  nand n20292(x20292, x20291, x20290);
  nand n20294(x20294, x18853, x20293);
  nand n20295(x20295, x18852, x20292);
  nand n20296(x20296, x20295, x20294);
  nand n20298(x20298, x20290, x20294);
  nand n20299(x20299, x18855, x18857);
  nand n20300(x20300, x18854, x18856);
  nand n20301(x20301, x20300, x20299);
  nand n20303(x20303, x18859, x20302);
  nand n20304(x20304, x18858, x20301);
  nand n20305(x20305, x20304, x20303);
  nand n20307(x20307, x20299, x20303);
  nand n20308(x20308, x18861, x18863);
  nand n20309(x20309, x18860, x18862);
  nand n20310(x20310, x20309, x20308);
  nand n20312(x20312, x18865, x20311);
  nand n20313(x20313, x18864, x20310);
  nand n20314(x20314, x20313, x20312);
  nand n20316(x20316, x20308, x20312);
  nand n20317(x20317, x18867, x18869);
  nand n20318(x20318, x18866, x18868);
  nand n20319(x20319, x20318, x20317);
  nand n20321(x20321, x18871, x20320);
  nand n20322(x20322, x18870, x20319);
  nand n20323(x20323, x20322, x20321);
  nand n20325(x20325, x20317, x20321);
  nand n20326(x20326, x18873, x18875);
  nand n20327(x20327, x18872, x18874);
  nand n20328(x20328, x20327, x20326);
  nand n20330(x20330, x18877, x20329);
  nand n20331(x20331, x18876, x20328);
  nand n20332(x20332, x20331, x20330);
  nand n20334(x20334, x20326, x20330);
  nand n20335(x20335, x18879, x18881);
  nand n20336(x20336, x18878, x18880);
  nand n20337(x20337, x20336, x20335);
  nand n20339(x20339, x18883, x20338);
  nand n20340(x20340, x18882, x20337);
  nand n20341(x20341, x20340, x20339);
  nand n20343(x20343, x20335, x20339);
  nand n20344(x20344, x18886, x18888);
  nand n20345(x20345, x18885, x18887);
  nand n20346(x20346, x20345, x20344);
  nand n20348(x20348, x18890, x20347);
  nand n20349(x20349, x18889, x20346);
  nand n20350(x20350, x20349, x20348);
  nand n20352(x20352, x18892, x18894);
  nand n20353(x20353, x18891, x18893);
  nand n20354(x20354, x20353, x20352);
  nand n20356(x20356, x18896, x20355);
  nand n20357(x20357, x18895, x20354);
  nand n20358(x20358, x20357, x20356);
  nand n20360(x20360, x18898, x18900);
  nand n20361(x20361, x18897, x18899);
  nand n20362(x20362, x20361, x20360);
  nand n20364(x20364, x18902, x20363);
  nand n20365(x20365, x18901, x20362);
  nand n20366(x20366, x20365, x20364);
  nand n20368(x20368, x18904, x18906);
  nand n20369(x20369, x18903, x18905);
  nand n20370(x20370, x20369, x20368);
  nand n20372(x20372, x18908, x20371);
  nand n20373(x20373, x18907, x20370);
  nand n20374(x20374, x20373, x20372);
  nand n20376(x20376, x18910, x18912);
  nand n20377(x20377, x18909, x18911);
  nand n20378(x20378, x20377, x20376);
  nand n20380(x20380, x18914, x20379);
  nand n20381(x20381, x18913, x20378);
  nand n20382(x20382, x20381, x20380);
  nand n20384(x20384, x18916, x18918);
  nand n20385(x20385, x18915, x18917);
  nand n20386(x20386, x20385, x20384);
  nand n20388(x20388, x18920, x20387);
  nand n20389(x20389, x18919, x20386);
  nand n20390(x20390, x20389, x20388);
  nand n20392(x20392, x18922, x18924);
  nand n20393(x20393, x18921, x18923);
  nand n20394(x20394, x20393, x20392);
  nand n20396(x20396, x18926, x20395);
  nand n20397(x20397, x18925, x20394);
  nand n20398(x20398, x20397, x20396);
  nand n20400(x20400, x18928, x18930);
  nand n20401(x20401, x18927, x18929);
  nand n20402(x20402, x20401, x20400);
  nand n20404(x20404, x18932, x20403);
  nand n20405(x20405, x18931, x20402);
  nand n20406(x20406, x20405, x20404);
  nand n20408(x20408, x18934, x18936);
  nand n20409(x20409, x18933, x18935);
  nand n20410(x20410, x20409, x20408);
  nand n20412(x20412, x18938, x20411);
  nand n20413(x20413, x18937, x20410);
  nand n20414(x20414, x20413, x20412);
  nand n20416(x20416, x18940, x18942);
  nand n20417(x20417, x18939, x18941);
  nand n20418(x20418, x20417, x20416);
  nand n20420(x20420, x18944, x20419);
  nand n20421(x20421, x18943, x20418);
  nand n20422(x20422, x20421, x20420);
  nand n20424(x20424, x18946, x18948);
  nand n20425(x20425, x18945, x18947);
  nand n20426(x20426, x20425, x20424);
  nand n20430(x20430, x18975, x83575);
  nand n20432(x20432, x20431, x18976);
  nand n20433(x20433, x20432, x20430);
  nand n20434(x20434, x18986, x18994);
  nand n20437(x20437, x20436, x20435);
  nand n20438(x20438, x20437, x20434);
  nand n20439(x20439, x19010, x83576);
  nand n20440(x20440, x19009, x17956);
  nand n20441(x20441, x20440, x20439);
  nand n20442(x20442, x19002, x19011);
  nand n20445(x20445, x20444, x20443);
  nand n20446(x20446, x20445, x20442);
  nand n20447(x20447, x19027, x83577);
  nand n20448(x20448, x19026, x19031);
  nand n20449(x20449, x20448, x20447);
  nand n20450(x20450, x19019, x19028);
  nand n20453(x20453, x20452, x20451);
  nand n20454(x20454, x20453, x20450);
  nand n20456(x20456, x83578, x20455);
  nand n20457(x20457, x19029, x20454);
  nand n20458(x20458, x20457, x20456);
  nand n20459(x20459, x20450, x20456);
  nand n20460(x20460, x19047, x19056);
  nand n20461(x20461, x19046, x19055);
  nand n20462(x20462, x20461, x20460);
  nand n20463(x20463, x19039, x19048);
  nand n20466(x20466, x20465, x20464);
  nand n20467(x20467, x20466, x20463);
  nand n20469(x20469, x19057, x20468);
  nand n20471(x20471, x20470, x20467);
  nand n20472(x20472, x20471, x20469);
  nand n20473(x20473, x20463, x20469);
  nand n20474(x20474, x19073, x19082);
  nand n20475(x20475, x19072, x19081);
  nand n20476(x20476, x20475, x20474);
  nand n20478(x20478, x83579, x20477);
  nand n20479(x20479, x18009, x20476);
  nand n20480(x20480, x20479, x20478);
  nand n20482(x20482, x20474, x20478);
  nand n20483(x20483, x19065, x19074);
  nand n20486(x20486, x20485, x20484);
  nand n20487(x20487, x20486, x20483);
  nand n20489(x20489, x19083, x20488);
  nand n20491(x20491, x20490, x20487);
  nand n20492(x20492, x20491, x20489);
  nand n20493(x20493, x20483, x20489);
  nand n20494(x20494, x19099, x19108);
  nand n20495(x20495, x19098, x19107);
  nand n20496(x20496, x20495, x20494);
  nand n20498(x20498, x83580, x20497);
  nand n20499(x20499, x19112, x20496);
  nand n20500(x20500, x20499, x20498);
  nand n20502(x20502, x20494, x20498);
  nand n20503(x20503, x19091, x19100);
  nand n20506(x20506, x20505, x20504);
  nand n20507(x20507, x20506, x20503);
  nand n20509(x20509, x19109, x20508);
  nand n20511(x20511, x20510, x20507);
  nand n20512(x20512, x20511, x20509);
  nand n20513(x20513, x20503, x20509);
  nand n20514(x20514, x19128, x19137);
  nand n20515(x20515, x19127, x19136);
  nand n20516(x20516, x20515, x20514);
  nand n20518(x20518, x19146, x20517);
  nand n20519(x20519, x19145, x20516);
  nand n20520(x20520, x20519, x20518);
  nand n20522(x20522, x20514, x20518);
  nand n20523(x20523, x19120, x19129);
  nand n20526(x20526, x20525, x20524);
  nand n20527(x20527, x20526, x20523);
  nand n20529(x20529, x19138, x20528);
  nand n20531(x20531, x20530, x20527);
  nand n20532(x20532, x20531, x20529);
  nand n20533(x20533, x20523, x20529);
  nand n20535(x20535, x19163, x19172);
  nand n20536(x20536, x19162, x19171);
  nand n20537(x20537, x20536, x20535);
  nand n20539(x20539, x19181, x20538);
  nand n20540(x20540, x19180, x20537);
  nand n20541(x20541, x20540, x20539);
  nand n20543(x20543, x20535, x20539);
  nand n20544(x20544, x19155, x19164);
  nand n20547(x20547, x20546, x20545);
  nand n20548(x20548, x20547, x20544);
  nand n20550(x20550, x19173, x20549);
  nand n20552(x20552, x20551, x20548);
  nand n20553(x20553, x20552, x20550);
  nand n20554(x20554, x20544, x20550);
  nand n20556(x20556, x19198, x19207);
  nand n20557(x20557, x19197, x19206);
  nand n20558(x20558, x20557, x20556);
  nand n20560(x20560, x19216, x20559);
  nand n20561(x20561, x19215, x20558);
  nand n20562(x20562, x20561, x20560);
  nand n20564(x20564, x20556, x20560);
  nand n20565(x20565, x19190, x19199);
  nand n20568(x20568, x20567, x20566);
  nand n20569(x20569, x20568, x20565);
  nand n20571(x20571, x19208, x20570);
  nand n20573(x20573, x20572, x20569);
  nand n20574(x20574, x20573, x20571);
  nand n20575(x20575, x20565, x20571);
  nand n20576(x20576, x19217, x83581);
  nand n20578(x20578, x20577, x19218);
  nand n20579(x20579, x20578, x20576);
  nand n20580(x20580, x19236, x19245);
  nand n20581(x20581, x19235, x19244);
  nand n20582(x20582, x20581, x20580);
  nand n20584(x20584, x19254, x20583);
  nand n20585(x20585, x19253, x20582);
  nand n20586(x20586, x20585, x20584);
  nand n20588(x20588, x20580, x20584);
  nand n20589(x20589, x19228, x19237);
  nand n20592(x20592, x20591, x20590);
  nand n20593(x20593, x20592, x20589);
  nand n20595(x20595, x19246, x20594);
  nand n20597(x20597, x20596, x20593);
  nand n20598(x20598, x20597, x20595);
  nand n20599(x20599, x20589, x20595);
  nand n20600(x20600, x19255, x19263);
  nand n20603(x20603, x20602, x20601);
  nand n20604(x20604, x20603, x20600);
  nand n20605(x20605, x19279, x19288);
  nand n20606(x20606, x19278, x19287);
  nand n20607(x20607, x20606, x20605);
  nand n20609(x20609, x19297, x20608);
  nand n20610(x20610, x19296, x20607);
  nand n20611(x20611, x20610, x20609);
  nand n20613(x20613, x20605, x20609);
  nand n20614(x20614, x19306, x83582);
  nand n20615(x20615, x19305, x18169);
  nand n20616(x20616, x20615, x20614);
  nand n20617(x20617, x19271, x19280);
  nand n20620(x20620, x20619, x20618);
  nand n20621(x20621, x20620, x20617);
  nand n20623(x20623, x19289, x20622);
  nand n20625(x20625, x20624, x20621);
  nand n20626(x20626, x20625, x20623);
  nand n20627(x20627, x20617, x20623);
  nand n20628(x20628, x19298, x19307);
  nand n20631(x20631, x20630, x20629);
  nand n20632(x20632, x20631, x20628);
  nand n20633(x20633, x19323, x19332);
  nand n20634(x20634, x19322, x19331);
  nand n20635(x20635, x20634, x20633);
  nand n20637(x20637, x19341, x20636);
  nand n20638(x20638, x19340, x20635);
  nand n20639(x20639, x20638, x20637);
  nand n20641(x20641, x20633, x20637);
  nand n20642(x20642, x19350, x83583);
  nand n20643(x20643, x19349, x19354);
  nand n20644(x20644, x20643, x20642);
  nand n20645(x20645, x19315, x19324);
  nand n20648(x20648, x20647, x20646);
  nand n20649(x20649, x20648, x20645);
  nand n20651(x20651, x19333, x20650);
  nand n20653(x20653, x20652, x20649);
  nand n20654(x20654, x20653, x20651);
  nand n20655(x20655, x20645, x20651);
  nand n20656(x20656, x19342, x19351);
  nand n20659(x20659, x20658, x20657);
  nand n20660(x20660, x20659, x20656);
  nand n20662(x20662, x83584, x20661);
  nand n20663(x20663, x19352, x20660);
  nand n20664(x20664, x20663, x20662);
  nand n20666(x20666, x20656, x20662);
  nand n20667(x20667, x19370, x19379);
  nand n20668(x20668, x19369, x19378);
  nand n20669(x20669, x20668, x20667);
  nand n20671(x20671, x19388, x20670);
  nand n20672(x20672, x19387, x20669);
  nand n20673(x20673, x20672, x20671);
  nand n20675(x20675, x20667, x20671);
  nand n20676(x20676, x19397, x19406);
  nand n20677(x20677, x19396, x19405);
  nand n20678(x20678, x20677, x20676);
  nand n20679(x20679, x19362, x19371);
  nand n20682(x20682, x20681, x20680);
  nand n20683(x20683, x20682, x20679);
  nand n20685(x20685, x19380, x20684);
  nand n20687(x20687, x20686, x20683);
  nand n20688(x20688, x20687, x20685);
  nand n20689(x20689, x20679, x20685);
  nand n20690(x20690, x19389, x19398);
  nand n20693(x20693, x20692, x20691);
  nand n20694(x20694, x20693, x20690);
  nand n20696(x20696, x19407, x20695);
  nand n20698(x20698, x20697, x20694);
  nand n20699(x20699, x20698, x20696);
  nand n20701(x20701, x20690, x20696);
  nand n20702(x20702, x19423, x19432);
  nand n20703(x20703, x19422, x19431);
  nand n20704(x20704, x20703, x20702);
  nand n20706(x20706, x19441, x20705);
  nand n20707(x20707, x19440, x20704);
  nand n20708(x20708, x20707, x20706);
  nand n20710(x20710, x20702, x20706);
  nand n20711(x20711, x19450, x19459);
  nand n20712(x20712, x19449, x19458);
  nand n20713(x20713, x20712, x20711);
  nand n20715(x20715, x83585, x20714);
  nand n20716(x20716, x18276, x20713);
  nand n20717(x20717, x20716, x20715);
  nand n20718(x20718, x20711, x20715);
  nand n20719(x20719, x19415, x19424);
  nand n20722(x20722, x20721, x20720);
  nand n20723(x20723, x20722, x20719);
  nand n20725(x20725, x19433, x20724);
  nand n20727(x20727, x20726, x20723);
  nand n20728(x20728, x20727, x20725);
  nand n20729(x20729, x20719, x20725);
  nand n20730(x20730, x19442, x19451);
  nand n20733(x20733, x20732, x20731);
  nand n20734(x20734, x20733, x20730);
  nand n20736(x20736, x19460, x20735);
  nand n20738(x20738, x20737, x20734);
  nand n20739(x20739, x20738, x20736);
  nand n20741(x20741, x20730, x20736);
  nand n20742(x20742, x19476, x19485);
  nand n20743(x20743, x19475, x19484);
  nand n20744(x20744, x20743, x20742);
  nand n20746(x20746, x19494, x20745);
  nand n20747(x20747, x19493, x20744);
  nand n20748(x20748, x20747, x20746);
  nand n20750(x20750, x20742, x20746);
  nand n20751(x20751, x19503, x19512);
  nand n20752(x20752, x19502, x19511);
  nand n20753(x20753, x20752, x20751);
  nand n20755(x20755, x83586, x20754);
  nand n20756(x20756, x19516, x20753);
  nand n20757(x20757, x20756, x20755);
  nand n20758(x20758, x20751, x20755);
  nand n20759(x20759, x19468, x19477);
  nand n20762(x20762, x20761, x20760);
  nand n20763(x20763, x20762, x20759);
  nand n20765(x20765, x19486, x20764);
  nand n20767(x20767, x20766, x20763);
  nand n20768(x20768, x20767, x20765);
  nand n20769(x20769, x20759, x20765);
  nand n20770(x20770, x19495, x19504);
  nand n20773(x20773, x20772, x20771);
  nand n20774(x20774, x20773, x20770);
  nand n20776(x20776, x19513, x20775);
  nand n20778(x20778, x20777, x20774);
  nand n20779(x20779, x20778, x20776);
  nand n20781(x20781, x20770, x20776);
  nand n20782(x20782, x19532, x19541);
  nand n20783(x20783, x19531, x19540);
  nand n20784(x20784, x20783, x20782);
  nand n20786(x20786, x19550, x20785);
  nand n20787(x20787, x19549, x20784);
  nand n20788(x20788, x20787, x20786);
  nand n20790(x20790, x20782, x20786);
  nand n20791(x20791, x19559, x19568);
  nand n20792(x20792, x19558, x19567);
  nand n20793(x20793, x20792, x20791);
  nand n20795(x20795, x19577, x20794);
  nand n20796(x20796, x19576, x20793);
  nand n20797(x20797, x20796, x20795);
  nand n20798(x20798, x20791, x20795);
  nand n20799(x20799, x19524, x19533);
  nand n20802(x20802, x20801, x20800);
  nand n20803(x20803, x20802, x20799);
  nand n20805(x20805, x19542, x20804);
  nand n20807(x20807, x20806, x20803);
  nand n20808(x20808, x20807, x20805);
  nand n20809(x20809, x20799, x20805);
  nand n20810(x20810, x19551, x19560);
  nand n20813(x20813, x20812, x20811);
  nand n20814(x20814, x20813, x20810);
  nand n20816(x20816, x19569, x20815);
  nand n20818(x20818, x20817, x20814);
  nand n20819(x20819, x20818, x20816);
  nand n20821(x20821, x20810, x20816);
  nand n20823(x20823, x19594, x19603);
  nand n20824(x20824, x19593, x19602);
  nand n20825(x20825, x20824, x20823);
  nand n20827(x20827, x19612, x20826);
  nand n20828(x20828, x19611, x20825);
  nand n20829(x20829, x20828, x20827);
  nand n20831(x20831, x20823, x20827);
  nand n20832(x20832, x19621, x19630);
  nand n20833(x20833, x19620, x19629);
  nand n20834(x20834, x20833, x20832);
  nand n20836(x20836, x19639, x20835);
  nand n20837(x20837, x19638, x20834);
  nand n20838(x20838, x20837, x20836);
  nand n20840(x20840, x20832, x20836);
  nand n20841(x20841, x19586, x19595);
  nand n20844(x20844, x20843, x20842);
  nand n20845(x20845, x20844, x20841);
  nand n20847(x20847, x19604, x20846);
  nand n20849(x20849, x20848, x20845);
  nand n20850(x20850, x20849, x20847);
  nand n20851(x20851, x20841, x20847);
  nand n20852(x20852, x19613, x19622);
  nand n20855(x20855, x20854, x20853);
  nand n20856(x20856, x20855, x20852);
  nand n20858(x20858, x19631, x20857);
  nand n20860(x20860, x20859, x20856);
  nand n20861(x20861, x20860, x20858);
  nand n20863(x20863, x20852, x20858);
  nand n20865(x20865, x19656, x19665);
  nand n20866(x20866, x19655, x19664);
  nand n20867(x20867, x20866, x20865);
  nand n20869(x20869, x19674, x20868);
  nand n20870(x20870, x19673, x20867);
  nand n20871(x20871, x20870, x20869);
  nand n20873(x20873, x20865, x20869);
  nand n20874(x20874, x19683, x19692);
  nand n20875(x20875, x19682, x19691);
  nand n20876(x20876, x20875, x20874);
  nand n20878(x20878, x19701, x20877);
  nand n20879(x20879, x19700, x20876);
  nand n20880(x20880, x20879, x20878);
  nand n20882(x20882, x20874, x20878);
  nand n20883(x20883, x19648, x19657);
  nand n20886(x20886, x20885, x20884);
  nand n20887(x20887, x20886, x20883);
  nand n20889(x20889, x19666, x20888);
  nand n20891(x20891, x20890, x20887);
  nand n20892(x20892, x20891, x20889);
  nand n20893(x20893, x20883, x20889);
  nand n20894(x20894, x19675, x19684);
  nand n20897(x20897, x20896, x20895);
  nand n20898(x20898, x20897, x20894);
  nand n20900(x20900, x19693, x20899);
  nand n20902(x20902, x20901, x20898);
  nand n20903(x20903, x20902, x20900);
  nand n20905(x20905, x20894, x20900);
  nand n20906(x20906, x19702, x83587);
  nand n20908(x20908, x20907, x19703);
  nand n20909(x20909, x20908, x20906);
  nand n20910(x20910, x19721, x19730);
  nand n20911(x20911, x19720, x19729);
  nand n20912(x20912, x20911, x20910);
  nand n20914(x20914, x19739, x20913);
  nand n20915(x20915, x19738, x20912);
  nand n20916(x20916, x20915, x20914);
  nand n20918(x20918, x20910, x20914);
  nand n20919(x20919, x19748, x19757);
  nand n20920(x20920, x19747, x19756);
  nand n20921(x20921, x20920, x20919);
  nand n20923(x20923, x19766, x20922);
  nand n20924(x20924, x19765, x20921);
  nand n20925(x20925, x20924, x20923);
  nand n20927(x20927, x20919, x20923);
  nand n20928(x20928, x19713, x19722);
  nand n20931(x20931, x20930, x20929);
  nand n20932(x20932, x20931, x20928);
  nand n20934(x20934, x19731, x20933);
  nand n20936(x20936, x20935, x20932);
  nand n20937(x20937, x20936, x20934);
  nand n20938(x20938, x20928, x20934);
  nand n20939(x20939, x19740, x19749);
  nand n20942(x20942, x20941, x20940);
  nand n20943(x20943, x20942, x20939);
  nand n20945(x20945, x19758, x20944);
  nand n20947(x20947, x20946, x20943);
  nand n20948(x20948, x20947, x20945);
  nand n20950(x20950, x20939, x20945);
  nand n20951(x20951, x19767, x19775);
  nand n20954(x20954, x20953, x20952);
  nand n20955(x20955, x20954, x20951);
  nand n20956(x20956, x19791, x19800);
  nand n20957(x20957, x19790, x19799);
  nand n20958(x20958, x20957, x20956);
  nand n20960(x20960, x19809, x20959);
  nand n20961(x20961, x19808, x20958);
  nand n20962(x20962, x20961, x20960);
  nand n20964(x20964, x20956, x20960);
  nand n20965(x20965, x19818, x19827);
  nand n20966(x20966, x19817, x19826);
  nand n20967(x20967, x20966, x20965);
  nand n20969(x20969, x19836, x20968);
  nand n20970(x20970, x19835, x20967);
  nand n20971(x20971, x20970, x20969);
  nand n20973(x20973, x20965, x20969);
  nand n20974(x20974, x19845, x83588);
  nand n20975(x20975, x19844, x18544);
  nand n20976(x20976, x20975, x20974);
  nand n20977(x20977, x19783, x19792);
  nand n20980(x20980, x20979, x20978);
  nand n20981(x20981, x20980, x20977);
  nand n20983(x20983, x19801, x20982);
  nand n20985(x20985, x20984, x20981);
  nand n20986(x20986, x20985, x20983);
  nand n20988(x20988, x20977, x20983);
  nand n20989(x20989, x19810, x19819);
  nand n20992(x20992, x20991, x20990);
  nand n20993(x20993, x20992, x20989);
  nand n20995(x20995, x19828, x20994);
  nand n20997(x20997, x20996, x20993);
  nand n20998(x20998, x20997, x20995);
  nand n21000(x21000, x20989, x20995);
  nand n21001(x21001, x19837, x19846);
  nand n21004(x21004, x21003, x21002);
  nand n21005(x21005, x21004, x21001);
  nand n21006(x21006, x19862, x19871);
  nand n21007(x21007, x19861, x19870);
  nand n21008(x21008, x21007, x21006);
  nand n21010(x21010, x19880, x21009);
  nand n21011(x21011, x19879, x21008);
  nand n21012(x21012, x21011, x21010);
  nand n21014(x21014, x21006, x21010);
  nand n21015(x21015, x19889, x19898);
  nand n21016(x21016, x19888, x19897);
  nand n21017(x21017, x21016, x21015);
  nand n21019(x21019, x19907, x21018);
  nand n21020(x21020, x19906, x21017);
  nand n21021(x21021, x21020, x21019);
  nand n21023(x21023, x21015, x21019);
  nand n21024(x21024, x19916, x83589);
  nand n21025(x21025, x19915, x19920);
  nand n21026(x21026, x21025, x21024);
  nand n21027(x21027, x19854, x19863);
  nand n21030(x21030, x21029, x21028);
  nand n21031(x21031, x21030, x21027);
  nand n21033(x21033, x19872, x21032);
  nand n21035(x21035, x21034, x21031);
  nand n21036(x21036, x21035, x21033);
  nand n21038(x21038, x21027, x21033);
  nand n21039(x21039, x19881, x19890);
  nand n21042(x21042, x21041, x21040);
  nand n21043(x21043, x21042, x21039);
  nand n21045(x21045, x19899, x21044);
  nand n21047(x21047, x21046, x21043);
  nand n21048(x21048, x21047, x21045);
  nand n21050(x21050, x21039, x21045);
  nand n21051(x21051, x19908, x19917);
  nand n21054(x21054, x21053, x21052);
  nand n21055(x21055, x21054, x21051);
  nand n21057(x21057, x83590, x21056);
  nand n21058(x21058, x19918, x21055);
  nand n21059(x21059, x21058, x21057);
  nand n21061(x21061, x21051, x21057);
  nand n21062(x21062, x19936, x19945);
  nand n21063(x21063, x19935, x19944);
  nand n21064(x21064, x21063, x21062);
  nand n21066(x21066, x19954, x21065);
  nand n21067(x21067, x19953, x21064);
  nand n21068(x21068, x21067, x21066);
  nand n21070(x21070, x21062, x21066);
  nand n21071(x21071, x19963, x19972);
  nand n21072(x21072, x19962, x19971);
  nand n21073(x21073, x21072, x21071);
  nand n21075(x21075, x19981, x21074);
  nand n21076(x21076, x19980, x21073);
  nand n21077(x21077, x21076, x21075);
  nand n21079(x21079, x21071, x21075);
  nand n21080(x21080, x19990, x19999);
  nand n21081(x21081, x19989, x19998);
  nand n21082(x21082, x21081, x21080);
  nand n21083(x21083, x19928, x19937);
  nand n21086(x21086, x21085, x21084);
  nand n21087(x21087, x21086, x21083);
  nand n21089(x21089, x19946, x21088);
  nand n21091(x21091, x21090, x21087);
  nand n21092(x21092, x21091, x21089);
  nand n21094(x21094, x21083, x21089);
  nand n21095(x21095, x19955, x19964);
  nand n21098(x21098, x21097, x21096);
  nand n21099(x21099, x21098, x21095);
  nand n21101(x21101, x19973, x21100);
  nand n21103(x21103, x21102, x21099);
  nand n21104(x21104, x21103, x21101);
  nand n21106(x21106, x21095, x21101);
  nand n21107(x21107, x19982, x19991);
  nand n21110(x21110, x21109, x21108);
  nand n21111(x21111, x21110, x21107);
  nand n21113(x21113, x20000, x21112);
  nand n21115(x21115, x21114, x21111);
  nand n21116(x21116, x21115, x21113);
  nand n21118(x21118, x21107, x21113);
  nand n21119(x21119, x20016, x20025);
  nand n21120(x21120, x20015, x20024);
  nand n21121(x21121, x21120, x21119);
  nand n21123(x21123, x20034, x21122);
  nand n21124(x21124, x20033, x21121);
  nand n21125(x21125, x21124, x21123);
  nand n21127(x21127, x21119, x21123);
  nand n21128(x21128, x20043, x20052);
  nand n21129(x21129, x20042, x20051);
  nand n21130(x21130, x21129, x21128);
  nand n21132(x21132, x20061, x21131);
  nand n21133(x21133, x20060, x21130);
  nand n21134(x21134, x21133, x21132);
  nand n21136(x21136, x21128, x21132);
  nand n21137(x21137, x20070, x20079);
  nand n21138(x21138, x20069, x20078);
  nand n21139(x21139, x21138, x21137);
  nand n21141(x21141, x83591, x21140);
  nand n21142(x21142, x18705, x21139);
  nand n21143(x21143, x21142, x21141);
  nand n21145(x21145, x21137, x21141);
  nand n21146(x21146, x20008, x20017);
  nand n21149(x21149, x21148, x21147);
  nand n21150(x21150, x21149, x21146);
  nand n21152(x21152, x20026, x21151);
  nand n21154(x21154, x21153, x21150);
  nand n21155(x21155, x21154, x21152);
  nand n21157(x21157, x21146, x21152);
  nand n21158(x21158, x20035, x20044);
  nand n21161(x21161, x21160, x21159);
  nand n21162(x21162, x21161, x21158);
  nand n21164(x21164, x20053, x21163);
  nand n21166(x21166, x21165, x21162);
  nand n21167(x21167, x21166, x21164);
  nand n21169(x21169, x21158, x21164);
  nand n21170(x21170, x20062, x20071);
  nand n21173(x21173, x21172, x21171);
  nand n21174(x21174, x21173, x21170);
  nand n21176(x21176, x20080, x21175);
  nand n21178(x21178, x21177, x21174);
  nand n21179(x21179, x21178, x21176);
  nand n21181(x21181, x21170, x21176);
  nand n21182(x21182, x20096, x20105);
  nand n21183(x21183, x20095, x20104);
  nand n21184(x21184, x21183, x21182);
  nand n21186(x21186, x20114, x21185);
  nand n21187(x21187, x20113, x21184);
  nand n21188(x21188, x21187, x21186);
  nand n21190(x21190, x21182, x21186);
  nand n21191(x21191, x20123, x20132);
  nand n21192(x21192, x20122, x20131);
  nand n21193(x21193, x21192, x21191);
  nand n21195(x21195, x20141, x21194);
  nand n21196(x21196, x20140, x21193);
  nand n21197(x21197, x21196, x21195);
  nand n21199(x21199, x21191, x21195);
  nand n21200(x21200, x20150, x20159);
  nand n21201(x21201, x20149, x20158);
  nand n21202(x21202, x21201, x21200);
  nand n21204(x21204, x83592, x21203);
  nand n21205(x21205, x20163, x21202);
  nand n21206(x21206, x21205, x21204);
  nand n21208(x21208, x21200, x21204);
  nand n21209(x21209, x20088, x20097);
  nand n21212(x21212, x21211, x21210);
  nand n21213(x21213, x21212, x21209);
  nand n21215(x21215, x20106, x21214);
  nand n21217(x21217, x21216, x21213);
  nand n21218(x21218, x21217, x21215);
  nand n21220(x21220, x21209, x21215);
  nand n21221(x21221, x20115, x20124);
  nand n21224(x21224, x21223, x21222);
  nand n21225(x21225, x21224, x21221);
  nand n21227(x21227, x20133, x21226);
  nand n21229(x21229, x21228, x21225);
  nand n21230(x21230, x21229, x21227);
  nand n21232(x21232, x21221, x21227);
  nand n21233(x21233, x20142, x20151);
  nand n21236(x21236, x21235, x21234);
  nand n21237(x21237, x21236, x21233);
  nand n21239(x21239, x20160, x21238);
  nand n21241(x21241, x21240, x21237);
  nand n21242(x21242, x21241, x21239);
  nand n21244(x21244, x21233, x21239);
  nand n21245(x21245, x20171, x83635);
  nand n21246(x21246, x20170, x20161);
  nand n21247(x21247, x21246, x21245);
  nand n21249(x21249, x20180, x20189);
  nand n21250(x21250, x20179, x20188);
  nand n21251(x21251, x21250, x21249);
  nand n21253(x21253, x20198, x21252);
  nand n21254(x21254, x20197, x21251);
  nand n21255(x21255, x21254, x21253);
  nand n21257(x21257, x21249, x21253);
  nand n21258(x21258, x20207, x20216);
  nand n21259(x21259, x20206, x20215);
  nand n21260(x21260, x21259, x21258);
  nand n21262(x21262, x20225, x21261);
  nand n21263(x21263, x20224, x21260);
  nand n21264(x21264, x21263, x21262);
  nand n21266(x21266, x21258, x21262);
  nand n21267(x21267, x20234, x20243);
  nand n21268(x21268, x20233, x20242);
  nand n21269(x21269, x21268, x21267);
  nand n21271(x21271, x20252, x21270);
  nand n21272(x21272, x20251, x21269);
  nand n21273(x21273, x21272, x21271);
  nand n21275(x21275, x21267, x21271);
  nand n21276(x21276, x20172, x20181);
  nand n21279(x21279, x21278, x21277);
  nand n21280(x21280, x21279, x21276);
  nand n21282(x21282, x20190, x21281);
  nand n21284(x21284, x21283, x21280);
  nand n21285(x21285, x21284, x21282);
  nand n21287(x21287, x21276, x21282);
  nand n21288(x21288, x20199, x20208);
  nand n21291(x21291, x21290, x21289);
  nand n21292(x21292, x21291, x21288);
  nand n21294(x21294, x20217, x21293);
  nand n21296(x21296, x21295, x21292);
  nand n21297(x21297, x21296, x21294);
  nand n21299(x21299, x21288, x21294);
  nand n21300(x21300, x20226, x20235);
  nand n21303(x21303, x21302, x21301);
  nand n21304(x21304, x21303, x21300);
  nand n21306(x21306, x20244, x21305);
  nand n21308(x21308, x21307, x21304);
  nand n21309(x21309, x21308, x21306);
  nand n21311(x21311, x21300, x21306);
  nand n21313(x21313, x20261, x20253);
  nand n21314(x21314, x20260, x21312);
  nand n21315(x21315, x21314, x21313);
  nand n21317(x21317, x20270, x20279);
  nand n21318(x21318, x20269, x20278);
  nand n21319(x21319, x21318, x21317);
  nand n21321(x21321, x20288, x21320);
  nand n21322(x21322, x20287, x21319);
  nand n21323(x21323, x21322, x21321);
  nand n21325(x21325, x21317, x21321);
  nand n21326(x21326, x20297, x20306);
  nand n21327(x21327, x20296, x20305);
  nand n21328(x21328, x21327, x21326);
  nand n21330(x21330, x20315, x21329);
  nand n21331(x21331, x20314, x21328);
  nand n21332(x21332, x21331, x21330);
  nand n21334(x21334, x21326, x21330);
  nand n21335(x21335, x20324, x20333);
  nand n21336(x21336, x20323, x20332);
  nand n21337(x21337, x21336, x21335);
  nand n21339(x21339, x20342, x21338);
  nand n21340(x21340, x20341, x21337);
  nand n21341(x21341, x21340, x21339);
  nand n21343(x21343, x21335, x21339);
  nand n21344(x21344, x20262, x20271);
  nand n21347(x21347, x21346, x21345);
  nand n21348(x21348, x21347, x21344);
  nand n21350(x21350, x20280, x21349);
  nand n21352(x21352, x21351, x21348);
  nand n21353(x21353, x21352, x21350);
  nand n21355(x21355, x20289, x20298);
  nand n21358(x21358, x21357, x21356);
  nand n21359(x21359, x21358, x21355);
  nand n21361(x21361, x20307, x21360);
  nand n21363(x21363, x21362, x21359);
  nand n21364(x21364, x21363, x21361);
  nand n21366(x21366, x20316, x20325);
  nand n21369(x21369, x21368, x21367);
  nand n21370(x21370, x21369, x21366);
  nand n21372(x21372, x20334, x21371);
  nand n21374(x21374, x21373, x21370);
  nand n21375(x21375, x21374, x21372);
  nand n21378(x21378, x20351, x20343);
  nand n21379(x21379, x20350, x21377);
  nand n21380(x21380, x21379, x21378);
  nand n21382(x21382, x20359, x20367);
  nand n21383(x21383, x20358, x20366);
  nand n21384(x21384, x21383, x21382);
  nand n21386(x21386, x20375, x21385);
  nand n21387(x21387, x20374, x21384);
  nand n21388(x21388, x21387, x21386);
  nand n21390(x21390, x20383, x20391);
  nand n21391(x21391, x20382, x20390);
  nand n21392(x21392, x21391, x21390);
  nand n21394(x21394, x20399, x21393);
  nand n21395(x21395, x20398, x21392);
  nand n21396(x21396, x21395, x21394);
  nand n21398(x21398, x20407, x20415);
  nand n21399(x21399, x20406, x20414);
  nand n21400(x21400, x21399, x21398);
  nand n21402(x21402, x20423, x21401);
  nand n21403(x21403, x20422, x21400);
  nand n21404(x21404, x21403, x21402);
  nand n21406(x21406, x83594, x83640);
  nand n21407(x21407, x17921, x18966);
  nand n21408(x21408, x21407, x21406);
  nand n21410(x21410, x83595, x83641);
  nand n21411(x21411, x18978, x18974);
  nand n21412(x21412, x21411, x21410);
  nand n21414(x21414, x83596, x83642);
  nand n21415(x21415, x18993, x18985);
  nand n21416(x21416, x21415, x21414);
  nand n21418(x21418, x83597, x83644);
  nand n21419(x21419, x20441, x19001);
  nand n21420(x21420, x21419, x21418);
  nand n21422(x21422, x83598, x83648);
  nand n21423(x21423, x20449, x19018);
  nand n21424(x21424, x21423, x21422);
  nand n21426(x21426, x83599, x83652);
  nand n21427(x21427, x20462, x19038);
  nand n21428(x21428, x21427, x21426);
  nand n21431(x21431, x20481, x83655);
  nand n21432(x21432, x20480, x19064);
  nand n21433(x21433, x21432, x21431);
  nand n21437(x21437, x20501, x83657);
  nand n21438(x21438, x20500, x19090);
  nand n21439(x21439, x21438, x21437);
  nand n21443(x21443, x83600, x83658);
  nand n21444(x21444, x19110, x20512);
  nand n21445(x21445, x21444, x21443);
  nand n21447(x21447, x20521, x83659);
  nand n21448(x21448, x20520, x19119);
  nand n21449(x21449, x21448, x21447);
  nand n21453(x21453, x19147, x83660);
  nand n21454(x21454, x20534, x20532);
  nand n21455(x21455, x21454, x21453);
  nand n21457(x21457, x20542, x83661);
  nand n21458(x21458, x20541, x19154);
  nand n21459(x21459, x21458, x21457);
  nand n21463(x21463, x19182, x83663);
  nand n21464(x21464, x20555, x20553);
  nand n21465(x21465, x21464, x21463);
  nand n21467(x21467, x20563, x83664);
  nand n21468(x21468, x20562, x19189);
  nand n21469(x21469, x21468, x21467);
  nand n21473(x21473, x83601, x83666);
  nand n21474(x21474, x20579, x20574);
  nand n21475(x21475, x21474, x21473);
  nand n21477(x21477, x20587, x83667);
  nand n21478(x21478, x20586, x19227);
  nand n21479(x21479, x21478, x21477);
  nand n21481(x21481, x20575, x83602);
  nand n21483(x21483, x21482, x20576);
  nand n21484(x21484, x21483, x21481);
  nand n21486(x21486, x83603, x83670);
  nand n21487(x21487, x20604, x20598);
  nand n21488(x21488, x21487, x21486);
  nand n21490(x21490, x20612, x83672);
  nand n21491(x21491, x20611, x19270);
  nand n21492(x21492, x21491, x21490);
  nand n21494(x21494, x20599, x83604);
  nand n21496(x21496, x21495, x20600);
  nand n21497(x21497, x21496, x21494);
  nand n21499(x21499, x83605, x20613);
  nand n21500(x21500, x20614, x21498);
  nand n21501(x21501, x21500, x21499);
  nand n21503(x21503, x83606, x83677);
  nand n21504(x21504, x20632, x20626);
  nand n21505(x21505, x21504, x21503);
  nand n21507(x21507, x20640, x83679);
  nand n21508(x21508, x20639, x19314);
  nand n21509(x21509, x21508, x21507);
  nand n21511(x21511, x20627, x83607);
  nand n21513(x21513, x21512, x20628);
  nand n21514(x21514, x21513, x21511);
  nand n21516(x21516, x83608, x20641);
  nand n21517(x21517, x20642, x21515);
  nand n21518(x21518, x21517, x21516);
  nand n21520(x21520, x20665, x83684);
  nand n21521(x21521, x20664, x20654);
  nand n21522(x21522, x21521, x21520);
  nand n21524(x21524, x20674, x83686);
  nand n21525(x21525, x20673, x19361);
  nand n21526(x21526, x21525, x21524);
  nand n21528(x21528, x20655, x20666);
  nand n21531(x21531, x21530, x21529);
  nand n21532(x21532, x21531, x21528);
  nand n21534(x21534, x83609, x20675);
  nand n21535(x21535, x20676, x21533);
  nand n21536(x21536, x21535, x21534);
  nand n21538(x21538, x20700, x83691);
  nand n21539(x21539, x20699, x20688);
  nand n21540(x21540, x21539, x21538);
  nand n21542(x21542, x20709, x83693);
  nand n21543(x21543, x20708, x19414);
  nand n21544(x21544, x21543, x21542);
  nand n21546(x21546, x20689, x20701);
  nand n21549(x21549, x21548, x21547);
  nand n21550(x21550, x21549, x21546);
  nand n21552(x21552, x20718, x20710);
  nand n21554(x21554, x21553, x21551);
  nand n21555(x21555, x21554, x21552);
  nand n21557(x21557, x20740, x83698);
  nand n21558(x21558, x20739, x20728);
  nand n21559(x21559, x21558, x21557);
  nand n21561(x21561, x20749, x83700);
  nand n21562(x21562, x20748, x19467);
  nand n21563(x21563, x21562, x21561);
  nand n21565(x21565, x20729, x20741);
  nand n21568(x21568, x21567, x21566);
  nand n21569(x21569, x21568, x21565);
  nand n21571(x21571, x20758, x20750);
  nand n21573(x21573, x21572, x21570);
  nand n21574(x21574, x21573, x21571);
  nand n21576(x21576, x20780, x83705);
  nand n21577(x21577, x20779, x20768);
  nand n21578(x21578, x21577, x21576);
  nand n21580(x21580, x83610, x83611);
  nand n21581(x21581, x19514, x19523);
  nand n21582(x21582, x21581, x21580);
  nand n21584(x21584, x20789, x21583);
  nand n21585(x21585, x20788, x21582);
  nand n21586(x21586, x21585, x21584);
  nand n21588(x21588, x21580, x21584);
  nand n21589(x21589, x20769, x20781);
  nand n21592(x21592, x21591, x21590);
  nand n21593(x21593, x21592, x21589);
  nand n21595(x21595, x20798, x20790);
  nand n21597(x21597, x21596, x21594);
  nand n21598(x21598, x21597, x21595);
  nand n21600(x21600, x20820, x83711);
  nand n21601(x21601, x20819, x20808);
  nand n21602(x21602, x21601, x21600);
  nand n21604(x21604, x19578, x83612);
  nand n21605(x21605, x20822, x19585);
  nand n21606(x21606, x21605, x21604);
  nand n21608(x21608, x20830, x21607);
  nand n21609(x21609, x20829, x21606);
  nand n21610(x21610, x21609, x21608);
  nand n21612(x21612, x21604, x21608);
  nand n21613(x21613, x20839, x83613);
  nand n21614(x21614, x20838, x18401);
  nand n21615(x21615, x21614, x21613);
  nand n21616(x21616, x20809, x20821);
  nand n21619(x21619, x21618, x21617);
  nand n21620(x21620, x21619, x21616);
  nand n21622(x21622, x20840, x20831);
  nand n21624(x21624, x21623, x21621);
  nand n21625(x21625, x21624, x21622);
  nand n21627(x21627, x20862, x83718);
  nand n21628(x21628, x20861, x20850);
  nand n21629(x21629, x21628, x21627);
  nand n21631(x21631, x19640, x83614);
  nand n21632(x21632, x20864, x19647);
  nand n21633(x21633, x21632, x21631);
  nand n21635(x21635, x20872, x21634);
  nand n21636(x21636, x20871, x21633);
  nand n21637(x21637, x21636, x21635);
  nand n21639(x21639, x21631, x21635);
  nand n21640(x21640, x20881, x83615);
  nand n21641(x21641, x20880, x19705);
  nand n21642(x21642, x21641, x21640);
  nand n21643(x21643, x20851, x20863);
  nand n21646(x21646, x21645, x21644);
  nand n21647(x21647, x21646, x21643);
  nand n21649(x21649, x20882, x20873);
  nand n21651(x21651, x21650, x21648);
  nand n21652(x21652, x21651, x21649);
  nand n21654(x21654, x20904, x83725);
  nand n21655(x21655, x20903, x20892);
  nand n21656(x21656, x21655, x21654);
  nand n21658(x21658, x83616, x83618);
  nand n21659(x21659, x20909, x19712);
  nand n21660(x21660, x21659, x21658);
  nand n21662(x21662, x20917, x21661);
  nand n21663(x21663, x20916, x21660);
  nand n21664(x21664, x21663, x21662);
  nand n21666(x21666, x21658, x21662);
  nand n21667(x21667, x20926, x83619);
  nand n21668(x21668, x20925, x19774);
  nand n21669(x21669, x21668, x21667);
  nand n21670(x21670, x20893, x20905);
  nand n21673(x21673, x21672, x21671);
  nand n21674(x21674, x21673, x21670);
  nand n21676(x21676, x83617, x21675);
  nand n21677(x21677, x20906, x21674);
  nand n21678(x21678, x21677, x21676);
  nand n21680(x21680, x21670, x21676);
  nand n21682(x21682, x20927, x20918);
  nand n21684(x21684, x21683, x21681);
  nand n21685(x21685, x21684, x21682);
  nand n21687(x21687, x20949, x83730);
  nand n21688(x21688, x20948, x20937);
  nand n21689(x21689, x21688, x21687);
  nand n21691(x21691, x83620, x83622);
  nand n21692(x21692, x20955, x19782);
  nand n21693(x21693, x21692, x21691);
  nand n21695(x21695, x20963, x21694);
  nand n21696(x21696, x20962, x21693);
  nand n21697(x21697, x21696, x21695);
  nand n21699(x21699, x21691, x21695);
  nand n21700(x21700, x20972, x83623);
  nand n21701(x21701, x20971, x20976);
  nand n21702(x21702, x21701, x21700);
  nand n21703(x21703, x20938, x20950);
  nand n21706(x21706, x21705, x21704);
  nand n21707(x21707, x21706, x21703);
  nand n21709(x21709, x83621, x21708);
  nand n21710(x21710, x20951, x21707);
  nand n21711(x21711, x21710, x21709);
  nand n21713(x21713, x21703, x21709);
  nand n21715(x21715, x20973, x20964);
  nand n21717(x21717, x21716, x21714);
  nand n21718(x21718, x21717, x21715);
  nand n21720(x21720, x83624, x20987);
  nand n21721(x21721, x20974, x20986);
  nand n21722(x21722, x21721, x21720);
  nand n21724(x21724, x20999, x21723);
  nand n21725(x21725, x20998, x21722);
  nand n21726(x21726, x21725, x21724);
  nand n21728(x21728, x21720, x21724);
  nand n21729(x21729, x83625, x83627);
  nand n21730(x21730, x21005, x19853);
  nand n21731(x21731, x21730, x21729);
  nand n21733(x21733, x21013, x21732);
  nand n21734(x21734, x21012, x21731);
  nand n21735(x21735, x21734, x21733);
  nand n21737(x21737, x21729, x21733);
  nand n21738(x21738, x21022, x83628);
  nand n21739(x21739, x21021, x21026);
  nand n21740(x21740, x21739, x21738);
  nand n21741(x21741, x20988, x21000);
  nand n21744(x21744, x21743, x21742);
  nand n21745(x21745, x21744, x21741);
  nand n21747(x21747, x83626, x21746);
  nand n21748(x21748, x21001, x21745);
  nand n21749(x21749, x21748, x21747);
  nand n21751(x21751, x21741, x21747);
  nand n21753(x21753, x21023, x21014);
  nand n21755(x21755, x21754, x21752);
  nand n21756(x21756, x21755, x21753);
  nand n21758(x21758, x83629, x21037);
  nand n21759(x21759, x21024, x21036);
  nand n21760(x21760, x21759, x21758);
  nand n21762(x21762, x21049, x21761);
  nand n21763(x21763, x21048, x21760);
  nand n21764(x21764, x21763, x21762);
  nand n21766(x21766, x21758, x21762);
  nand n21767(x21767, x21060, x83630);
  nand n21768(x21768, x21059, x19927);
  nand n21769(x21769, x21768, x21767);
  nand n21771(x21771, x21069, x21770);
  nand n21772(x21772, x21068, x21769);
  nand n21773(x21773, x21772, x21771);
  nand n21775(x21775, x21767, x21771);
  nand n21776(x21776, x21078, x83631);
  nand n21777(x21777, x21077, x21082);
  nand n21778(x21778, x21777, x21776);
  nand n21779(x21779, x21038, x21050);
  nand n21782(x21782, x21781, x21780);
  nand n21783(x21783, x21782, x21779);
  nand n21785(x21785, x21061, x21784);
  nand n21787(x21787, x21786, x21783);
  nand n21788(x21788, x21787, x21785);
  nand n21790(x21790, x21779, x21785);
  nand n21792(x21792, x21079, x21070);
  nand n21794(x21794, x21793, x21791);
  nand n21795(x21795, x21794, x21792);
  nand n21797(x21797, x83632, x21093);
  nand n21798(x21798, x21080, x21092);
  nand n21799(x21799, x21798, x21797);
  nand n21801(x21801, x21105, x21800);
  nand n21802(x21802, x21104, x21799);
  nand n21803(x21803, x21802, x21801);
  nand n21805(x21805, x21797, x21801);
  nand n21806(x21806, x21117, x83633);
  nand n21807(x21807, x21116, x20007);
  nand n21808(x21808, x21807, x21806);
  nand n21810(x21810, x21126, x21809);
  nand n21811(x21811, x21125, x21808);
  nand n21812(x21812, x21811, x21810);
  nand n21814(x21814, x21806, x21810);
  nand n21815(x21815, x21135, x21144);
  nand n21816(x21816, x21134, x21143);
  nand n21817(x21817, x21816, x21815);
  nand n21818(x21818, x21094, x21106);
  nand n21821(x21821, x21820, x21819);
  nand n21822(x21822, x21821, x21818);
  nand n21824(x21824, x21118, x21823);
  nand n21826(x21826, x21825, x21822);
  nand n21827(x21827, x21826, x21824);
  nand n21829(x21829, x21818, x21824);
  nand n21831(x21831, x21136, x21127);
  nand n21833(x21833, x21832, x21830);
  nand n21834(x21834, x21833, x21831);
  nand n21836(x21836, x21145, x21156);
  nand n21838(x21838, x21837, x21155);
  nand n21839(x21839, x21838, x21836);
  nand n21841(x21841, x21168, x21840);
  nand n21842(x21842, x21167, x21839);
  nand n21843(x21843, x21842, x21841);
  nand n21845(x21845, x21836, x21841);
  nand n21846(x21846, x21180, x83634);
  nand n21847(x21847, x21179, x20087);
  nand n21848(x21848, x21847, x21846);
  nand n21850(x21850, x21189, x21849);
  nand n21851(x21851, x21188, x21848);
  nand n21852(x21852, x21851, x21850);
  nand n21854(x21854, x21846, x21850);
  nand n21855(x21855, x21198, x21207);
  nand n21856(x21856, x21197, x21206);
  nand n21857(x21857, x21856, x21855);
  nand n21858(x21858, x21157, x21169);
  nand n21861(x21861, x21860, x21859);
  nand n21862(x21862, x21861, x21858);
  nand n21864(x21864, x21181, x21863);
  nand n21866(x21866, x21865, x21862);
  nand n21867(x21867, x21866, x21864);
  nand n21869(x21869, x21858, x21864);
  nand n21871(x21871, x21199, x21190);
  nand n21873(x21873, x21872, x21870);
  nand n21874(x21874, x21873, x21871);
  nand n21876(x21876, x21208, x21219);
  nand n21878(x21878, x21877, x21218);
  nand n21879(x21879, x21878, x21876);
  nand n21881(x21881, x21231, x21880);
  nand n21882(x21882, x21230, x21879);
  nand n21883(x21883, x21882, x21881);
  nand n21885(x21885, x21876, x21881);
  nand n21886(x21886, x21243, x21248);
  nand n21887(x21887, x21242, x21247);
  nand n21888(x21888, x21887, x21886);
  nand n21890(x21890, x21256, x21889);
  nand n21891(x21891, x21255, x21888);
  nand n21892(x21892, x21891, x21890);
  nand n21894(x21894, x21886, x21890);
  nand n21895(x21895, x21265, x21274);
  nand n21896(x21896, x21264, x21273);
  nand n21897(x21897, x21896, x21895);
  nand n21898(x21898, x21220, x21232);
  nand n21901(x21901, x21900, x21899);
  nand n21902(x21902, x21901, x21898);
  nand n21904(x21904, x21244, x21903);
  nand n21906(x21906, x21905, x21902);
  nand n21907(x21907, x21906, x21904);
  nand n21909(x21909, x21898, x21904);
  nand n21910(x21910, x83636, x21257);
  nand n21912(x21912, x21245, x21911);
  nand n21913(x21913, x21912, x21910);
  nand n21915(x21915, x21266, x21914);
  nand n21917(x21917, x21916, x21913);
  nand n21918(x21918, x21917, x21915);
  nand n21920(x21920, x21910, x21915);
  nand n21921(x21921, x21275, x21286);
  nand n21923(x21923, x21922, x21285);
  nand n21924(x21924, x21923, x21921);
  nand n21926(x21926, x21298, x21925);
  nand n21927(x21927, x21297, x21924);
  nand n21928(x21928, x21927, x21926);
  nand n21930(x21930, x21921, x21926);
  nand n21931(x21931, x21310, x21316);
  nand n21932(x21932, x21309, x21315);
  nand n21933(x21933, x21932, x21931);
  nand n21935(x21935, x21324, x21934);
  nand n21936(x21936, x21323, x21933);
  nand n21937(x21937, x21936, x21935);
  nand n21939(x21939, x21931, x21935);
  nand n21940(x21940, x21333, x21342);
  nand n21941(x21941, x21332, x21341);
  nand n21942(x21942, x21941, x21940);
  nand n21944(x21944, x83593, x21943);
  nand n21945(x21945, x18884, x21942);
  nand n21946(x21946, x21945, x21944);
  nand n21948(x21948, x21940, x21944);
  nand n21949(x21949, x21287, x21299);
  nand n21952(x21952, x21951, x21950);
  nand n21953(x21953, x21952, x21949);
  nand n21955(x21955, x21311, x21954);
  nand n21957(x21957, x21956, x21953);
  nand n21958(x21958, x21957, x21955);
  nand n21960(x21960, x83637, x21325);
  nand n21962(x21962, x21313, x21961);
  nand n21963(x21963, x21962, x21960);
  nand n21965(x21965, x21334, x21964);
  nand n21967(x21967, x21966, x21963);
  nand n21968(x21968, x21967, x21965);
  nand n21970(x21970, x21343, x21354);
  nand n21972(x21972, x21971, x21353);
  nand n21973(x21973, x21972, x21970);
  nand n21975(x21975, x21365, x21974);
  nand n21976(x21976, x21364, x21973);
  nand n21977(x21977, x21976, x21975);
  nand n21979(x21979, x21376, x21381);
  nand n21980(x21980, x21375, x21380);
  nand n21981(x21981, x21980, x21979);
  nand n21983(x21983, x21389, x21982);
  nand n21984(x21984, x21388, x21981);
  nand n21985(x21985, x21984, x21983);
  nand n21987(x21987, x21397, x21405);
  nand n21988(x21988, x21396, x21404);
  nand n21989(x21989, x21988, x21987);
  nand n21991(x21991, x20427, x21990);
  nand n21992(x21992, x20426, x21989);
  nand n21993(x21993, x21992, x21991);
  nand n21995(x21995, x83638, x83639);
  nand n21996(x21996, x18949, x18958);
  nand n21997(x21997, x21996, x21995);
  nand n21998(x21998, x21409, x18959);
  nand n21999(x21999, x21408, x20428);
  nand n22000(x22000, x21999, x21998);
  nand n22001(x22001, x21413, x18967);
  nand n22002(x22002, x21412, x20429);
  nand n22003(x22003, x22002, x22001);
  nand n22005(x22005, x21417, x83749);
  nand n22006(x22006, x21416, x20433);
  nand n22007(x22007, x22006, x22005);
  nand n22009(x22009, x83643, x83750);
  nand n22010(x22010, x20430, x21414);
  nand n22011(x22011, x22010, x22009);
  nand n22012(x22012, x21421, x83751);
  nand n22013(x22013, x21420, x20438);
  nand n22014(x22014, x22013, x22012);
  nand n22016(x22016, x83645, x83753);
  nand n22017(x22017, x20434, x21418);
  nand n22018(x22018, x22017, x22016);
  nand n22019(x22019, x83646, x83647);
  nand n22020(x22020, x20439, x20446);
  nand n22021(x22021, x22020, x22019);
  nand n22023(x22023, x21425, x22022);
  nand n22024(x22024, x21424, x22021);
  nand n22025(x22025, x22024, x22023);
  nand n22027(x22027, x22019, x22023);
  nand n22028(x22028, x83649, x83754);
  nand n22029(x22029, x20442, x21422);
  nand n22030(x22030, x22029, x22028);
  nand n22031(x22031, x83650, x83651);
  nand n22032(x22032, x20447, x20458);
  nand n22033(x22033, x22032, x22031);
  nand n22035(x22035, x21429, x22034);
  nand n22036(x22036, x21428, x22033);
  nand n22037(x22037, x22036, x22035);
  nand n22039(x22039, x22031, x22035);
  nand n22040(x22040, x20459, x83755);
  nand n22041(x22041, x21430, x21426);
  nand n22042(x22042, x22041, x22040);
  nand n22043(x22043, x83653, x83654);
  nand n22044(x22044, x20460, x20472);
  nand n22045(x22045, x22044, x22043);
  nand n22047(x22047, x21434, x22046);
  nand n22048(x22048, x21433, x22045);
  nand n22049(x22049, x22048, x22047);
  nand n22051(x22051, x22043, x22047);
  nand n22052(x22052, x20473, x83756);
  nand n22053(x22053, x21435, x21431);
  nand n22054(x22054, x22053, x22052);
  nand n22055(x22055, x20482, x83656);
  nand n22056(x22056, x21436, x20492);
  nand n22057(x22057, x22056, x22055);
  nand n22059(x22059, x21440, x22058);
  nand n22060(x22060, x21439, x22057);
  nand n22061(x22061, x22060, x22059);
  nand n22063(x22063, x22055, x22059);
  nand n22064(x22064, x20493, x83757);
  nand n22065(x22065, x21441, x21437);
  nand n22066(x22066, x22065, x22064);
  nand n22067(x22067, x20502, x21446);
  nand n22068(x22068, x21442, x21445);
  nand n22069(x22069, x22068, x22067);
  nand n22071(x22071, x21450, x22070);
  nand n22072(x22072, x21449, x22069);
  nand n22073(x22073, x22072, x22071);
  nand n22075(x22075, x22067, x22071);
  nand n22076(x22076, x20513, x83759);
  nand n22077(x22077, x21451, x21447);
  nand n22078(x22078, x22077, x22076);
  nand n22080(x22080, x20522, x21456);
  nand n22081(x22081, x21452, x21455);
  nand n22082(x22082, x22081, x22080);
  nand n22084(x22084, x21460, x22083);
  nand n22085(x22085, x21459, x22082);
  nand n22086(x22086, x22085, x22084);
  nand n22088(x22088, x22080, x22084);
  nand n22089(x22089, x20533, x83761);
  nand n22090(x22090, x21461, x21457);
  nand n22091(x22091, x22090, x22089);
  nand n22093(x22093, x20543, x21466);
  nand n22094(x22094, x21462, x21465);
  nand n22095(x22095, x22094, x22093);
  nand n22097(x22097, x21470, x22096);
  nand n22098(x22098, x21469, x22095);
  nand n22099(x22099, x22098, x22097);
  nand n22101(x22101, x22093, x22097);
  nand n22102(x22102, x20554, x83763);
  nand n22103(x22103, x21471, x21467);
  nand n22104(x22104, x22103, x22102);
  nand n22106(x22106, x20564, x21476);
  nand n22107(x22107, x21472, x21475);
  nand n22108(x22108, x22107, x22106);
  nand n22110(x22110, x21480, x22109);
  nand n22111(x22111, x21479, x22108);
  nand n22112(x22112, x22111, x22110);
  nand n22114(x22114, x22106, x22110);
  nand n22115(x22115, x83669, x83765);
  nand n22116(x22116, x21484, x21477);
  nand n22117(x22117, x22116, x22115);
  nand n22119(x22119, x20588, x21489);
  nand n22120(x22120, x21485, x21488);
  nand n22121(x22121, x22120, x22119);
  nand n22123(x22123, x21493, x22122);
  nand n22124(x22124, x21492, x22121);
  nand n22125(x22125, x22124, x22123);
  nand n22127(x22127, x22119, x22123);
  nand n22128(x22128, x83671, x83766);
  nand n22129(x22129, x21486, x21481);
  nand n22130(x22130, x22129, x22128);
  nand n22132(x22132, x83674, x83768);
  nand n22133(x22133, x21497, x21490);
  nand n22134(x22134, x22133, x22132);
  nand n22136(x22136, x21502, x21506);
  nand n22137(x22137, x21501, x21505);
  nand n22138(x22138, x22137, x22136);
  nand n22140(x22140, x21510, x22139);
  nand n22141(x22141, x21509, x22138);
  nand n22142(x22142, x22141, x22140);
  nand n22144(x22144, x22136, x22140);
  nand n22145(x22145, x83675, x83676);
  nand n22146(x22146, x21494, x21499);
  nand n22147(x22147, x22146, x22145);
  nand n22149(x22149, x83678, x22148);
  nand n22150(x22150, x21503, x22147);
  nand n22151(x22151, x22150, x22149);
  nand n22153(x22153, x22145, x22149);
  nand n22154(x22154, x83681, x83770);
  nand n22155(x22155, x21514, x21507);
  nand n22156(x22156, x22155, x22154);
  nand n22158(x22158, x21519, x21523);
  nand n22159(x22159, x21518, x21522);
  nand n22160(x22160, x22159, x22158);
  nand n22162(x22162, x21527, x22161);
  nand n22163(x22163, x21526, x22160);
  nand n22164(x22164, x22163, x22162);
  nand n22166(x22166, x22158, x22162);
  nand n22167(x22167, x83682, x83683);
  nand n22168(x22168, x21511, x21516);
  nand n22169(x22169, x22168, x22167);
  nand n22171(x22171, x83685, x22170);
  nand n22172(x22172, x21520, x22169);
  nand n22173(x22173, x22172, x22171);
  nand n22175(x22175, x22167, x22171);
  nand n22176(x22176, x83688, x83772);
  nand n22177(x22177, x21532, x21524);
  nand n22178(x22178, x22177, x22176);
  nand n22180(x22180, x21537, x21541);
  nand n22181(x22181, x21536, x21540);
  nand n22182(x22182, x22181, x22180);
  nand n22184(x22184, x21545, x22183);
  nand n22185(x22185, x21544, x22182);
  nand n22186(x22186, x22185, x22184);
  nand n22188(x22188, x22180, x22184);
  nand n22189(x22189, x83689, x83690);
  nand n22190(x22190, x21528, x21534);
  nand n22191(x22191, x22190, x22189);
  nand n22193(x22193, x83692, x22192);
  nand n22194(x22194, x21538, x22191);
  nand n22195(x22195, x22194, x22193);
  nand n22197(x22197, x22189, x22193);
  nand n22198(x22198, x83695, x83774);
  nand n22199(x22199, x21550, x21542);
  nand n22200(x22200, x22199, x22198);
  nand n22202(x22202, x21556, x21560);
  nand n22203(x22203, x21555, x21559);
  nand n22204(x22204, x22203, x22202);
  nand n22206(x22206, x21564, x22205);
  nand n22207(x22207, x21563, x22204);
  nand n22208(x22208, x22207, x22206);
  nand n22210(x22210, x22202, x22206);
  nand n22211(x22211, x83696, x83697);
  nand n22212(x22212, x21546, x21552);
  nand n22213(x22213, x22212, x22211);
  nand n22215(x22215, x83699, x22214);
  nand n22216(x22216, x21557, x22213);
  nand n22217(x22217, x22216, x22215);
  nand n22219(x22219, x22211, x22215);
  nand n22220(x22220, x83702, x83776);
  nand n22221(x22221, x21569, x21561);
  nand n22222(x22222, x22221, x22220);
  nand n22224(x22224, x21575, x21579);
  nand n22225(x22225, x21574, x21578);
  nand n22226(x22226, x22225, x22224);
  nand n22228(x22228, x21587, x22227);
  nand n22229(x22229, x21586, x22226);
  nand n22230(x22230, x22229, x22228);
  nand n22232(x22232, x22224, x22228);
  nand n22233(x22233, x83703, x83704);
  nand n22234(x22234, x21565, x21571);
  nand n22235(x22235, x22234, x22233);
  nand n22237(x22237, x83706, x22236);
  nand n22238(x22238, x21576, x22235);
  nand n22239(x22239, x22238, x22237);
  nand n22241(x22241, x22233, x22237);
  nand n22243(x22243, x83708, x21588);
  nand n22244(x22244, x21593, x22242);
  nand n22245(x22245, x22244, x22243);
  nand n22247(x22247, x21599, x21603);
  nand n22248(x22248, x21598, x21602);
  nand n22249(x22249, x22248, x22247);
  nand n22251(x22251, x21611, x22250);
  nand n22252(x22252, x21610, x22249);
  nand n22253(x22253, x22252, x22251);
  nand n22255(x22255, x22247, x22251);
  nand n22256(x22256, x83709, x83710);
  nand n22257(x22257, x21589, x21595);
  nand n22258(x22258, x22257, x22256);
  nand n22260(x22260, x83712, x22259);
  nand n22261(x22261, x21600, x22258);
  nand n22262(x22262, x22261, x22260);
  nand n22264(x22264, x22256, x22260);
  nand n22265(x22265, x21612, x83714);
  nand n22267(x22267, x22266, x21613);
  nand n22268(x22268, x22267, x22265);
  nand n22270(x22270, x83715, x22269);
  nand n22271(x22271, x21620, x22268);
  nand n22272(x22272, x22271, x22270);
  nand n22274(x22274, x22265, x22270);
  nand n22275(x22275, x21626, x21630);
  nand n22276(x22276, x21625, x21629);
  nand n22277(x22277, x22276, x22275);
  nand n22279(x22279, x21638, x22278);
  nand n22280(x22280, x21637, x22277);
  nand n22281(x22281, x22280, x22279);
  nand n22283(x22283, x22275, x22279);
  nand n22284(x22284, x83716, x83717);
  nand n22285(x22285, x21616, x21622);
  nand n22286(x22286, x22285, x22284);
  nand n22288(x22288, x83719, x22287);
  nand n22289(x22289, x21627, x22286);
  nand n22290(x22290, x22289, x22288);
  nand n22292(x22292, x22284, x22288);
  nand n22293(x22293, x21639, x83721);
  nand n22295(x22295, x22294, x21640);
  nand n22296(x22296, x22295, x22293);
  nand n22298(x22298, x83722, x22297);
  nand n22299(x22299, x21647, x22296);
  nand n22300(x22300, x22299, x22298);
  nand n22302(x22302, x22293, x22298);
  nand n22303(x22303, x21653, x21657);
  nand n22304(x22304, x21652, x21656);
  nand n22305(x22305, x22304, x22303);
  nand n22307(x22307, x21665, x22306);
  nand n22308(x22308, x21664, x22305);
  nand n22309(x22309, x22308, x22307);
  nand n22311(x22311, x22303, x22307);
  nand n22312(x22312, x83723, x83724);
  nand n22313(x22313, x21643, x21649);
  nand n22314(x22314, x22313, x22312);
  nand n22316(x22316, x83726, x22315);
  nand n22317(x22317, x21654, x22314);
  nand n22318(x22318, x22317, x22316);
  nand n22320(x22320, x22312, x22316);
  nand n22321(x22321, x21666, x83728);
  nand n22323(x22323, x22322, x21667);
  nand n22324(x22324, x22323, x22321);
  nand n22326(x22326, x21679, x22325);
  nand n22327(x22327, x21678, x22324);
  nand n22328(x22328, x22327, x22326);
  nand n22330(x22330, x22321, x22326);
  nand n22331(x22331, x21686, x21690);
  nand n22332(x22332, x21685, x21689);
  nand n22333(x22333, x22332, x22331);
  nand n22335(x22335, x21698, x22334);
  nand n22336(x22336, x21697, x22333);
  nand n22337(x22337, x22336, x22335);
  nand n22339(x22339, x22331, x22335);
  nand n22340(x22340, x21680, x83729);
  nand n22342(x22342, x22341, x21682);
  nand n22343(x22343, x22342, x22340);
  nand n22345(x22345, x83731, x22344);
  nand n22346(x22346, x21687, x22343);
  nand n22347(x22347, x22346, x22345);
  nand n22349(x22349, x22340, x22345);
  nand n22350(x22350, x21699, x83733);
  nand n22352(x22352, x22351, x21700);
  nand n22353(x22353, x22352, x22350);
  nand n22355(x22355, x21712, x22354);
  nand n22356(x22356, x21711, x22353);
  nand n22357(x22357, x22356, x22355);
  nand n22359(x22359, x22350, x22355);
  nand n22360(x22360, x21719, x21727);
  nand n22361(x22361, x21718, x21726);
  nand n22362(x22362, x22361, x22360);
  nand n22364(x22364, x21736, x22363);
  nand n22365(x22365, x21735, x22362);
  nand n22366(x22366, x22365, x22364);
  nand n22368(x22368, x22360, x22364);
  nand n22369(x22369, x21713, x83734);
  nand n22371(x22371, x22370, x21715);
  nand n22372(x22372, x22371, x22369);
  nand n22374(x22374, x21728, x22373);
  nand n22376(x22376, x22375, x22372);
  nand n22377(x22377, x22376, x22374);
  nand n22379(x22379, x22369, x22374);
  nand n22380(x22380, x21737, x83736);
  nand n22382(x22382, x22381, x21738);
  nand n22383(x22383, x22382, x22380);
  nand n22385(x22385, x21750, x22384);
  nand n22386(x22386, x21749, x22383);
  nand n22387(x22387, x22386, x22385);
  nand n22389(x22389, x22380, x22385);
  nand n22390(x22390, x21757, x21765);
  nand n22391(x22391, x21756, x21764);
  nand n22392(x22392, x22391, x22390);
  nand n22394(x22394, x21774, x22393);
  nand n22395(x22395, x21773, x22392);
  nand n22396(x22396, x22395, x22394);
  nand n22398(x22398, x22390, x22394);
  nand n22399(x22399, x21751, x83737);
  nand n22401(x22401, x22400, x21753);
  nand n22402(x22402, x22401, x22399);
  nand n22404(x22404, x21766, x22403);
  nand n22406(x22406, x22405, x22402);
  nand n22407(x22407, x22406, x22404);
  nand n22409(x22409, x22399, x22404);
  nand n22410(x22410, x21775, x83739);
  nand n22412(x22412, x22411, x21776);
  nand n22413(x22413, x22412, x22410);
  nand n22415(x22415, x21789, x22414);
  nand n22416(x22416, x21788, x22413);
  nand n22417(x22417, x22416, x22415);
  nand n22419(x22419, x22410, x22415);
  nand n22420(x22420, x21796, x21804);
  nand n22421(x22421, x21795, x21803);
  nand n22422(x22422, x22421, x22420);
  nand n22424(x22424, x21813, x22423);
  nand n22425(x22425, x21812, x22422);
  nand n22426(x22426, x22425, x22424);
  nand n22428(x22428, x22420, x22424);
  nand n22429(x22429, x21790, x83740);
  nand n22431(x22431, x22430, x21792);
  nand n22432(x22432, x22431, x22429);
  nand n22434(x22434, x21805, x22433);
  nand n22436(x22436, x22435, x22432);
  nand n22437(x22437, x22436, x22434);
  nand n22439(x22439, x22429, x22434);
  nand n22440(x22440, x21814, x83742);
  nand n22442(x22442, x22441, x21815);
  nand n22443(x22443, x22442, x22440);
  nand n22445(x22445, x21828, x22444);
  nand n22446(x22446, x21827, x22443);
  nand n22447(x22447, x22446, x22445);
  nand n22449(x22449, x22440, x22445);
  nand n22450(x22450, x21835, x21844);
  nand n22451(x22451, x21834, x21843);
  nand n22452(x22452, x22451, x22450);
  nand n22454(x22454, x21853, x22453);
  nand n22455(x22455, x21852, x22452);
  nand n22456(x22456, x22455, x22454);
  nand n22458(x22458, x22450, x22454);
  nand n22459(x22459, x21829, x83743);
  nand n22461(x22461, x22460, x21831);
  nand n22462(x22462, x22461, x22459);
  nand n22464(x22464, x21845, x22463);
  nand n22466(x22466, x22465, x22462);
  nand n22467(x22467, x22466, x22464);
  nand n22469(x22469, x22459, x22464);
  nand n22470(x22470, x21854, x83745);
  nand n22472(x22472, x22471, x21855);
  nand n22473(x22473, x22472, x22470);
  nand n22475(x22475, x21868, x22474);
  nand n22476(x22476, x21867, x22473);
  nand n22477(x22477, x22476, x22475);
  nand n22479(x22479, x22470, x22475);
  nand n22480(x22480, x21875, x21884);
  nand n22481(x22481, x21874, x21883);
  nand n22482(x22482, x22481, x22480);
  nand n22484(x22484, x21893, x22483);
  nand n22485(x22485, x21892, x22482);
  nand n22486(x22486, x22485, x22484);
  nand n22488(x22488, x22480, x22484);
  nand n22489(x22489, x21869, x83746);
  nand n22491(x22491, x22490, x21871);
  nand n22492(x22492, x22491, x22489);
  nand n22494(x22494, x21885, x22493);
  nand n22496(x22496, x22495, x22492);
  nand n22497(x22497, x22496, x22494);
  nand n22499(x22499, x22489, x22494);
  nand n22500(x22500, x21894, x83748);
  nand n22502(x22502, x22501, x21895);
  nand n22503(x22503, x22502, x22500);
  nand n22505(x22505, x21908, x22504);
  nand n22506(x22506, x21907, x22503);
  nand n22507(x22507, x22506, x22505);
  nand n22509(x22509, x22500, x22505);
  nand n22510(x22510, x21919, x21929);
  nand n22511(x22511, x21918, x21928);
  nand n22512(x22512, x22511, x22510);
  nand n22514(x22514, x21938, x22513);
  nand n22515(x22515, x21937, x22512);
  nand n22516(x22516, x22515, x22514);
  nand n22518(x22518, x22510, x22514);
  nand n22519(x22519, x21909, x21920);
  nand n22522(x22522, x22521, x22520);
  nand n22523(x22523, x22522, x22519);
  nand n22525(x22525, x21930, x22524);
  nand n22527(x22527, x22526, x22523);
  nand n22528(x22528, x22527, x22525);
  nand n22530(x22530, x21939, x21948);
  nand n22533(x22533, x22532, x22531);
  nand n22534(x22534, x22533, x22530);
  nand n22536(x22536, x21959, x22535);
  nand n22537(x22537, x21958, x22534);
  nand n22538(x22538, x22537, x22536);
  nand n22540(x22540, x21969, x21978);
  nand n22541(x22541, x21968, x21977);
  nand n22542(x22542, x22541, x22540);
  nand n22544(x22544, x21986, x22543);
  nand n22545(x22545, x21985, x22542);
  nand n22546(x22546, x22545, x22544);
  nand n22548(x22548, x22004, x83779);
  nand n22549(x22549, x22003, x21406);
  nand n22550(x22550, x22549, x22548);
  nand n22551(x22551, x22008, x83781);
  nand n22552(x22552, x22007, x21410);
  nand n22553(x22553, x22552, x22551);
  nand n22554(x22554, x22015, x83783);
  nand n22555(x22555, x22014, x22011);
  nand n22556(x22556, x22555, x22554);
  nand n22557(x22557, x83752, x83784);
  nand n22558(x22558, x22012, x22009);
  nand n22559(x22559, x22558, x22557);
  nand n22561(x22561, x22026, x83786);
  nand n22562(x22562, x22025, x22018);
  nand n22563(x22563, x22562, x22561);
  nand n22564(x22564, x22027, x83788);
  nand n22566(x22566, x22565, x22016);
  nand n22567(x22567, x22566, x22564);
  nand n22569(x22569, x22038, x83790);
  nand n22570(x22570, x22037, x22030);
  nand n22571(x22571, x22570, x22569);
  nand n22572(x22572, x22039, x83792);
  nand n22574(x22574, x22573, x22028);
  nand n22575(x22575, x22574, x22572);
  nand n22577(x22577, x22050, x83794);
  nand n22578(x22578, x22049, x22042);
  nand n22579(x22579, x22578, x22577);
  nand n22580(x22580, x22051, x83796);
  nand n22582(x22582, x22581, x22040);
  nand n22583(x22583, x22582, x22580);
  nand n22585(x22585, x22062, x83798);
  nand n22586(x22586, x22061, x22054);
  nand n22587(x22587, x22586, x22585);
  nand n22588(x22588, x22063, x83800);
  nand n22590(x22590, x22589, x22052);
  nand n22591(x22591, x22590, x22588);
  nand n22593(x22593, x22074, x83802);
  nand n22594(x22594, x22073, x22066);
  nand n22595(x22595, x22594, x22593);
  nand n22596(x22596, x22075, x83804);
  nand n22598(x22598, x22597, x22064);
  nand n22599(x22599, x22598, x22596);
  nand n22601(x22601, x83758, x22079);
  nand n22602(x22602, x21443, x22078);
  nand n22603(x22603, x22602, x22601);
  nand n22605(x22605, x22087, x22604);
  nand n22606(x22606, x22086, x22603);
  nand n22607(x22607, x22606, x22605);
  nand n22609(x22609, x22601, x22605);
  nand n22610(x22610, x22088, x83806);
  nand n22612(x22612, x22611, x22076);
  nand n22613(x22613, x22612, x22610);
  nand n22615(x22615, x83760, x22092);
  nand n22616(x22616, x21453, x22091);
  nand n22617(x22617, x22616, x22615);
  nand n22619(x22619, x22100, x22618);
  nand n22620(x22620, x22099, x22617);
  nand n22621(x22621, x22620, x22619);
  nand n22623(x22623, x22615, x22619);
  nand n22624(x22624, x22101, x83808);
  nand n22626(x22626, x22625, x22089);
  nand n22627(x22627, x22626, x22624);
  nand n22629(x22629, x83762, x22105);
  nand n22630(x22630, x21463, x22104);
  nand n22631(x22631, x22630, x22629);
  nand n22633(x22633, x22113, x22632);
  nand n22634(x22634, x22112, x22631);
  nand n22635(x22635, x22634, x22633);
  nand n22637(x22637, x22629, x22633);
  nand n22638(x22638, x22114, x83810);
  nand n22640(x22640, x22639, x22102);
  nand n22641(x22641, x22640, x22638);
  nand n22643(x22643, x83764, x22118);
  nand n22644(x22644, x21473, x22117);
  nand n22645(x22645, x22644, x22643);
  nand n22647(x22647, x22126, x22646);
  nand n22648(x22648, x22125, x22645);
  nand n22649(x22649, x22648, x22647);
  nand n22651(x22651, x22643, x22647);
  nand n22652(x22652, x22127, x83812);
  nand n22654(x22654, x22653, x22115);
  nand n22655(x22655, x22654, x22652);
  nand n22657(x22657, x22131, x22135);
  nand n22658(x22658, x22130, x22134);
  nand n22659(x22659, x22658, x22657);
  nand n22661(x22661, x22143, x22660);
  nand n22662(x22662, x22142, x22659);
  nand n22663(x22663, x22662, x22661);
  nand n22665(x22665, x22657, x22661);
  nand n22666(x22666, x83767, x83769);
  nand n22667(x22667, x22128, x22132);
  nand n22668(x22668, x22667, x22666);
  nand n22670(x22670, x22144, x22669);
  nand n22672(x22672, x22671, x22668);
  nand n22673(x22673, x22672, x22670);
  nand n22675(x22675, x22666, x22670);
  nand n22676(x22676, x22152, x22157);
  nand n22677(x22677, x22151, x22156);
  nand n22678(x22678, x22677, x22676);
  nand n22680(x22680, x22165, x22679);
  nand n22681(x22681, x22164, x22678);
  nand n22682(x22682, x22681, x22680);
  nand n22684(x22684, x22676, x22680);
  nand n22685(x22685, x22153, x83771);
  nand n22687(x22687, x22686, x22154);
  nand n22688(x22688, x22687, x22685);
  nand n22690(x22690, x22166, x22689);
  nand n22692(x22692, x22691, x22688);
  nand n22693(x22693, x22692, x22690);
  nand n22695(x22695, x22685, x22690);
  nand n22696(x22696, x22174, x22179);
  nand n22697(x22697, x22173, x22178);
  nand n22698(x22698, x22697, x22696);
  nand n22700(x22700, x22187, x22699);
  nand n22701(x22701, x22186, x22698);
  nand n22702(x22702, x22701, x22700);
  nand n22704(x22704, x22696, x22700);
  nand n22705(x22705, x22175, x83773);
  nand n22707(x22707, x22706, x22176);
  nand n22708(x22708, x22707, x22705);
  nand n22710(x22710, x22188, x22709);
  nand n22712(x22712, x22711, x22708);
  nand n22713(x22713, x22712, x22710);
  nand n22715(x22715, x22705, x22710);
  nand n22716(x22716, x22196, x22201);
  nand n22717(x22717, x22195, x22200);
  nand n22718(x22718, x22717, x22716);
  nand n22720(x22720, x22209, x22719);
  nand n22721(x22721, x22208, x22718);
  nand n22722(x22722, x22721, x22720);
  nand n22724(x22724, x22716, x22720);
  nand n22725(x22725, x22197, x83775);
  nand n22727(x22727, x22726, x22198);
  nand n22728(x22728, x22727, x22725);
  nand n22730(x22730, x22210, x22729);
  nand n22732(x22732, x22731, x22728);
  nand n22733(x22733, x22732, x22730);
  nand n22735(x22735, x22725, x22730);
  nand n22736(x22736, x22218, x22223);
  nand n22737(x22737, x22217, x22222);
  nand n22738(x22738, x22737, x22736);
  nand n22740(x22740, x22231, x22739);
  nand n22741(x22741, x22230, x22738);
  nand n22742(x22742, x22741, x22740);
  nand n22744(x22744, x22736, x22740);
  nand n22745(x22745, x22219, x83777);
  nand n22747(x22747, x22746, x22220);
  nand n22748(x22748, x22747, x22745);
  nand n22750(x22750, x22232, x22749);
  nand n22752(x22752, x22751, x22748);
  nand n22753(x22753, x22752, x22750);
  nand n22755(x22755, x22745, x22750);
  nand n22756(x22756, x22240, x22246);
  nand n22757(x22757, x22239, x22245);
  nand n22758(x22758, x22757, x22756);
  nand n22760(x22760, x22254, x22759);
  nand n22761(x22761, x22253, x22758);
  nand n22762(x22762, x22761, x22760);
  nand n22764(x22764, x22756, x22760);
  nand n22765(x22765, x22241, x83778);
  nand n22767(x22767, x22766, x22243);
  nand n22768(x22768, x22767, x22765);
  nand n22770(x22770, x22255, x22769);
  nand n22772(x22772, x22771, x22768);
  nand n22773(x22773, x22772, x22770);
  nand n22775(x22775, x22765, x22770);
  nand n22776(x22776, x22263, x22273);
  nand n22777(x22777, x22262, x22272);
  nand n22778(x22778, x22777, x22776);
  nand n22780(x22780, x22282, x22779);
  nand n22781(x22781, x22281, x22778);
  nand n22782(x22782, x22781, x22780);
  nand n22784(x22784, x22776, x22780);
  nand n22785(x22785, x22264, x22274);
  nand n22788(x22788, x22787, x22786);
  nand n22789(x22789, x22788, x22785);
  nand n22791(x22791, x22283, x22790);
  nand n22793(x22793, x22792, x22789);
  nand n22794(x22794, x22793, x22791);
  nand n22796(x22796, x22785, x22791);
  nand n22797(x22797, x22291, x22301);
  nand n22798(x22798, x22290, x22300);
  nand n22799(x22799, x22798, x22797);
  nand n22801(x22801, x22310, x22800);
  nand n22802(x22802, x22309, x22799);
  nand n22803(x22803, x22802, x22801);
  nand n22805(x22805, x22797, x22801);
  nand n22806(x22806, x22292, x22302);
  nand n22809(x22809, x22808, x22807);
  nand n22810(x22810, x22809, x22806);
  nand n22812(x22812, x22311, x22811);
  nand n22814(x22814, x22813, x22810);
  nand n22815(x22815, x22814, x22812);
  nand n22817(x22817, x22806, x22812);
  nand n22818(x22818, x22319, x22329);
  nand n22819(x22819, x22318, x22328);
  nand n22820(x22820, x22819, x22818);
  nand n22822(x22822, x22338, x22821);
  nand n22823(x22823, x22337, x22820);
  nand n22824(x22824, x22823, x22822);
  nand n22826(x22826, x22818, x22822);
  nand n22827(x22827, x22320, x22330);
  nand n22830(x22830, x22829, x22828);
  nand n22831(x22831, x22830, x22827);
  nand n22833(x22833, x22339, x22832);
  nand n22835(x22835, x22834, x22831);
  nand n22836(x22836, x22835, x22833);
  nand n22838(x22838, x22827, x22833);
  nand n22839(x22839, x22348, x22358);
  nand n22840(x22840, x22347, x22357);
  nand n22841(x22841, x22840, x22839);
  nand n22843(x22843, x22367, x22842);
  nand n22844(x22844, x22366, x22841);
  nand n22845(x22845, x22844, x22843);
  nand n22847(x22847, x22839, x22843);
  nand n22848(x22848, x22349, x22359);
  nand n22851(x22851, x22850, x22849);
  nand n22852(x22852, x22851, x22848);
  nand n22854(x22854, x22368, x22853);
  nand n22856(x22856, x22855, x22852);
  nand n22857(x22857, x22856, x22854);
  nand n22859(x22859, x22848, x22854);
  nand n22860(x22860, x22378, x22388);
  nand n22861(x22861, x22377, x22387);
  nand n22862(x22862, x22861, x22860);
  nand n22864(x22864, x22397, x22863);
  nand n22865(x22865, x22396, x22862);
  nand n22866(x22866, x22865, x22864);
  nand n22868(x22868, x22860, x22864);
  nand n22869(x22869, x22379, x22389);
  nand n22872(x22872, x22871, x22870);
  nand n22873(x22873, x22872, x22869);
  nand n22875(x22875, x22398, x22874);
  nand n22877(x22877, x22876, x22873);
  nand n22878(x22878, x22877, x22875);
  nand n22880(x22880, x22869, x22875);
  nand n22881(x22881, x22408, x22418);
  nand n22882(x22882, x22407, x22417);
  nand n22883(x22883, x22882, x22881);
  nand n22885(x22885, x22427, x22884);
  nand n22886(x22886, x22426, x22883);
  nand n22887(x22887, x22886, x22885);
  nand n22889(x22889, x22881, x22885);
  nand n22890(x22890, x22409, x22419);
  nand n22893(x22893, x22892, x22891);
  nand n22894(x22894, x22893, x22890);
  nand n22896(x22896, x22428, x22895);
  nand n22898(x22898, x22897, x22894);
  nand n22899(x22899, x22898, x22896);
  nand n22901(x22901, x22890, x22896);
  nand n22902(x22902, x22438, x22448);
  nand n22903(x22903, x22437, x22447);
  nand n22904(x22904, x22903, x22902);
  nand n22906(x22906, x22457, x22905);
  nand n22907(x22907, x22456, x22904);
  nand n22908(x22908, x22907, x22906);
  nand n22910(x22910, x22902, x22906);
  nand n22911(x22911, x22439, x22449);
  nand n22914(x22914, x22913, x22912);
  nand n22915(x22915, x22914, x22911);
  nand n22917(x22917, x22458, x22916);
  nand n22919(x22919, x22918, x22915);
  nand n22920(x22920, x22919, x22917);
  nand n22922(x22922, x22911, x22917);
  nand n22923(x22923, x22468, x22478);
  nand n22924(x22924, x22467, x22477);
  nand n22925(x22925, x22924, x22923);
  nand n22927(x22927, x22487, x22926);
  nand n22928(x22928, x22486, x22925);
  nand n22929(x22929, x22928, x22927);
  nand n22931(x22931, x22923, x22927);
  nand n22932(x22932, x22469, x22479);
  nand n22935(x22935, x22934, x22933);
  nand n22936(x22936, x22935, x22932);
  nand n22938(x22938, x22488, x22937);
  nand n22940(x22940, x22939, x22936);
  nand n22941(x22941, x22940, x22938);
  nand n22943(x22943, x22932, x22938);
  nand n22944(x22944, x22498, x22508);
  nand n22945(x22945, x22497, x22507);
  nand n22946(x22946, x22945, x22944);
  nand n22948(x22948, x22517, x22947);
  nand n22949(x22949, x22516, x22946);
  nand n22950(x22950, x22949, x22948);
  nand n22952(x22952, x22944, x22948);
  nand n22953(x22953, x22499, x22509);
  nand n22956(x22956, x22955, x22954);
  nand n22957(x22957, x22956, x22953);
  nand n22959(x22959, x22518, x22958);
  nand n22961(x22961, x22960, x22957);
  nand n22962(x22962, x22961, x22959);
  nand n22964(x22964, x22529, x22539);
  nand n22965(x22965, x22528, x22538);
  nand n22966(x22966, x22965, x22964);
  nand n22968(x22968, x22547, x22967);
  nand n22969(x22969, x22546, x22966);
  nand n22970(x22970, x22969, x22968);
  nand n22972(x22972, x83780, x83816);
  nand n22973(x22973, x22001, x22548);
  nand n22974(x22974, x22973, x22972);
  nand n22975(x22975, x83782, x83818);
  nand n22976(x22976, x22005, x22551);
  nand n22977(x22977, x22976, x22975);
  nand n22979(x22979, x22560, x83820);
  nand n22980(x22980, x22559, x22554);
  nand n22981(x22981, x22980, x22979);
  nand n22983(x22983, x83785, x83787);
  nand n22984(x22984, x22557, x22561);
  nand n22985(x22985, x22984, x22983);
  nand n22987(x22987, x22568, x22986);
  nand n22988(x22988, x22567, x22985);
  nand n22989(x22989, x22988, x22987);
  nand n22991(x22991, x22983, x22987);
  nand n22992(x22992, x83789, x83791);
  nand n22993(x22993, x22564, x22569);
  nand n22994(x22994, x22993, x22992);
  nand n22996(x22996, x22576, x22995);
  nand n22997(x22997, x22575, x22994);
  nand n22998(x22998, x22997, x22996);
  nand n23000(x23000, x22992, x22996);
  nand n23001(x23001, x83793, x83795);
  nand n23002(x23002, x22572, x22577);
  nand n23003(x23003, x23002, x23001);
  nand n23005(x23005, x22584, x23004);
  nand n23006(x23006, x22583, x23003);
  nand n23007(x23007, x23006, x23005);
  nand n23009(x23009, x23001, x23005);
  nand n23010(x23010, x83797, x83799);
  nand n23011(x23011, x22580, x22585);
  nand n23012(x23012, x23011, x23010);
  nand n23014(x23014, x22592, x23013);
  nand n23015(x23015, x22591, x23012);
  nand n23016(x23016, x23015, x23014);
  nand n23018(x23018, x23010, x23014);
  nand n23019(x23019, x83801, x83803);
  nand n23020(x23020, x22588, x22593);
  nand n23021(x23021, x23020, x23019);
  nand n23023(x23023, x22600, x23022);
  nand n23024(x23024, x22599, x23021);
  nand n23025(x23025, x23024, x23023);
  nand n23027(x23027, x23019, x23023);
  nand n23028(x23028, x22608, x83662);
  nand n23029(x23029, x22607, x18080);
  nand n23030(x23030, x23029, x23028);
  nand n23033(x23033, x83805, x22609);
  nand n23035(x23035, x22596, x23034);
  nand n23036(x23036, x23035, x23033);
  nand n23038(x23038, x22614, x23037);
  nand n23039(x23039, x22613, x23036);
  nand n23040(x23040, x23039, x23038);
  nand n23042(x23042, x23033, x23038);
  nand n23043(x23043, x22622, x83665);
  nand n23044(x23044, x22621, x19220);
  nand n23045(x23045, x23044, x23043);
  nand n23048(x23048, x83807, x22623);
  nand n23050(x23050, x22610, x23049);
  nand n23051(x23051, x23050, x23048);
  nand n23053(x23053, x22628, x23052);
  nand n23054(x23054, x22627, x23051);
  nand n23055(x23055, x23054, x23053);
  nand n23057(x23057, x23048, x23053);
  nand n23058(x23058, x22636, x83668);
  nand n23059(x23059, x22635, x19262);
  nand n23060(x23060, x23059, x23058);
  nand n23063(x23063, x83809, x22637);
  nand n23065(x23065, x22624, x23064);
  nand n23066(x23066, x23065, x23063);
  nand n23068(x23068, x22642, x23067);
  nand n23069(x23069, x22641, x23066);
  nand n23070(x23070, x23069, x23068);
  nand n23072(x23072, x23063, x23068);
  nand n23073(x23073, x22650, x83673);
  nand n23074(x23074, x22649, x20616);
  nand n23075(x23075, x23074, x23073);
  nand n23078(x23078, x83811, x22651);
  nand n23080(x23080, x22638, x23079);
  nand n23081(x23081, x23080, x23078);
  nand n23083(x23083, x22656, x23082);
  nand n23084(x23084, x22655, x23081);
  nand n23085(x23085, x23084, x23083);
  nand n23087(x23087, x23078, x23083);
  nand n23088(x23088, x22664, x83680);
  nand n23089(x23089, x22663, x20644);
  nand n23090(x23090, x23089, x23088);
  nand n23093(x23093, x83813, x22665);
  nand n23095(x23095, x22652, x23094);
  nand n23096(x23096, x23095, x23093);
  nand n23098(x23098, x22674, x23097);
  nand n23099(x23099, x22673, x23096);
  nand n23100(x23100, x23099, x23098);
  nand n23102(x23102, x23093, x23098);
  nand n23103(x23103, x22683, x83687);
  nand n23104(x23104, x22682, x20678);
  nand n23105(x23105, x23104, x23103);
  nand n23108(x23108, x22675, x22684);
  nand n23111(x23111, x23110, x23109);
  nand n23112(x23112, x23111, x23108);
  nand n23114(x23114, x22694, x23113);
  nand n23115(x23115, x22693, x23112);
  nand n23116(x23116, x23115, x23114);
  nand n23118(x23118, x23108, x23114);
  nand n23119(x23119, x22703, x83694);
  nand n23120(x23120, x22702, x20717);
  nand n23121(x23121, x23120, x23119);
  nand n23124(x23124, x22695, x22704);
  nand n23127(x23127, x23126, x23125);
  nand n23128(x23128, x23127, x23124);
  nand n23130(x23130, x22714, x23129);
  nand n23131(x23131, x22713, x23128);
  nand n23132(x23132, x23131, x23130);
  nand n23134(x23134, x23124, x23130);
  nand n23135(x23135, x22723, x83701);
  nand n23136(x23136, x22722, x20757);
  nand n23137(x23137, x23136, x23135);
  nand n23140(x23140, x22715, x22724);
  nand n23143(x23143, x23142, x23141);
  nand n23144(x23144, x23143, x23140);
  nand n23146(x23146, x22734, x23145);
  nand n23147(x23147, x22733, x23144);
  nand n23148(x23148, x23147, x23146);
  nand n23150(x23150, x23140, x23146);
  nand n23151(x23151, x22743, x83707);
  nand n23152(x23152, x22742, x20797);
  nand n23153(x23153, x23152, x23151);
  nand n23156(x23156, x22735, x22744);
  nand n23159(x23159, x23158, x23157);
  nand n23160(x23160, x23159, x23156);
  nand n23162(x23162, x22754, x23161);
  nand n23163(x23163, x22753, x23160);
  nand n23164(x23164, x23163, x23162);
  nand n23166(x23166, x23156, x23162);
  nand n23167(x23167, x22763, x83713);
  nand n23168(x23168, x22762, x21615);
  nand n23169(x23169, x23168, x23167);
  nand n23172(x23172, x22755, x22764);
  nand n23175(x23175, x23174, x23173);
  nand n23176(x23176, x23175, x23172);
  nand n23178(x23178, x22774, x23177);
  nand n23179(x23179, x22773, x23176);
  nand n23180(x23180, x23179, x23178);
  nand n23182(x23182, x23172, x23178);
  nand n23183(x23183, x22783, x83720);
  nand n23184(x23184, x22782, x21642);
  nand n23185(x23185, x23184, x23183);
  nand n23188(x23188, x22775, x22784);
  nand n23191(x23191, x23190, x23189);
  nand n23192(x23192, x23191, x23188);
  nand n23194(x23194, x22795, x23193);
  nand n23195(x23195, x22794, x23192);
  nand n23196(x23196, x23195, x23194);
  nand n23198(x23198, x23188, x23194);
  nand n23199(x23199, x22804, x83727);
  nand n23200(x23200, x22803, x21669);
  nand n23201(x23201, x23200, x23199);
  nand n23204(x23204, x22796, x22805);
  nand n23207(x23207, x23206, x23205);
  nand n23208(x23208, x23207, x23204);
  nand n23210(x23210, x22816, x23209);
  nand n23211(x23211, x22815, x23208);
  nand n23212(x23212, x23211, x23210);
  nand n23214(x23214, x23204, x23210);
  nand n23215(x23215, x22825, x83732);
  nand n23216(x23216, x22824, x21702);
  nand n23217(x23217, x23216, x23215);
  nand n23220(x23220, x22817, x22826);
  nand n23223(x23223, x23222, x23221);
  nand n23224(x23224, x23223, x23220);
  nand n23226(x23226, x22837, x23225);
  nand n23227(x23227, x22836, x23224);
  nand n23228(x23228, x23227, x23226);
  nand n23230(x23230, x23220, x23226);
  nand n23231(x23231, x22846, x83735);
  nand n23232(x23232, x22845, x21740);
  nand n23233(x23233, x23232, x23231);
  nand n23236(x23236, x22838, x22847);
  nand n23239(x23239, x23238, x23237);
  nand n23240(x23240, x23239, x23236);
  nand n23242(x23242, x22858, x23241);
  nand n23243(x23243, x22857, x23240);
  nand n23244(x23244, x23243, x23242);
  nand n23246(x23246, x23236, x23242);
  nand n23247(x23247, x22867, x83738);
  nand n23248(x23248, x22866, x21778);
  nand n23249(x23249, x23248, x23247);
  nand n23252(x23252, x22859, x22868);
  nand n23255(x23255, x23254, x23253);
  nand n23256(x23256, x23255, x23252);
  nand n23258(x23258, x22879, x23257);
  nand n23259(x23259, x22878, x23256);
  nand n23260(x23260, x23259, x23258);
  nand n23262(x23262, x23252, x23258);
  nand n23263(x23263, x22888, x83741);
  nand n23264(x23264, x22887, x21817);
  nand n23265(x23265, x23264, x23263);
  nand n23268(x23268, x22880, x22889);
  nand n23271(x23271, x23270, x23269);
  nand n23272(x23272, x23271, x23268);
  nand n23274(x23274, x22900, x23273);
  nand n23275(x23275, x22899, x23272);
  nand n23276(x23276, x23275, x23274);
  nand n23278(x23278, x23268, x23274);
  nand n23279(x23279, x22909, x83744);
  nand n23280(x23280, x22908, x21857);
  nand n23281(x23281, x23280, x23279);
  nand n23284(x23284, x22901, x22910);
  nand n23287(x23287, x23286, x23285);
  nand n23288(x23288, x23287, x23284);
  nand n23290(x23290, x22921, x23289);
  nand n23291(x23291, x22920, x23288);
  nand n23292(x23292, x23291, x23290);
  nand n23294(x23294, x23284, x23290);
  nand n23295(x23295, x22930, x83747);
  nand n23296(x23296, x22929, x21897);
  nand n23297(x23297, x23296, x23295);
  nand n23300(x23300, x22922, x22931);
  nand n23303(x23303, x23302, x23301);
  nand n23304(x23304, x23303, x23300);
  nand n23306(x23306, x22942, x23305);
  nand n23307(x23307, x22941, x23304);
  nand n23308(x23308, x23307, x23306);
  nand n23310(x23310, x23300, x23306);
  nand n23311(x23311, x22951, x21947);
  nand n23312(x23312, x22950, x21946);
  nand n23313(x23313, x23312, x23311);
  nand n23316(x23316, x22943, x22952);
  nand n23319(x23319, x23318, x23317);
  nand n23320(x23320, x23319, x23316);
  nand n23322(x23322, x22963, x23321);
  nand n23323(x23323, x22962, x23320);
  nand n23324(x23324, x23323, x23322);
  nand n23326(x23326, x22971, x21994);
  nand n23327(x23327, x22970, x21993);
  nand n23328(x23328, x23327, x23326);
  nand n23330(x23330, x83814, x83826);
  nand n23331(x23331, x22000, x21995);
  nand n23332(x23332, x23331, x23330);
  nand n23333(x23333, x22978, x83829);
  nand n23334(x23334, x22977, x22972);
  nand n23335(x23335, x23334, x23333);
  nand n23336(x23336, x22982, x83831);
  nand n23337(x23337, x22981, x22975);
  nand n23338(x23338, x23337, x23336);
  nand n23340(x23340, x22990, x83833);
  nand n23341(x23341, x22989, x22979);
  nand n23342(x23342, x23341, x23340);
  nand n23345(x23345, x22999, x22991);
  nand n23346(x23346, x22998, x23344);
  nand n23347(x23347, x23346, x23345);
  nand n23350(x23350, x23008, x23000);
  nand n23351(x23351, x23007, x23349);
  nand n23352(x23352, x23351, x23350);
  nand n23355(x23355, x23017, x23009);
  nand n23356(x23356, x23016, x23354);
  nand n23357(x23357, x23356, x23355);
  nand n23360(x23360, x23026, x23018);
  nand n23361(x23361, x23025, x23359);
  nand n23362(x23362, x23361, x23360);
  nand n23364(x23364, x23027, x23032);
  nand n23366(x23366, x23365, x23028);
  nand n23367(x23367, x23366, x23364);
  nand n23369(x23369, x23041, x23368);
  nand n23370(x23370, x23040, x23367);
  nand n23371(x23371, x23370, x23369);
  nand n23373(x23373, x23364, x23369);
  nand n23374(x23374, x23042, x23047);
  nand n23376(x23376, x23375, x23043);
  nand n23377(x23377, x23376, x23374);
  nand n23379(x23379, x23056, x23378);
  nand n23380(x23380, x23055, x23377);
  nand n23381(x23381, x23380, x23379);
  nand n23383(x23383, x23374, x23379);
  nand n23384(x23384, x23057, x23062);
  nand n23386(x23386, x23385, x23058);
  nand n23387(x23387, x23386, x23384);
  nand n23389(x23389, x23071, x23388);
  nand n23390(x23390, x23070, x23387);
  nand n23391(x23391, x23390, x23389);
  nand n23393(x23393, x23384, x23389);
  nand n23394(x23394, x23072, x23077);
  nand n23396(x23396, x23395, x23073);
  nand n23397(x23397, x23396, x23394);
  nand n23399(x23399, x23086, x23398);
  nand n23400(x23400, x23085, x23397);
  nand n23401(x23401, x23400, x23399);
  nand n23403(x23403, x23394, x23399);
  nand n23404(x23404, x23087, x23092);
  nand n23406(x23406, x23405, x23088);
  nand n23407(x23407, x23406, x23404);
  nand n23409(x23409, x23101, x23408);
  nand n23410(x23410, x23100, x23407);
  nand n23411(x23411, x23410, x23409);
  nand n23413(x23413, x23404, x23409);
  nand n23414(x23414, x23102, x23107);
  nand n23416(x23416, x23415, x23103);
  nand n23417(x23417, x23416, x23414);
  nand n23419(x23419, x23117, x23418);
  nand n23420(x23420, x23116, x23417);
  nand n23421(x23421, x23420, x23419);
  nand n23423(x23423, x23414, x23419);
  nand n23424(x23424, x23118, x23123);
  nand n23426(x23426, x23425, x23119);
  nand n23427(x23427, x23426, x23424);
  nand n23429(x23429, x23133, x23428);
  nand n23430(x23430, x23132, x23427);
  nand n23431(x23431, x23430, x23429);
  nand n23433(x23433, x23424, x23429);
  nand n23434(x23434, x23134, x23139);
  nand n23436(x23436, x23435, x23135);
  nand n23437(x23437, x23436, x23434);
  nand n23439(x23439, x23149, x23438);
  nand n23440(x23440, x23148, x23437);
  nand n23441(x23441, x23440, x23439);
  nand n23443(x23443, x23434, x23439);
  nand n23444(x23444, x23150, x23155);
  nand n23446(x23446, x23445, x23151);
  nand n23447(x23447, x23446, x23444);
  nand n23449(x23449, x23165, x23448);
  nand n23450(x23450, x23164, x23447);
  nand n23451(x23451, x23450, x23449);
  nand n23453(x23453, x23444, x23449);
  nand n23454(x23454, x23166, x23171);
  nand n23456(x23456, x23455, x23167);
  nand n23457(x23457, x23456, x23454);
  nand n23459(x23459, x23181, x23458);
  nand n23460(x23460, x23180, x23457);
  nand n23461(x23461, x23460, x23459);
  nand n23463(x23463, x23454, x23459);
  nand n23464(x23464, x23182, x23187);
  nand n23466(x23466, x23465, x23183);
  nand n23467(x23467, x23466, x23464);
  nand n23469(x23469, x23197, x23468);
  nand n23470(x23470, x23196, x23467);
  nand n23471(x23471, x23470, x23469);
  nand n23473(x23473, x23464, x23469);
  nand n23474(x23474, x23198, x23203);
  nand n23476(x23476, x23475, x23199);
  nand n23477(x23477, x23476, x23474);
  nand n23479(x23479, x23213, x23478);
  nand n23480(x23480, x23212, x23477);
  nand n23481(x23481, x23480, x23479);
  nand n23483(x23483, x23474, x23479);
  nand n23484(x23484, x23214, x23219);
  nand n23486(x23486, x23485, x23215);
  nand n23487(x23487, x23486, x23484);
  nand n23489(x23489, x23229, x23488);
  nand n23490(x23490, x23228, x23487);
  nand n23491(x23491, x23490, x23489);
  nand n23493(x23493, x23484, x23489);
  nand n23494(x23494, x23230, x23235);
  nand n23496(x23496, x23495, x23231);
  nand n23497(x23497, x23496, x23494);
  nand n23499(x23499, x23245, x23498);
  nand n23500(x23500, x23244, x23497);
  nand n23501(x23501, x23500, x23499);
  nand n23503(x23503, x23494, x23499);
  nand n23504(x23504, x23246, x23251);
  nand n23506(x23506, x23505, x23247);
  nand n23507(x23507, x23506, x23504);
  nand n23509(x23509, x23261, x23508);
  nand n23510(x23510, x23260, x23507);
  nand n23511(x23511, x23510, x23509);
  nand n23513(x23513, x23504, x23509);
  nand n23514(x23514, x23262, x23267);
  nand n23516(x23516, x23515, x23263);
  nand n23517(x23517, x23516, x23514);
  nand n23519(x23519, x23277, x23518);
  nand n23520(x23520, x23276, x23517);
  nand n23521(x23521, x23520, x23519);
  nand n23523(x23523, x23514, x23519);
  nand n23524(x23524, x23278, x23283);
  nand n23526(x23526, x23525, x23279);
  nand n23527(x23527, x23526, x23524);
  nand n23529(x23529, x23293, x23528);
  nand n23530(x23530, x23292, x23527);
  nand n23531(x23531, x23530, x23529);
  nand n23533(x23533, x23524, x23529);
  nand n23534(x23534, x23294, x23299);
  nand n23536(x23536, x23535, x23295);
  nand n23537(x23537, x23536, x23534);
  nand n23539(x23539, x23309, x23538);
  nand n23540(x23540, x23308, x23537);
  nand n23541(x23541, x23540, x23539);
  nand n23543(x23543, x23534, x23539);
  nand n23544(x23544, x23310, x23315);
  nand n23546(x23546, x23545, x23311);
  nand n23547(x23547, x23546, x23544);
  nand n23549(x23549, x23325, x23548);
  nand n23550(x23550, x23324, x23547);
  nand n23551(x23551, x23550, x23549);
  nand n23553(x23553, x83827, x83828);
  nand n23554(x23554, x23330, x21998);
  nand n23555(x23555, x23554, x23553);
  nand n23557(x23557, x83815, x23556);
  nand n23558(x23558, x22550, x23555);
  nand n23559(x23559, x23558, x23557);
  nand n23560(x23560, x23553, x23557);
  nand n23561(x23561, x83817, x83839);
  nand n23562(x23562, x22553, x22974);
  nand n23563(x23563, x23562, x23561);
  nand n23565(x23565, x83819, x83841);
  nand n23566(x23566, x22556, x23335);
  nand n23567(x23567, x23566, x23565);
  nand n23569(x23569, x83830, x23339);
  nand n23570(x23570, x23333, x23338);
  nand n23571(x23571, x23570, x23569);
  nand n23573(x23573, x83821, x23572);
  nand n23574(x23574, x22563, x23571);
  nand n23575(x23575, x23574, x23573);
  nand n23577(x23577, x23569, x23573);
  nand n23578(x23578, x83832, x23343);
  nand n23579(x23579, x23336, x23342);
  nand n23580(x23580, x23579, x23578);
  nand n23582(x23582, x83822, x23581);
  nand n23583(x23583, x22571, x23580);
  nand n23584(x23584, x23583, x23582);
  nand n23586(x23586, x23578, x23582);
  nand n23587(x23587, x83834, x23348);
  nand n23588(x23588, x23340, x23347);
  nand n23589(x23589, x23588, x23587);
  nand n23591(x23591, x83823, x23590);
  nand n23592(x23592, x22579, x23589);
  nand n23593(x23593, x23592, x23591);
  nand n23595(x23595, x23587, x23591);
  nand n23596(x23596, x83835, x23353);
  nand n23597(x23597, x23345, x23352);
  nand n23598(x23598, x23597, x23596);
  nand n23600(x23600, x83824, x23599);
  nand n23601(x23601, x22587, x23598);
  nand n23602(x23602, x23601, x23600);
  nand n23604(x23604, x23596, x23600);
  nand n23605(x23605, x83836, x23358);
  nand n23606(x23606, x23350, x23357);
  nand n23607(x23607, x23606, x23605);
  nand n23609(x23609, x83825, x23608);
  nand n23610(x23610, x22595, x23607);
  nand n23611(x23611, x23610, x23609);
  nand n23613(x23613, x23605, x23609);
  nand n23614(x23614, x83837, x23363);
  nand n23615(x23615, x23355, x23362);
  nand n23616(x23616, x23615, x23614);
  nand n23618(x23618, x23031, x23617);
  nand n23619(x23619, x23030, x23616);
  nand n23620(x23620, x23619, x23618);
  nand n23622(x23622, x23614, x23618);
  nand n23623(x23623, x83838, x23372);
  nand n23624(x23624, x23360, x23371);
  nand n23625(x23625, x23624, x23623);
  nand n23627(x23627, x23046, x23626);
  nand n23628(x23628, x23045, x23625);
  nand n23629(x23629, x23628, x23627);
  nand n23631(x23631, x23623, x23627);
  nand n23632(x23632, x23373, x23382);
  nand n23634(x23634, x23633, x23381);
  nand n23635(x23635, x23634, x23632);
  nand n23637(x23637, x23061, x23636);
  nand n23638(x23638, x23060, x23635);
  nand n23639(x23639, x23638, x23637);
  nand n23641(x23641, x23632, x23637);
  nand n23642(x23642, x23383, x23392);
  nand n23644(x23644, x23643, x23391);
  nand n23645(x23645, x23644, x23642);
  nand n23647(x23647, x23076, x23646);
  nand n23648(x23648, x23075, x23645);
  nand n23649(x23649, x23648, x23647);
  nand n23651(x23651, x23642, x23647);
  nand n23652(x23652, x23393, x23402);
  nand n23654(x23654, x23653, x23401);
  nand n23655(x23655, x23654, x23652);
  nand n23657(x23657, x23091, x23656);
  nand n23658(x23658, x23090, x23655);
  nand n23659(x23659, x23658, x23657);
  nand n23661(x23661, x23652, x23657);
  nand n23662(x23662, x23403, x23412);
  nand n23664(x23664, x23663, x23411);
  nand n23665(x23665, x23664, x23662);
  nand n23667(x23667, x23106, x23666);
  nand n23668(x23668, x23105, x23665);
  nand n23669(x23669, x23668, x23667);
  nand n23671(x23671, x23662, x23667);
  nand n23672(x23672, x23413, x23422);
  nand n23674(x23674, x23673, x23421);
  nand n23675(x23675, x23674, x23672);
  nand n23677(x23677, x23122, x23676);
  nand n23678(x23678, x23121, x23675);
  nand n23679(x23679, x23678, x23677);
  nand n23681(x23681, x23672, x23677);
  nand n23682(x23682, x23423, x23432);
  nand n23684(x23684, x23683, x23431);
  nand n23685(x23685, x23684, x23682);
  nand n23687(x23687, x23138, x23686);
  nand n23688(x23688, x23137, x23685);
  nand n23689(x23689, x23688, x23687);
  nand n23691(x23691, x23682, x23687);
  nand n23692(x23692, x23433, x23442);
  nand n23694(x23694, x23693, x23441);
  nand n23695(x23695, x23694, x23692);
  nand n23697(x23697, x23154, x23696);
  nand n23698(x23698, x23153, x23695);
  nand n23699(x23699, x23698, x23697);
  nand n23701(x23701, x23692, x23697);
  nand n23702(x23702, x23443, x23452);
  nand n23704(x23704, x23703, x23451);
  nand n23705(x23705, x23704, x23702);
  nand n23707(x23707, x23170, x23706);
  nand n23708(x23708, x23169, x23705);
  nand n23709(x23709, x23708, x23707);
  nand n23711(x23711, x23702, x23707);
  nand n23712(x23712, x23453, x23462);
  nand n23714(x23714, x23713, x23461);
  nand n23715(x23715, x23714, x23712);
  nand n23717(x23717, x23186, x23716);
  nand n23718(x23718, x23185, x23715);
  nand n23719(x23719, x23718, x23717);
  nand n23721(x23721, x23712, x23717);
  nand n23722(x23722, x23463, x23472);
  nand n23724(x23724, x23723, x23471);
  nand n23725(x23725, x23724, x23722);
  nand n23727(x23727, x23202, x23726);
  nand n23728(x23728, x23201, x23725);
  nand n23729(x23729, x23728, x23727);
  nand n23731(x23731, x23722, x23727);
  nand n23732(x23732, x23473, x23482);
  nand n23734(x23734, x23733, x23481);
  nand n23735(x23735, x23734, x23732);
  nand n23737(x23737, x23218, x23736);
  nand n23738(x23738, x23217, x23735);
  nand n23739(x23739, x23738, x23737);
  nand n23741(x23741, x23732, x23737);
  nand n23742(x23742, x23483, x23492);
  nand n23744(x23744, x23743, x23491);
  nand n23745(x23745, x23744, x23742);
  nand n23747(x23747, x23234, x23746);
  nand n23748(x23748, x23233, x23745);
  nand n23749(x23749, x23748, x23747);
  nand n23751(x23751, x23742, x23747);
  nand n23752(x23752, x23493, x23502);
  nand n23754(x23754, x23753, x23501);
  nand n23755(x23755, x23754, x23752);
  nand n23757(x23757, x23250, x23756);
  nand n23758(x23758, x23249, x23755);
  nand n23759(x23759, x23758, x23757);
  nand n23761(x23761, x23752, x23757);
  nand n23762(x23762, x23503, x23512);
  nand n23764(x23764, x23763, x23511);
  nand n23765(x23765, x23764, x23762);
  nand n23767(x23767, x23266, x23766);
  nand n23768(x23768, x23265, x23765);
  nand n23769(x23769, x23768, x23767);
  nand n23771(x23771, x23762, x23767);
  nand n23772(x23772, x23513, x23522);
  nand n23774(x23774, x23773, x23521);
  nand n23775(x23775, x23774, x23772);
  nand n23777(x23777, x23282, x23776);
  nand n23778(x23778, x23281, x23775);
  nand n23779(x23779, x23778, x23777);
  nand n23781(x23781, x23772, x23777);
  nand n23782(x23782, x23523, x23532);
  nand n23784(x23784, x23783, x23531);
  nand n23785(x23785, x23784, x23782);
  nand n23787(x23787, x23298, x23786);
  nand n23788(x23788, x23297, x23785);
  nand n23789(x23789, x23788, x23787);
  nand n23791(x23791, x23782, x23787);
  nand n23792(x23792, x23533, x23542);
  nand n23794(x23794, x23793, x23541);
  nand n23795(x23795, x23794, x23792);
  nand n23797(x23797, x23314, x23796);
  nand n23798(x23798, x23313, x23795);
  nand n23799(x23799, x23798, x23797);
  nand n23801(x23801, x23792, x23797);
  nand n23802(x23802, x23543, x23552);
  nand n23804(x23804, x23803, x23551);
  nand n23805(x23805, x23804, x23802);
  nand n23807(x23807, x23329, x23806);
  nand n23808(x23808, x23328, x23805);
  nand n23809(x23809, x23808, x23807);
  nand n23811(x23811, x23560, x23564);
  nand n23813(x23813, x23812, x23563);
  nand n23814(x23814, x23813, x23811);
  nand n23815(x23815, x83840, x23568);
  nand n23816(x23816, x23561, x23567);
  nand n23817(x23817, x23816, x23815);
  nand n23819(x23819, x83842, x23576);
  nand n23820(x23820, x23565, x23575);
  nand n23821(x23821, x23820, x23819);
  nand n23823(x23823, x23577, x23585);
  nand n23825(x23825, x23824, x23584);
  nand n23826(x23826, x23825, x23823);
  nand n23828(x23828, x23586, x23594);
  nand n23830(x23830, x23829, x23593);
  nand n23831(x23831, x23830, x23828);
  nand n23833(x23833, x23595, x23603);
  nand n23835(x23835, x23834, x23602);
  nand n23836(x23836, x23835, x23833);
  nand n23838(x23838, x23604, x23612);
  nand n23840(x23840, x23839, x23611);
  nand n23841(x23841, x23840, x23838);
  nand n23843(x23843, x23613, x23621);
  nand n23845(x23845, x23844, x23620);
  nand n23846(x23846, x23845, x23843);
  nand n23848(x23848, x23622, x23630);
  nand n23850(x23850, x23849, x23629);
  nand n23851(x23851, x23850, x23848);
  nand n23853(x23853, x23631, x23640);
  nand n23855(x23855, x23854, x23639);
  nand n23856(x23856, x23855, x23853);
  nand n23858(x23858, x23641, x23650);
  nand n23860(x23860, x23859, x23649);
  nand n23861(x23861, x23860, x23858);
  nand n23863(x23863, x23651, x23660);
  nand n23865(x23865, x23864, x23659);
  nand n23866(x23866, x23865, x23863);
  nand n23868(x23868, x23661, x23670);
  nand n23870(x23870, x23869, x23669);
  nand n23871(x23871, x23870, x23868);
  nand n23873(x23873, x23671, x23680);
  nand n23875(x23875, x23874, x23679);
  nand n23876(x23876, x23875, x23873);
  nand n23878(x23878, x23681, x23690);
  nand n23880(x23880, x23879, x23689);
  nand n23881(x23881, x23880, x23878);
  nand n23883(x23883, x23691, x23700);
  nand n23885(x23885, x23884, x23699);
  nand n23886(x23886, x23885, x23883);
  nand n23888(x23888, x23701, x23710);
  nand n23890(x23890, x23889, x23709);
  nand n23891(x23891, x23890, x23888);
  nand n23893(x23893, x23711, x23720);
  nand n23895(x23895, x23894, x23719);
  nand n23896(x23896, x23895, x23893);
  nand n23898(x23898, x23721, x23730);
  nand n23900(x23900, x23899, x23729);
  nand n23901(x23901, x23900, x23898);
  nand n23903(x23903, x23731, x23740);
  nand n23905(x23905, x23904, x23739);
  nand n23906(x23906, x23905, x23903);
  nand n23908(x23908, x23741, x23750);
  nand n23910(x23910, x23909, x23749);
  nand n23911(x23911, x23910, x23908);
  nand n23913(x23913, x23751, x23760);
  nand n23915(x23915, x23914, x23759);
  nand n23916(x23916, x23915, x23913);
  nand n23918(x23918, x23761, x23770);
  nand n23920(x23920, x23919, x23769);
  nand n23921(x23921, x23920, x23918);
  nand n23923(x23923, x23771, x23780);
  nand n23925(x23925, x23924, x23779);
  nand n23926(x23926, x23925, x23923);
  nand n23928(x23928, x23781, x23790);
  nand n23930(x23930, x23929, x23789);
  nand n23931(x23931, x23930, x23928);
  nand n23933(x23933, x23791, x23800);
  nand n23935(x23935, x23934, x23799);
  nand n23936(x23936, x23935, x23933);
  nand n23938(x23938, x23801, x23810);
  nand n23940(x23940, x23939, x23809);
  nand n23941(x23941, x23940, x23938);
  nand n23968(x23968, x23818, x23943);
  nand n23969(x23969, x23968, x23815);
  nand n23970(x23970, x23822, x23944);
  nand n23971(x23971, x23970, x23819);
  nand n23972(x23972, x23822, x23818);
  nand n23974(x23974, x23827, x23945);
  nand n23975(x23975, x23974, x23823);
  nand n23976(x23976, x23827, x23822);
  nand n23978(x23978, x23832, x23946);
  nand n23979(x23979, x23978, x23828);
  nand n23980(x23980, x23832, x23827);
  nand n23982(x23982, x23837, x23947);
  nand n23983(x23983, x23982, x23833);
  nand n23984(x23984, x23837, x23832);
  nand n23986(x23986, x23842, x23948);
  nand n23987(x23987, x23986, x23838);
  nand n23988(x23988, x23842, x23837);
  nand n23990(x23990, x23847, x23949);
  nand n23991(x23991, x23990, x23843);
  nand n23992(x23992, x23847, x23842);
  nand n23994(x23994, x23852, x23950);
  nand n23995(x23995, x23994, x23848);
  nand n23996(x23996, x23852, x23847);
  nand n23998(x23998, x23857, x23951);
  nand n23999(x23999, x23998, x23853);
  nand n24000(x24000, x23857, x23852);
  nand n24002(x24002, x23862, x23952);
  nand n24003(x24003, x24002, x23858);
  nand n24004(x24004, x23862, x23857);
  nand n24006(x24006, x23867, x23953);
  nand n24007(x24007, x24006, x23863);
  nand n24008(x24008, x23867, x23862);
  nand n24010(x24010, x23872, x23954);
  nand n24011(x24011, x24010, x23868);
  nand n24012(x24012, x23872, x23867);
  nand n24014(x24014, x23877, x23955);
  nand n24015(x24015, x24014, x23873);
  nand n24016(x24016, x23877, x23872);
  nand n24018(x24018, x23882, x23956);
  nand n24019(x24019, x24018, x23878);
  nand n24020(x24020, x23882, x23877);
  nand n24022(x24022, x23887, x23957);
  nand n24023(x24023, x24022, x23883);
  nand n24024(x24024, x23887, x23882);
  nand n24026(x24026, x23892, x23958);
  nand n24027(x24027, x24026, x23888);
  nand n24028(x24028, x23892, x23887);
  nand n24030(x24030, x23897, x23959);
  nand n24031(x24031, x24030, x23893);
  nand n24032(x24032, x23897, x23892);
  nand n24034(x24034, x23902, x23960);
  nand n24035(x24035, x24034, x23898);
  nand n24036(x24036, x23902, x23897);
  nand n24038(x24038, x23907, x23961);
  nand n24039(x24039, x24038, x23903);
  nand n24040(x24040, x23907, x23902);
  nand n24042(x24042, x23912, x23962);
  nand n24043(x24043, x24042, x23908);
  nand n24044(x24044, x23912, x23907);
  nand n24046(x24046, x23917, x23963);
  nand n24047(x24047, x24046, x23913);
  nand n24048(x24048, x23917, x23912);
  nand n24050(x24050, x23922, x23964);
  nand n24051(x24051, x24050, x23918);
  nand n24052(x24052, x23922, x23917);
  nand n24054(x24054, x23927, x23965);
  nand n24055(x24055, x24054, x23923);
  nand n24056(x24056, x23927, x23922);
  nand n24058(x24058, x23932, x23966);
  nand n24059(x24059, x24058, x23928);
  nand n24060(x24060, x23932, x23927);
  nand n24062(x24062, x23937, x23967);
  nand n24063(x24063, x24062, x23933);
  nand n24064(x24064, x23937, x23932);
  nand n24067(x24067, x23973, x23943);
  nand n24069(x24069, x24067, x24068);
  nand n24070(x24070, x23977, x23969);
  nand n24072(x24072, x24070, x24071);
  nand n24073(x24073, x23981, x23971);
  nand n24075(x24075, x24073, x24074);
  nand n24076(x24076, x23981, x23973);
  nand n24078(x24078, x23985, x23975);
  nand n24080(x24080, x24078, x24079);
  nand n24081(x24081, x23985, x23977);
  nand n24083(x24083, x23989, x23979);
  nand n24085(x24085, x24083, x24084);
  nand n24086(x24086, x23989, x23981);
  nand n24088(x24088, x23993, x23983);
  nand n24090(x24090, x24088, x24089);
  nand n24091(x24091, x23993, x23985);
  nand n24093(x24093, x23997, x23987);
  nand n24095(x24095, x24093, x24094);
  nand n24096(x24096, x23997, x23989);
  nand n24098(x24098, x24001, x23991);
  nand n24100(x24100, x24098, x24099);
  nand n24101(x24101, x24001, x23993);
  nand n24103(x24103, x24005, x23995);
  nand n24105(x24105, x24103, x24104);
  nand n24106(x24106, x24005, x23997);
  nand n24108(x24108, x24009, x23999);
  nand n24110(x24110, x24108, x24109);
  nand n24111(x24111, x24009, x24001);
  nand n24113(x24113, x24013, x24003);
  nand n24115(x24115, x24113, x24114);
  nand n24116(x24116, x24013, x24005);
  nand n24118(x24118, x24017, x24007);
  nand n24120(x24120, x24118, x24119);
  nand n24121(x24121, x24017, x24009);
  nand n24123(x24123, x24021, x24011);
  nand n24125(x24125, x24123, x24124);
  nand n24126(x24126, x24021, x24013);
  nand n24128(x24128, x24025, x24015);
  nand n24130(x24130, x24128, x24129);
  nand n24131(x24131, x24025, x24017);
  nand n24133(x24133, x24029, x24019);
  nand n24135(x24135, x24133, x24134);
  nand n24136(x24136, x24029, x24021);
  nand n24138(x24138, x24033, x24023);
  nand n24140(x24140, x24138, x24139);
  nand n24141(x24141, x24033, x24025);
  nand n24143(x24143, x24037, x24027);
  nand n24145(x24145, x24143, x24144);
  nand n24146(x24146, x24037, x24029);
  nand n24148(x24148, x24041, x24031);
  nand n24150(x24150, x24148, x24149);
  nand n24151(x24151, x24041, x24033);
  nand n24153(x24153, x24045, x24035);
  nand n24155(x24155, x24153, x24154);
  nand n24156(x24156, x24045, x24037);
  nand n24158(x24158, x24049, x24039);
  nand n24160(x24160, x24158, x24159);
  nand n24161(x24161, x24049, x24041);
  nand n24163(x24163, x24053, x24043);
  nand n24165(x24165, x24163, x24164);
  nand n24166(x24166, x24053, x24045);
  nand n24168(x24168, x24057, x24047);
  nand n24170(x24170, x24168, x24169);
  nand n24171(x24171, x24057, x24049);
  nand n24173(x24173, x24061, x24051);
  nand n24175(x24175, x24173, x24174);
  nand n24176(x24176, x24061, x24053);
  nand n24178(x24178, x24065, x24055);
  nand n24180(x24180, x24178, x24179);
  nand n24181(x24181, x24065, x24057);
  nand n24185(x24185, x24077, x23943);
  nand n24187(x24187, x24185, x24186);
  nand n24188(x24188, x24082, x23969);
  nand n24190(x24190, x24188, x24189);
  nand n24191(x24191, x24087, x24069);
  nand n24193(x24193, x24191, x24192);
  nand n24194(x24194, x24092, x24072);
  nand n24196(x24196, x24194, x24195);
  nand n24197(x24197, x24097, x24075);
  nand n24199(x24199, x24197, x24198);
  nand n24200(x24200, x24097, x24077);
  nand n24202(x24202, x24102, x24080);
  nand n24204(x24204, x24202, x24203);
  nand n24205(x24205, x24102, x24082);
  nand n24207(x24207, x24107, x24085);
  nand n24209(x24209, x24207, x24208);
  nand n24210(x24210, x24107, x24087);
  nand n24212(x24212, x24112, x24090);
  nand n24214(x24214, x24212, x24213);
  nand n24215(x24215, x24112, x24092);
  nand n24217(x24217, x24117, x24095);
  nand n24219(x24219, x24217, x24218);
  nand n24220(x24220, x24117, x24097);
  nand n24222(x24222, x24122, x24100);
  nand n24224(x24224, x24222, x24223);
  nand n24225(x24225, x24122, x24102);
  nand n24227(x24227, x24127, x24105);
  nand n24229(x24229, x24227, x24228);
  nand n24230(x24230, x24127, x24107);
  nand n24232(x24232, x24132, x24110);
  nand n24234(x24234, x24232, x24233);
  nand n24235(x24235, x24132, x24112);
  nand n24237(x24237, x24137, x24115);
  nand n24239(x24239, x24237, x24238);
  nand n24240(x24240, x24137, x24117);
  nand n24242(x24242, x24142, x24120);
  nand n24244(x24244, x24242, x24243);
  nand n24245(x24245, x24142, x24122);
  nand n24247(x24247, x24147, x24125);
  nand n24249(x24249, x24247, x24248);
  nand n24250(x24250, x24147, x24127);
  nand n24252(x24252, x24152, x24130);
  nand n24254(x24254, x24252, x24253);
  nand n24255(x24255, x24152, x24132);
  nand n24257(x24257, x24157, x24135);
  nand n24259(x24259, x24257, x24258);
  nand n24260(x24260, x24157, x24137);
  nand n24262(x24262, x24162, x24140);
  nand n24264(x24264, x24262, x24263);
  nand n24265(x24265, x24162, x24142);
  nand n24267(x24267, x24167, x24145);
  nand n24269(x24269, x24267, x24268);
  nand n24270(x24270, x24167, x24147);
  nand n24272(x24272, x24172, x24150);
  nand n24274(x24274, x24272, x24273);
  nand n24275(x24275, x24172, x24152);
  nand n24277(x24277, x24177, x24155);
  nand n24279(x24279, x24277, x24278);
  nand n24280(x24280, x24177, x24157);
  nand n24282(x24282, x24182, x24160);
  nand n24284(x24284, x24282, x24283);
  nand n24285(x24285, x24182, x24162);
  nand n24291(x24291, x24201, x23943);
  nand n24293(x24293, x24291, x24292);
  nand n24294(x24294, x24206, x23969);
  nand n24296(x24296, x24294, x24295);
  nand n24297(x24297, x24211, x24069);
  nand n24299(x24299, x24297, x24298);
  nand n24300(x24300, x24216, x24072);
  nand n24302(x24302, x24300, x24301);
  nand n24303(x24303, x24221, x24187);
  nand n24305(x24305, x24303, x24304);
  nand n24306(x24306, x24226, x24190);
  nand n24308(x24308, x24306, x24307);
  nand n24309(x24309, x24231, x24193);
  nand n24311(x24311, x24309, x24310);
  nand n24312(x24312, x24236, x24196);
  nand n24314(x24314, x24312, x24313);
  nand n24315(x24315, x24241, x24199);
  nand n24317(x24317, x24315, x24316);
  nand n24318(x24318, x24241, x24201);
  nand n24320(x24320, x24246, x24204);
  nand n24322(x24322, x24320, x24321);
  nand n24323(x24323, x24246, x24206);
  nand n24325(x24325, x24251, x24209);
  nand n24327(x24327, x24325, x24326);
  nand n24328(x24328, x24251, x24211);
  nand n24330(x24330, x24256, x24214);
  nand n24332(x24332, x24330, x24331);
  nand n24333(x24333, x24256, x24216);
  nand n24335(x24335, x24261, x24219);
  nand n24337(x24337, x24335, x24336);
  nand n24338(x24338, x24261, x24221);
  nand n24340(x24340, x24266, x24224);
  nand n24342(x24342, x24340, x24341);
  nand n24343(x24343, x24266, x24226);
  nand n24345(x24345, x24271, x24229);
  nand n24347(x24347, x24345, x24346);
  nand n24348(x24348, x24271, x24231);
  nand n24350(x24350, x24276, x24234);
  nand n24352(x24352, x24350, x24351);
  nand n24353(x24353, x24276, x24236);
  nand n24355(x24355, x24281, x24239);
  nand n24357(x24357, x24355, x24356);
  nand n24358(x24358, x24281, x24241);
  nand n24360(x24360, x24286, x24244);
  nand n24362(x24362, x24360, x24361);
  nand n24363(x24363, x24286, x24246);
  nand n24371(x24371, x24319, x23943);
  nand n24373(x24373, x24371, x24372);
  nand n24374(x24374, x24324, x23969);
  nand n24376(x24376, x24374, x24375);
  nand n24377(x24377, x24329, x24069);
  nand n24379(x24379, x24377, x24378);
  nand n24380(x24380, x24334, x24072);
  nand n24382(x24382, x24380, x24381);
  nand n24383(x24383, x24339, x24187);
  nand n24385(x24385, x24383, x24384);
  nand n24386(x24386, x24344, x24190);
  nand n24388(x24388, x24386, x24387);
  nand n24389(x24389, x24349, x24193);
  nand n24391(x24391, x24389, x24390);
  nand n24392(x24392, x24354, x24196);
  nand n24394(x24394, x24392, x24393);
  nand n24395(x24395, x24359, x24293);
  nand n24397(x24397, x24395, x24396);
  nand n24398(x24398, x24364, x24296);
  nand n24400(x24400, x24398, x24399);
  nand n24401(x24401, x23817, x23811);
  nand n24402(x24402, x24401, x23968);
  nand n24404(x24404, x23822, x23969);
  nand n24405(x24405, x23821, x24066);
  nand n24406(x24406, x24405, x24404);
  nand n24408(x24408, x23827, x24069);
  nand n24409(x24409, x23826, x24183);
  nand n24410(x24410, x24409, x24408);
  nand n24412(x24412, x23832, x24072);
  nand n24413(x24413, x23831, x24184);
  nand n24414(x24414, x24413, x24412);
  nand n24416(x24416, x23837, x24187);
  nand n24417(x24417, x23836, x24287);
  nand n24418(x24418, x24417, x24416);
  nand n24420(x24420, x23842, x24190);
  nand n24421(x24421, x23841, x24288);
  nand n24422(x24422, x24421, x24420);
  nand n24424(x24424, x23847, x24193);
  nand n24425(x24425, x23846, x24289);
  nand n24426(x24426, x24425, x24424);
  nand n24428(x24428, x23852, x24196);
  nand n24429(x24429, x23851, x24290);
  nand n24430(x24430, x24429, x24428);
  nand n24432(x24432, x23857, x24293);
  nand n24434(x24434, x23856, x24433);
  nand n24435(x24435, x24434, x24432);
  nand n24437(x24437, x23862, x24296);
  nand n24439(x24439, x23861, x24438);
  nand n24440(x24440, x24439, x24437);
  nand n24442(x24442, x23867, x24299);
  nand n24443(x24443, x23866, x24365);
  nand n24444(x24444, x24443, x24442);
  nand n24446(x24446, x23872, x24302);
  nand n24447(x24447, x23871, x24366);
  nand n24448(x24448, x24447, x24446);
  nand n24450(x24450, x23877, x24305);
  nand n24451(x24451, x23876, x24367);
  nand n24452(x24452, x24451, x24450);
  nand n24454(x24454, x23882, x24308);
  nand n24455(x24455, x23881, x24368);
  nand n24456(x24456, x24455, x24454);
  nand n24458(x24458, x23887, x24311);
  nand n24459(x24459, x23886, x24369);
  nand n24460(x24460, x24459, x24458);
  nand n24462(x24462, x23892, x24314);
  nand n24463(x24463, x23891, x24370);
  nand n24464(x24464, x24463, x24462);
  nand n24466(x24466, x23897, x24373);
  nand n24468(x24468, x23896, x24467);
  nand n24469(x24469, x24468, x24466);
  nand n24471(x24471, x23902, x24376);
  nand n24473(x24473, x23901, x24472);
  nand n24474(x24474, x24473, x24471);
  nand n24476(x24476, x23907, x24379);
  nand n24478(x24478, x23906, x24477);
  nand n24479(x24479, x24478, x24476);
  nand n24481(x24481, x23912, x24382);
  nand n24483(x24483, x23911, x24482);
  nand n24484(x24484, x24483, x24481);
  nand n24486(x24486, x23917, x24385);
  nand n24488(x24488, x23916, x24487);
  nand n24489(x24489, x24488, x24486);
  nand n24491(x24491, x23922, x24388);
  nand n24493(x24493, x23921, x24492);
  nand n24494(x24494, x24493, x24491);
  nand n24496(x24496, x23927, x24391);
  nand n24498(x24498, x23926, x24497);
  nand n24499(x24499, x24498, x24496);
  nand n24501(x24501, x23932, x24394);
  nand n24503(x24503, x23931, x24502);
  nand n24504(x24504, x24503, x24501);
  nand n24506(x24506, x23937, x24397);
  nand n24508(x24508, x23936, x24507);
  nand n24509(x24509, x24508, x24506);
  nand n24511(x24511, x23942, x24400);
  nand n24513(x24513, x23941, x24512);
  nand n24514(x24514, x24513, x24511);
  nand n24516(x24516, x16980, x16974);
  nand n24518(x24518, x16986, x16980);
  nand n24520(x24520, x16992, x16986);
  nand n24522(x24522, x16998, x16992);
  nand n24524(x24524, x17004, x16998);
  nand n24526(x24526, x17010, x17004);
  nand n24528(x24528, x17016, x17010);
  nand n24530(x24530, x17022, x17016);
  nand n24532(x24532, x17028, x17022);
  nand n24534(x24534, x17034, x17028);
  nand n24536(x24536, x17040, x17034);
  nand n24538(x24538, x17046, x17040);
  nand n24540(x24540, x17052, x17046);
  nand n24542(x24542, x17058, x17052);
  nand n24544(x24544, x17064, x17058);
  nand n24546(x24546, x17070, x17064);
  nand n24548(x24548, x17076, x17070);
  nand n24550(x24550, x17082, x17076);
  nand n24552(x24552, x17088, x17082);
  nand n24554(x24554, x17094, x17088);
  nand n24556(x24556, x17100, x17094);
  nand n24558(x24558, x17106, x17100);
  nand n24560(x24560, x17112, x17106);
  nand n24562(x24562, x17118, x17112);
  nand n24564(x24564, x17124, x17118);
  nand n24566(x24566, x17130, x17124);
  nand n24568(x24568, x17136, x17130);
  nand n24570(x24570, x17142, x17136);
  nand n24572(x24572, x17148, x17142);
  nand n24574(x24574, x17154, x17148);
  nand n24576(x24576, x24519, x16974);
  nand n24577(x24577, x24521, x24517);
  nand n24579(x24579, x24523, x24519);
  nand n24581(x24581, x24525, x24521);
  nand n24583(x24583, x24527, x24523);
  nand n24585(x24585, x24529, x24525);
  nand n24587(x24587, x24531, x24527);
  nand n24589(x24589, x24533, x24529);
  nand n24591(x24591, x24535, x24531);
  nand n24593(x24593, x24537, x24533);
  nand n24595(x24595, x24539, x24535);
  nand n24597(x24597, x24541, x24537);
  nand n24599(x24599, x24543, x24539);
  nand n24601(x24601, x24545, x24541);
  nand n24603(x24603, x24547, x24543);
  nand n24605(x24605, x24549, x24545);
  nand n24607(x24607, x24551, x24547);
  nand n24609(x24609, x24553, x24549);
  nand n24611(x24611, x24555, x24551);
  nand n24613(x24613, x24557, x24553);
  nand n24615(x24615, x24559, x24555);
  nand n24617(x24617, x24561, x24557);
  nand n24619(x24619, x24563, x24559);
  nand n24621(x24621, x24565, x24561);
  nand n24623(x24623, x24567, x24563);
  nand n24625(x24625, x24569, x24565);
  nand n24627(x24627, x24571, x24567);
  nand n24629(x24629, x24573, x24569);
  nand n24631(x24631, x24575, x24571);
  nand n24633(x24633, x24580, x16974);
  nand n24634(x24634, x24582, x24517);
  nand n24635(x24635, x24584, x83848);
  nand n24636(x24636, x24586, x24578);
  nand n24638(x24638, x24588, x24580);
  nand n24640(x24640, x24590, x24582);
  nand n24642(x24642, x24592, x24584);
  nand n24644(x24644, x24594, x24586);
  nand n24646(x24646, x24596, x24588);
  nand n24648(x24648, x24598, x24590);
  nand n24650(x24650, x24600, x24592);
  nand n24652(x24652, x24602, x24594);
  nand n24654(x24654, x24604, x24596);
  nand n24656(x24656, x24606, x24598);
  nand n24658(x24658, x24608, x24600);
  nand n24660(x24660, x24610, x24602);
  nand n24662(x24662, x24612, x24604);
  nand n24664(x24664, x24614, x24606);
  nand n24666(x24666, x24616, x24608);
  nand n24668(x24668, x24618, x24610);
  nand n24670(x24670, x24620, x24612);
  nand n24672(x24672, x24622, x24614);
  nand n24674(x24674, x24624, x24616);
  nand n24676(x24676, x24626, x24618);
  nand n24678(x24678, x24628, x24620);
  nand n24680(x24680, x24630, x24622);
  nand n24682(x24682, x24632, x24624);
  nand n24684(x24684, x24639, x16974);
  nand n24685(x24685, x24641, x24517);
  nand n24686(x24686, x24643, x83848);
  nand n24687(x24687, x24645, x24578);
  nand n24688(x24688, x24647, x83849);
  nand n24689(x24689, x24649, x83850);
  nand n24690(x24690, x24651, x83851);
  nand n24691(x24691, x24653, x24637);
  nand n24692(x24692, x24655, x24639);
  nand n24694(x24694, x24657, x24641);
  nand n24696(x24696, x24659, x24643);
  nand n24698(x24698, x24661, x24645);
  nand n24700(x24700, x24663, x24647);
  nand n24702(x24702, x24665, x24649);
  nand n24704(x24704, x24667, x24651);
  nand n24706(x24706, x24669, x24653);
  nand n24708(x24708, x24671, x24655);
  nand n24710(x24710, x24673, x24657);
  nand n24712(x24712, x24675, x24659);
  nand n24714(x24714, x24677, x24661);
  nand n24716(x24716, x24679, x24663);
  nand n24718(x24718, x24681, x24665);
  nand n24720(x24720, x24683, x24667);
  nand n24722(x24722, x24693, x16974);
  nand n24723(x24723, x24695, x24517);
  nand n24724(x24724, x24697, x83848);
  nand n24725(x24725, x24699, x24578);
  nand n24726(x24726, x24701, x83849);
  nand n24727(x24727, x24703, x83850);
  nand n24728(x24728, x24705, x83851);
  nand n24729(x24729, x24707, x24637);
  nand n24730(x24730, x24709, x83852);
  nand n24731(x24731, x24711, x83853);
  nand n24732(x24732, x24713, x83854);
  nand n24733(x24733, x24715, x83855);
  nand n24734(x24734, x24717, x83856);
  nand n24735(x24735, x24719, x83857);
  nand n24736(x24736, x24721, x83858);
  nand n24737(x24737, x72052, x72047);
  nand n24738(x24738, x24737, x24516);
  nand n24740(x24740, x16986, x24517);
  nand n24741(x24741, x72057, x24516);
  nand n24742(x24742, x24741, x24740);
  nand n24744(x24744, x16992, x83848);
  nand n24745(x24745, x72062, x24576);
  nand n24746(x24746, x24745, x24744);
  nand n24748(x24748, x16998, x24578);
  nand n24749(x24749, x72067, x24577);
  nand n24750(x24750, x24749, x24748);
  nand n24752(x24752, x17004, x83849);
  nand n24753(x24753, x72072, x24633);
  nand n24754(x24754, x24753, x24752);
  nand n24756(x24756, x17010, x83850);
  nand n24757(x24757, x72077, x24634);
  nand n24758(x24758, x24757, x24756);
  nand n24760(x24760, x17016, x83851);
  nand n24761(x24761, x72082, x24635);
  nand n24762(x24762, x24761, x24760);
  nand n24764(x24764, x17022, x24637);
  nand n24765(x24765, x72087, x24636);
  nand n24766(x24766, x24765, x24764);
  nand n24768(x24768, x17028, x83852);
  nand n24769(x24769, x72092, x24684);
  nand n24770(x24770, x24769, x24768);
  nand n24772(x24772, x17034, x83853);
  nand n24773(x24773, x72097, x24685);
  nand n24774(x24774, x24773, x24772);
  nand n24776(x24776, x17040, x83854);
  nand n24777(x24777, x72102, x24686);
  nand n24778(x24778, x24777, x24776);
  nand n24780(x24780, x17046, x83855);
  nand n24781(x24781, x72107, x24687);
  nand n24782(x24782, x24781, x24780);
  nand n24784(x24784, x17052, x83856);
  nand n24785(x24785, x72112, x24688);
  nand n24786(x24786, x24785, x24784);
  nand n24788(x24788, x17058, x83857);
  nand n24789(x24789, x72117, x24689);
  nand n24790(x24790, x24789, x24788);
  nand n24792(x24792, x17064, x83858);
  nand n24793(x24793, x72122, x24690);
  nand n24794(x24794, x24793, x24792);
  nand n24796(x24796, x17070, x83859);
  nand n24797(x24797, x72127, x24691);
  nand n24798(x24798, x24797, x24796);
  nand n24800(x24800, x17076, x83860);
  nand n24801(x24801, x72132, x24722);
  nand n24802(x24802, x24801, x24800);
  nand n24804(x24804, x17082, x83861);
  nand n24805(x24805, x72137, x24723);
  nand n24806(x24806, x24805, x24804);
  nand n24808(x24808, x17088, x83862);
  nand n24809(x24809, x72142, x24724);
  nand n24810(x24810, x24809, x24808);
  nand n24812(x24812, x17094, x83863);
  nand n24813(x24813, x72147, x24725);
  nand n24814(x24814, x24813, x24812);
  nand n24816(x24816, x17100, x83864);
  nand n24817(x24817, x72152, x24726);
  nand n24818(x24818, x24817, x24816);
  nand n24820(x24820, x17106, x83865);
  nand n24821(x24821, x72157, x24727);
  nand n24822(x24822, x24821, x24820);
  nand n24824(x24824, x17112, x83866);
  nand n24825(x24825, x72162, x24728);
  nand n24826(x24826, x24825, x24824);
  nand n24828(x24828, x17118, x83867);
  nand n24829(x24829, x72167, x24729);
  nand n24830(x24830, x24829, x24828);
  nand n24832(x24832, x17124, x83868);
  nand n24833(x24833, x72172, x24730);
  nand n24834(x24834, x24833, x24832);
  nand n24836(x24836, x17130, x83869);
  nand n24837(x24837, x72177, x24731);
  nand n24838(x24838, x24837, x24836);
  nand n24840(x24840, x17136, x83870);
  nand n24841(x24841, x72182, x24732);
  nand n24842(x24842, x24841, x24840);
  nand n24844(x24844, x17142, x83871);
  nand n24845(x24845, x72187, x24733);
  nand n24846(x24846, x24845, x24844);
  nand n24848(x24848, x17148, x83872);
  nand n24849(x24849, x72192, x24734);
  nand n24850(x24850, x24849, x24848);
  nand n24852(x24852, x17154, x83873);
  nand n24853(x24853, x72197, x24735);
  nand n24854(x24854, x24853, x24852);
  nand n24856(x24856, x17160, x83874);
  nand n24857(x24857, x72202, x24736);
  nand n24858(x24858, x24857, x24856);
  nand n24861(x24861, x72127, x16797);
  nand n24863(x24863, x72132, x16800);
  nand n24865(x24865, x72137, x16803);
  nand n24867(x24867, x72142, x16806);
  nand n24869(x24869, x72147, x16809);
  nand n24871(x24871, x72152, x16812);
  nand n24873(x24873, x72157, x16815);
  nand n24875(x24875, x72162, x16818);
  nand n24877(x24877, x72167, x16821);
  nand n24879(x24879, x72172, x16824);
  nand n24881(x24881, x72177, x16827);
  nand n24883(x24883, x72182, x16830);
  nand n24885(x24885, x72187, x16833);
  nand n24887(x24887, x72192, x16836);
  nand n24889(x24889, x72197, x16839);
  nand n24891(x24891, x72202, x16842);
  nand n24893(x24893, x16974, x16843);
  nand n24894(x24894, x16980, x16844);
  nand n24895(x24895, x16986, x16845);
  nand n24896(x24896, x16992, x16846);
  nand n24897(x24897, x16998, x16847);
  nand n24898(x24898, x17004, x16848);
  nand n24899(x24899, x17010, x16849);
  nand n24900(x24900, x17016, x16850);
  nand n24901(x24901, x17022, x16851);
  nand n24902(x24902, x17028, x16852);
  nand n24903(x24903, x17034, x16853);
  nand n24904(x24904, x17040, x16854);
  nand n24905(x24905, x17046, x16855);
  nand n24906(x24906, x17052, x16856);
  nand n24907(x24907, x17058, x16857);
  nand n24908(x24908, x17064, x16858);
  nand n24909(x24909, x17070, x16859);
  nand n24910(x24910, x17076, x16860);
  nand n24911(x24911, x17082, x16861);
  nand n24912(x24912, x17088, x16862);
  nand n24913(x24913, x17094, x16863);
  nand n24914(x24914, x17100, x16864);
  nand n24915(x24915, x17106, x16865);
  nand n24916(x24916, x17112, x16866);
  nand n24917(x24917, x17118, x16867);
  nand n24918(x24918, x17124, x16868);
  nand n24919(x24919, x17130, x16869);
  nand n24920(x24920, x17136, x16870);
  nand n24921(x24921, x17142, x16871);
  nand n24922(x24922, x17148, x16872);
  nand n24923(x24923, x17154, x16873);
  nand n24924(x24924, x17160, x16874);
  nand n24925(x24925, x24893, x17904);
  nand n24927(x24927, x24894, x17911);
  nand n24929(x24929, x24895, x17926);
  nand n24931(x24931, x24896, x17950);
  nand n24933(x24933, x24897, x17981);
  nand n24935(x24935, x24898, x18020);
  nand n24937(x24937, x24899, x18068);
  nand n24939(x24939, x24900, x18123);
  nand n24941(x24941, x24901, x18186);
  nand n24943(x24943, x24902, x18258);
  nand n24945(x24945, x24903, x18337);
  nand n24947(x24947, x24904, x18424);
  nand n24949(x24949, x24905, x18520);
  nand n24951(x24951, x24906, x18623);
  nand n24953(x24953, x24907, x18734);
  nand n24955(x24955, x24908, x18854);
  nand n24957(x24957, x24909, x24861);
  nand n24959(x24959, x24910, x24863);
  nand n24961(x24961, x24911, x24865);
  nand n24963(x24963, x24912, x24867);
  nand n24965(x24965, x24913, x24869);
  nand n24967(x24967, x24914, x24871);
  nand n24969(x24969, x24915, x24873);
  nand n24971(x24971, x24916, x24875);
  nand n24973(x24973, x24917, x24877);
  nand n24975(x24975, x24918, x24879);
  nand n24977(x24977, x24919, x24881);
  nand n24979(x24979, x24920, x24883);
  nand n24981(x24981, x24921, x24885);
  nand n24983(x24983, x24922, x24887);
  nand n24985(x24985, x24923, x24889);
  nand n24987(x24987, x24924, x24891);
  nand n24989(x24989, x16843, x72047);
  nand n24990(x24990, x16843, x72052);
  nand n24991(x24991, x24990, x17904);
  nand n24992(x24992, x16843, x72057);
  nand n24993(x24993, x24992, x17905);
  nand n24994(x24994, x16843, x72062);
  nand n24995(x24995, x24994, x17909);
  nand n24996(x24996, x16843, x72067);
  nand n24997(x24997, x24996, x17915);
  nand n24998(x24998, x16843, x72072);
  nand n24999(x24999, x24998, x17922);
  nand n25000(x25000, x16843, x72077);
  nand n25001(x25001, x25000, x17932);
  nand n25002(x25002, x16843, x72082);
  nand n25003(x25003, x25002, x17944);
  nand n25004(x25004, x16843, x72087);
  nand n25005(x25005, x25004, x17957);
  nand n25006(x25006, x16843, x72092);
  nand n25007(x25007, x25006, x17973);
  nand n25008(x25008, x16843, x72097);
  nand n25009(x25009, x25008, x17991);
  nand n25010(x25010, x16843, x72102);
  nand n25011(x25011, x25010, x18010);
  nand n25012(x25012, x16843, x72107);
  nand n25013(x25013, x25012, x18032);
  nand n25014(x25014, x16843, x72112);
  nand n25015(x25015, x25014, x18056);
  nand n25016(x25016, x16843, x72117);
  nand n25017(x25017, x25016, x18081);
  nand n25018(x25018, x16843, x72122);
  nand n25019(x25019, x25018, x18109);
  nand n25020(x25020, x16843, x72127);
  nand n25021(x25021, x25020, x18139);
  nand n25022(x25022, x16843, x72132);
  nand n25023(x25023, x25022, x18170);
  nand n25024(x25024, x16843, x72137);
  nand n25025(x25025, x25024, x18204);
  nand n25026(x25026, x16843, x72142);
  nand n25027(x25027, x25026, x18240);
  nand n25028(x25028, x16843, x72147);
  nand n25029(x25029, x25028, x18277);
  nand n25030(x25030, x16843, x72152);
  nand n25031(x25031, x25030, x18317);
  nand n25032(x25032, x16843, x72157);
  nand n25033(x25033, x25032, x18359);
  nand n25034(x25034, x16843, x72162);
  nand n25035(x25035, x25034, x18402);
  nand n25036(x25036, x16843, x72167);
  nand n25037(x25037, x25036, x18448);
  nand n25038(x25038, x16843, x72172);
  nand n25039(x25039, x25038, x18496);
  nand n25040(x25040, x16843, x72177);
  nand n25041(x25041, x25040, x18545);
  nand n25042(x25042, x16843, x72182);
  nand n25043(x25043, x25042, x18597);
  nand n25044(x25044, x16843, x72187);
  nand n25045(x25045, x25044, x18651);
  nand n25046(x25046, x16843, x72192);
  nand n25047(x25047, x25046, x18706);
  nand n25048(x25048, x16843, x72197);
  nand n25049(x25049, x25048, x18764);
  nand n25050(x25050, x16843, x72202);
  nand n25051(x25051, x25050, x18824);
  nand n25052(x25052, x16844, x83875);
  nand n25053(x25053, x16844, x24991);
  nand n25054(x25054, x16752, x83875);
  nand n25055(x25055, x16844, x24993);
  nand n25056(x25056, x25055, x25054);
  nand n25057(x25057, x16752, x24991);
  nand n25058(x25058, x16844, x24995);
  nand n25059(x25059, x25058, x25057);
  nand n25060(x25060, x16752, x24993);
  nand n25061(x25061, x16844, x24997);
  nand n25062(x25062, x25061, x25060);
  nand n25063(x25063, x16752, x24995);
  nand n25064(x25064, x16844, x24999);
  nand n25065(x25065, x25064, x25063);
  nand n25066(x25066, x16752, x24997);
  nand n25067(x25067, x16844, x25001);
  nand n25068(x25068, x25067, x25066);
  nand n25069(x25069, x16752, x24999);
  nand n25070(x25070, x16844, x25003);
  nand n25071(x25071, x25070, x25069);
  nand n25072(x25072, x16752, x25001);
  nand n25073(x25073, x16844, x25005);
  nand n25074(x25074, x25073, x25072);
  nand n25075(x25075, x16752, x25003);
  nand n25076(x25076, x16844, x25007);
  nand n25077(x25077, x25076, x25075);
  nand n25078(x25078, x16752, x25005);
  nand n25079(x25079, x16844, x25009);
  nand n25080(x25080, x25079, x25078);
  nand n25081(x25081, x16752, x25007);
  nand n25082(x25082, x16844, x25011);
  nand n25083(x25083, x25082, x25081);
  nand n25084(x25084, x16752, x25009);
  nand n25085(x25085, x16844, x25013);
  nand n25086(x25086, x25085, x25084);
  nand n25087(x25087, x16752, x25011);
  nand n25088(x25088, x16844, x25015);
  nand n25089(x25089, x25088, x25087);
  nand n25090(x25090, x16752, x25013);
  nand n25091(x25091, x16844, x25017);
  nand n25092(x25092, x25091, x25090);
  nand n25093(x25093, x16752, x25015);
  nand n25094(x25094, x16844, x25019);
  nand n25095(x25095, x25094, x25093);
  nand n25096(x25096, x16752, x25017);
  nand n25097(x25097, x16844, x25021);
  nand n25098(x25098, x25097, x25096);
  nand n25099(x25099, x16752, x25019);
  nand n25100(x25100, x16844, x25023);
  nand n25101(x25101, x25100, x25099);
  nand n25102(x25102, x16752, x25021);
  nand n25103(x25103, x16844, x25025);
  nand n25104(x25104, x25103, x25102);
  nand n25105(x25105, x16752, x25023);
  nand n25106(x25106, x16844, x25027);
  nand n25107(x25107, x25106, x25105);
  nand n25108(x25108, x16752, x25025);
  nand n25109(x25109, x16844, x25029);
  nand n25110(x25110, x25109, x25108);
  nand n25111(x25111, x16752, x25027);
  nand n25112(x25112, x16844, x25031);
  nand n25113(x25113, x25112, x25111);
  nand n25114(x25114, x16752, x25029);
  nand n25115(x25115, x16844, x25033);
  nand n25116(x25116, x25115, x25114);
  nand n25117(x25117, x16752, x25031);
  nand n25118(x25118, x16844, x25035);
  nand n25119(x25119, x25118, x25117);
  nand n25120(x25120, x16752, x25033);
  nand n25121(x25121, x16844, x25037);
  nand n25122(x25122, x25121, x25120);
  nand n25123(x25123, x16752, x25035);
  nand n25124(x25124, x16844, x25039);
  nand n25125(x25125, x25124, x25123);
  nand n25126(x25126, x16752, x25037);
  nand n25127(x25127, x16844, x25041);
  nand n25128(x25128, x25127, x25126);
  nand n25129(x25129, x16752, x25039);
  nand n25130(x25130, x16844, x25043);
  nand n25131(x25131, x25130, x25129);
  nand n25132(x25132, x16752, x25041);
  nand n25133(x25133, x16844, x25045);
  nand n25134(x25134, x25133, x25132);
  nand n25135(x25135, x16752, x25043);
  nand n25136(x25136, x16844, x25047);
  nand n25137(x25137, x25136, x25135);
  nand n25138(x25138, x16752, x25045);
  nand n25139(x25139, x16844, x25049);
  nand n25140(x25140, x25139, x25138);
  nand n25141(x25141, x16752, x25047);
  nand n25142(x25142, x16844, x25051);
  nand n25143(x25143, x25142, x25141);
  nand n25144(x25144, x16845, x83876);
  nand n25145(x25145, x16845, x83877);
  nand n25146(x25146, x16845, x25056);
  nand n25147(x25147, x16845, x25059);
  nand n25148(x25148, x16755, x83876);
  nand n25149(x25149, x16845, x25062);
  nand n25150(x25150, x25149, x25148);
  nand n25151(x25151, x16755, x83877);
  nand n25152(x25152, x16845, x25065);
  nand n25153(x25153, x25152, x25151);
  nand n25154(x25154, x16755, x25056);
  nand n25155(x25155, x16845, x25068);
  nand n25156(x25156, x25155, x25154);
  nand n25157(x25157, x16755, x25059);
  nand n25158(x25158, x16845, x25071);
  nand n25159(x25159, x25158, x25157);
  nand n25160(x25160, x16755, x25062);
  nand n25161(x25161, x16845, x25074);
  nand n25162(x25162, x25161, x25160);
  nand n25163(x25163, x16755, x25065);
  nand n25164(x25164, x16845, x25077);
  nand n25165(x25165, x25164, x25163);
  nand n25166(x25166, x16755, x25068);
  nand n25167(x25167, x16845, x25080);
  nand n25168(x25168, x25167, x25166);
  nand n25169(x25169, x16755, x25071);
  nand n25170(x25170, x16845, x25083);
  nand n25171(x25171, x25170, x25169);
  nand n25172(x25172, x16755, x25074);
  nand n25173(x25173, x16845, x25086);
  nand n25174(x25174, x25173, x25172);
  nand n25175(x25175, x16755, x25077);
  nand n25176(x25176, x16845, x25089);
  nand n25177(x25177, x25176, x25175);
  nand n25178(x25178, x16755, x25080);
  nand n25179(x25179, x16845, x25092);
  nand n25180(x25180, x25179, x25178);
  nand n25181(x25181, x16755, x25083);
  nand n25182(x25182, x16845, x25095);
  nand n25183(x25183, x25182, x25181);
  nand n25184(x25184, x16755, x25086);
  nand n25185(x25185, x16845, x25098);
  nand n25186(x25186, x25185, x25184);
  nand n25187(x25187, x16755, x25089);
  nand n25188(x25188, x16845, x25101);
  nand n25189(x25189, x25188, x25187);
  nand n25190(x25190, x16755, x25092);
  nand n25191(x25191, x16845, x25104);
  nand n25192(x25192, x25191, x25190);
  nand n25193(x25193, x16755, x25095);
  nand n25194(x25194, x16845, x25107);
  nand n25195(x25195, x25194, x25193);
  nand n25196(x25196, x16755, x25098);
  nand n25197(x25197, x16845, x25110);
  nand n25198(x25198, x25197, x25196);
  nand n25199(x25199, x16755, x25101);
  nand n25200(x25200, x16845, x25113);
  nand n25201(x25201, x25200, x25199);
  nand n25202(x25202, x16755, x25104);
  nand n25203(x25203, x16845, x25116);
  nand n25204(x25204, x25203, x25202);
  nand n25205(x25205, x16755, x25107);
  nand n25206(x25206, x16845, x25119);
  nand n25207(x25207, x25206, x25205);
  nand n25208(x25208, x16755, x25110);
  nand n25209(x25209, x16845, x25122);
  nand n25210(x25210, x25209, x25208);
  nand n25211(x25211, x16755, x25113);
  nand n25212(x25212, x16845, x25125);
  nand n25213(x25213, x25212, x25211);
  nand n25214(x25214, x16755, x25116);
  nand n25215(x25215, x16845, x25128);
  nand n25216(x25216, x25215, x25214);
  nand n25217(x25217, x16755, x25119);
  nand n25218(x25218, x16845, x25131);
  nand n25219(x25219, x25218, x25217);
  nand n25220(x25220, x16755, x25122);
  nand n25221(x25221, x16845, x25134);
  nand n25222(x25222, x25221, x25220);
  nand n25223(x25223, x16755, x25125);
  nand n25224(x25224, x16845, x25137);
  nand n25225(x25225, x25224, x25223);
  nand n25226(x25226, x16755, x25128);
  nand n25227(x25227, x16845, x25140);
  nand n25228(x25228, x25227, x25226);
  nand n25229(x25229, x16755, x25131);
  nand n25230(x25230, x16845, x25143);
  nand n25231(x25231, x25230, x25229);
  nand n25232(x25232, x16846, x83878);
  nand n25233(x25233, x16846, x83879);
  nand n25234(x25234, x16846, x83880);
  nand n25235(x25235, x16846, x83881);
  nand n25236(x25236, x16846, x25150);
  nand n25237(x25237, x16846, x25153);
  nand n25238(x25238, x16846, x25156);
  nand n25239(x25239, x16846, x25159);
  nand n25240(x25240, x16758, x83878);
  nand n25241(x25241, x16846, x25162);
  nand n25242(x25242, x25241, x25240);
  nand n25243(x25243, x16758, x83879);
  nand n25244(x25244, x16846, x25165);
  nand n25245(x25245, x25244, x25243);
  nand n25246(x25246, x16758, x83880);
  nand n25247(x25247, x16846, x25168);
  nand n25248(x25248, x25247, x25246);
  nand n25249(x25249, x16758, x83881);
  nand n25250(x25250, x16846, x25171);
  nand n25251(x25251, x25250, x25249);
  nand n25252(x25252, x16758, x25150);
  nand n25253(x25253, x16846, x25174);
  nand n25254(x25254, x25253, x25252);
  nand n25255(x25255, x16758, x25153);
  nand n25256(x25256, x16846, x25177);
  nand n25257(x25257, x25256, x25255);
  nand n25258(x25258, x16758, x25156);
  nand n25259(x25259, x16846, x25180);
  nand n25260(x25260, x25259, x25258);
  nand n25261(x25261, x16758, x25159);
  nand n25262(x25262, x16846, x25183);
  nand n25263(x25263, x25262, x25261);
  nand n25264(x25264, x16758, x25162);
  nand n25265(x25265, x16846, x25186);
  nand n25266(x25266, x25265, x25264);
  nand n25267(x25267, x16758, x25165);
  nand n25268(x25268, x16846, x25189);
  nand n25269(x25269, x25268, x25267);
  nand n25270(x25270, x16758, x25168);
  nand n25271(x25271, x16846, x25192);
  nand n25272(x25272, x25271, x25270);
  nand n25273(x25273, x16758, x25171);
  nand n25274(x25274, x16846, x25195);
  nand n25275(x25275, x25274, x25273);
  nand n25276(x25276, x16758, x25174);
  nand n25277(x25277, x16846, x25198);
  nand n25278(x25278, x25277, x25276);
  nand n25279(x25279, x16758, x25177);
  nand n25280(x25280, x16846, x25201);
  nand n25281(x25281, x25280, x25279);
  nand n25282(x25282, x16758, x25180);
  nand n25283(x25283, x16846, x25204);
  nand n25284(x25284, x25283, x25282);
  nand n25285(x25285, x16758, x25183);
  nand n25286(x25286, x16846, x25207);
  nand n25287(x25287, x25286, x25285);
  nand n25288(x25288, x16758, x25186);
  nand n25289(x25289, x16846, x25210);
  nand n25290(x25290, x25289, x25288);
  nand n25291(x25291, x16758, x25189);
  nand n25292(x25292, x16846, x25213);
  nand n25293(x25293, x25292, x25291);
  nand n25294(x25294, x16758, x25192);
  nand n25295(x25295, x16846, x25216);
  nand n25296(x25296, x25295, x25294);
  nand n25297(x25297, x16758, x25195);
  nand n25298(x25298, x16846, x25219);
  nand n25299(x25299, x25298, x25297);
  nand n25300(x25300, x16758, x25198);
  nand n25301(x25301, x16846, x25222);
  nand n25302(x25302, x25301, x25300);
  nand n25303(x25303, x16758, x25201);
  nand n25304(x25304, x16846, x25225);
  nand n25305(x25305, x25304, x25303);
  nand n25306(x25306, x16758, x25204);
  nand n25307(x25307, x16846, x25228);
  nand n25308(x25308, x25307, x25306);
  nand n25309(x25309, x16758, x25207);
  nand n25310(x25310, x16846, x25231);
  nand n25311(x25311, x25310, x25309);
  nand n25312(x25312, x16847, x83882);
  nand n25313(x25313, x16847, x83883);
  nand n25314(x25314, x16847, x83884);
  nand n25315(x25315, x16847, x83885);
  nand n25316(x25316, x16847, x83886);
  nand n25317(x25317, x16847, x83887);
  nand n25318(x25318, x16847, x83888);
  nand n25319(x25319, x16847, x83889);
  nand n25320(x25320, x16847, x25242);
  nand n25321(x25321, x16847, x25245);
  nand n25322(x25322, x16847, x25248);
  nand n25323(x25323, x16847, x25251);
  nand n25324(x25324, x16847, x25254);
  nand n25325(x25325, x16847, x25257);
  nand n25326(x25326, x16847, x25260);
  nand n25327(x25327, x16847, x25263);
  nand n25328(x25328, x16761, x83882);
  nand n25329(x25329, x16847, x25266);
  nand n25330(x25330, x25329, x25328);
  nand n25331(x25331, x16761, x83883);
  nand n25332(x25332, x16847, x25269);
  nand n25333(x25333, x25332, x25331);
  nand n25334(x25334, x16761, x83884);
  nand n25335(x25335, x16847, x25272);
  nand n25336(x25336, x25335, x25334);
  nand n25337(x25337, x16761, x83885);
  nand n25338(x25338, x16847, x25275);
  nand n25339(x25339, x25338, x25337);
  nand n25340(x25340, x16761, x83886);
  nand n25341(x25341, x16847, x25278);
  nand n25342(x25342, x25341, x25340);
  nand n25343(x25343, x16761, x83887);
  nand n25344(x25344, x16847, x25281);
  nand n25345(x25345, x25344, x25343);
  nand n25346(x25346, x16761, x83888);
  nand n25347(x25347, x16847, x25284);
  nand n25348(x25348, x25347, x25346);
  nand n25349(x25349, x16761, x83889);
  nand n25350(x25350, x16847, x25287);
  nand n25351(x25351, x25350, x25349);
  nand n25352(x25352, x16761, x25242);
  nand n25353(x25353, x16847, x25290);
  nand n25354(x25354, x25353, x25352);
  nand n25355(x25355, x16761, x25245);
  nand n25356(x25356, x16847, x25293);
  nand n25357(x25357, x25356, x25355);
  nand n25358(x25358, x16761, x25248);
  nand n25359(x25359, x16847, x25296);
  nand n25360(x25360, x25359, x25358);
  nand n25361(x25361, x16761, x25251);
  nand n25362(x25362, x16847, x25299);
  nand n25363(x25363, x25362, x25361);
  nand n25364(x25364, x16761, x25254);
  nand n25365(x25365, x16847, x25302);
  nand n25366(x25366, x25365, x25364);
  nand n25367(x25367, x16761, x25257);
  nand n25368(x25368, x16847, x25305);
  nand n25369(x25369, x25368, x25367);
  nand n25370(x25370, x16761, x25260);
  nand n25371(x25371, x16847, x25308);
  nand n25372(x25372, x25371, x25370);
  nand n25373(x25373, x16761, x25263);
  nand n25374(x25374, x16847, x25311);
  nand n25375(x25375, x25374, x25373);
  nand n25376(x25376, x24989, x17905);
  nand n25377(x25377, x24990, x17909);
  nand n25378(x25378, x24992, x17915);
  nand n25379(x25379, x24994, x17922);
  nand n25380(x25380, x24996, x17932);
  nand n25381(x25381, x24998, x17944);
  nand n25382(x25382, x25000, x17957);
  nand n25383(x25383, x25002, x17973);
  nand n25384(x25384, x25004, x17991);
  nand n25385(x25385, x25006, x18010);
  nand n25386(x25386, x25008, x18032);
  nand n25387(x25387, x25010, x18056);
  nand n25388(x25388, x25012, x18081);
  nand n25389(x25389, x25014, x18109);
  nand n25390(x25390, x25016, x18139);
  nand n25391(x25391, x25018, x18170);
  nand n25392(x25392, x25020, x18204);
  nand n25393(x25393, x25022, x18240);
  nand n25394(x25394, x25024, x18277);
  nand n25395(x25395, x25026, x18317);
  nand n25396(x25396, x25028, x18359);
  nand n25397(x25397, x25030, x18402);
  nand n25398(x25398, x25032, x18448);
  nand n25399(x25399, x25034, x18496);
  nand n25400(x25400, x25036, x18545);
  nand n25401(x25401, x25038, x18597);
  nand n25402(x25402, x25040, x18651);
  nand n25403(x25403, x25042, x18706);
  nand n25404(x25404, x25044, x18764);
  nand n25405(x25405, x25046, x18824);
  nand n25406(x25406, x25048, x18885);
  nand n25407(x25407, x16752, x25378);
  nand n25408(x25408, x16844, x25376);
  nand n25409(x25409, x25408, x25407);
  nand n25410(x25410, x16752, x25379);
  nand n25411(x25411, x16844, x25377);
  nand n25412(x25412, x25411, x25410);
  nand n25413(x25413, x16752, x25380);
  nand n25414(x25414, x16844, x25378);
  nand n25415(x25415, x25414, x25413);
  nand n25416(x25416, x16752, x25381);
  nand n25417(x25417, x16844, x25379);
  nand n25418(x25418, x25417, x25416);
  nand n25419(x25419, x16752, x25382);
  nand n25420(x25420, x16844, x25380);
  nand n25421(x25421, x25420, x25419);
  nand n25422(x25422, x16752, x25383);
  nand n25423(x25423, x16844, x25381);
  nand n25424(x25424, x25423, x25422);
  nand n25425(x25425, x16752, x25384);
  nand n25426(x25426, x16844, x25382);
  nand n25427(x25427, x25426, x25425);
  nand n25428(x25428, x16752, x25385);
  nand n25429(x25429, x16844, x25383);
  nand n25430(x25430, x25429, x25428);
  nand n25431(x25431, x16752, x25386);
  nand n25432(x25432, x16844, x25384);
  nand n25433(x25433, x25432, x25431);
  nand n25434(x25434, x16752, x25387);
  nand n25435(x25435, x16844, x25385);
  nand n25436(x25436, x25435, x25434);
  nand n25437(x25437, x16752, x25388);
  nand n25438(x25438, x16844, x25386);
  nand n25439(x25439, x25438, x25437);
  nand n25440(x25440, x16752, x25389);
  nand n25441(x25441, x16844, x25387);
  nand n25442(x25442, x25441, x25440);
  nand n25443(x25443, x16752, x25390);
  nand n25444(x25444, x16844, x25388);
  nand n25445(x25445, x25444, x25443);
  nand n25446(x25446, x16752, x25391);
  nand n25447(x25447, x16844, x25389);
  nand n25448(x25448, x25447, x25446);
  nand n25449(x25449, x16752, x25392);
  nand n25450(x25450, x16844, x25390);
  nand n25451(x25451, x25450, x25449);
  nand n25452(x25452, x16752, x25393);
  nand n25453(x25453, x16844, x25391);
  nand n25454(x25454, x25453, x25452);
  nand n25455(x25455, x16752, x25394);
  nand n25456(x25456, x16844, x25392);
  nand n25457(x25457, x25456, x25455);
  nand n25458(x25458, x16752, x25395);
  nand n25459(x25459, x16844, x25393);
  nand n25460(x25460, x25459, x25458);
  nand n25461(x25461, x16752, x25396);
  nand n25462(x25462, x16844, x25394);
  nand n25463(x25463, x25462, x25461);
  nand n25464(x25464, x16752, x25397);
  nand n25465(x25465, x16844, x25395);
  nand n25466(x25466, x25465, x25464);
  nand n25467(x25467, x16752, x25398);
  nand n25468(x25468, x16844, x25396);
  nand n25469(x25469, x25468, x25467);
  nand n25470(x25470, x16752, x25399);
  nand n25471(x25471, x16844, x25397);
  nand n25472(x25472, x25471, x25470);
  nand n25473(x25473, x16752, x25400);
  nand n25474(x25474, x16844, x25398);
  nand n25475(x25475, x25474, x25473);
  nand n25476(x25476, x16752, x25401);
  nand n25477(x25477, x16844, x25399);
  nand n25478(x25478, x25477, x25476);
  nand n25479(x25479, x16752, x25402);
  nand n25480(x25480, x16844, x25400);
  nand n25481(x25481, x25480, x25479);
  nand n25482(x25482, x16752, x25403);
  nand n25483(x25483, x16844, x25401);
  nand n25484(x25484, x25483, x25482);
  nand n25485(x25485, x16752, x25404);
  nand n25486(x25486, x16844, x25402);
  nand n25487(x25487, x25486, x25485);
  nand n25488(x25488, x16752, x25405);
  nand n25489(x25489, x16844, x25403);
  nand n25490(x25490, x25489, x25488);
  nand n25491(x25491, x16752, x25406);
  nand n25492(x25492, x16844, x25404);
  nand n25493(x25493, x25492, x25491);
  nand n25494(x25494, x16752, x83906);
  nand n25495(x25495, x16844, x25405);
  nand n25496(x25496, x25495, x25494);
  nand n25497(x25497, x16844, x25406);
  nand n25498(x25498, x16844, x83906);
  nand n25499(x25499, x16755, x25421);
  nand n25500(x25500, x16845, x25409);
  nand n25501(x25501, x25500, x25499);
  nand n25502(x25502, x16755, x25424);
  nand n25503(x25503, x16845, x25412);
  nand n25504(x25504, x25503, x25502);
  nand n25505(x25505, x16755, x25427);
  nand n25506(x25506, x16845, x25415);
  nand n25507(x25507, x25506, x25505);
  nand n25508(x25508, x16755, x25430);
  nand n25509(x25509, x16845, x25418);
  nand n25510(x25510, x25509, x25508);
  nand n25511(x25511, x16755, x25433);
  nand n25512(x25512, x16845, x25421);
  nand n25513(x25513, x25512, x25511);
  nand n25514(x25514, x16755, x25436);
  nand n25515(x25515, x16845, x25424);
  nand n25516(x25516, x25515, x25514);
  nand n25517(x25517, x16755, x25439);
  nand n25518(x25518, x16845, x25427);
  nand n25519(x25519, x25518, x25517);
  nand n25520(x25520, x16755, x25442);
  nand n25521(x25521, x16845, x25430);
  nand n25522(x25522, x25521, x25520);
  nand n25523(x25523, x16755, x25445);
  nand n25524(x25524, x16845, x25433);
  nand n25525(x25525, x25524, x25523);
  nand n25526(x25526, x16755, x25448);
  nand n25527(x25527, x16845, x25436);
  nand n25528(x25528, x25527, x25526);
  nand n25529(x25529, x16755, x25451);
  nand n25530(x25530, x16845, x25439);
  nand n25531(x25531, x25530, x25529);
  nand n25532(x25532, x16755, x25454);
  nand n25533(x25533, x16845, x25442);
  nand n25534(x25534, x25533, x25532);
  nand n25535(x25535, x16755, x25457);
  nand n25536(x25536, x16845, x25445);
  nand n25537(x25537, x25536, x25535);
  nand n25538(x25538, x16755, x25460);
  nand n25539(x25539, x16845, x25448);
  nand n25540(x25540, x25539, x25538);
  nand n25541(x25541, x16755, x25463);
  nand n25542(x25542, x16845, x25451);
  nand n25543(x25543, x25542, x25541);
  nand n25544(x25544, x16755, x25466);
  nand n25545(x25545, x16845, x25454);
  nand n25546(x25546, x25545, x25544);
  nand n25547(x25547, x16755, x25469);
  nand n25548(x25548, x16845, x25457);
  nand n25549(x25549, x25548, x25547);
  nand n25550(x25550, x16755, x25472);
  nand n25551(x25551, x16845, x25460);
  nand n25552(x25552, x25551, x25550);
  nand n25553(x25553, x16755, x25475);
  nand n25554(x25554, x16845, x25463);
  nand n25555(x25555, x25554, x25553);
  nand n25556(x25556, x16755, x25478);
  nand n25557(x25557, x16845, x25466);
  nand n25558(x25558, x25557, x25556);
  nand n25559(x25559, x16755, x25481);
  nand n25560(x25560, x16845, x25469);
  nand n25561(x25561, x25560, x25559);
  nand n25562(x25562, x16755, x25484);
  nand n25563(x25563, x16845, x25472);
  nand n25564(x25564, x25563, x25562);
  nand n25565(x25565, x16755, x25487);
  nand n25566(x25566, x16845, x25475);
  nand n25567(x25567, x25566, x25565);
  nand n25568(x25568, x16755, x25490);
  nand n25569(x25569, x16845, x25478);
  nand n25570(x25570, x25569, x25568);
  nand n25571(x25571, x16755, x25493);
  nand n25572(x25572, x16845, x25481);
  nand n25573(x25573, x25572, x25571);
  nand n25574(x25574, x16755, x25496);
  nand n25575(x25575, x16845, x25484);
  nand n25576(x25576, x25575, x25574);
  nand n25577(x25577, x16755, x83907);
  nand n25578(x25578, x16845, x25487);
  nand n25579(x25579, x25578, x25577);
  nand n25580(x25580, x16755, x83908);
  nand n25581(x25581, x16845, x25490);
  nand n25582(x25582, x25581, x25580);
  nand n25583(x25583, x16845, x25493);
  nand n25584(x25584, x16845, x25496);
  nand n25585(x25585, x16845, x83907);
  nand n25586(x25586, x16845, x83908);
  nand n25587(x25587, x16758, x25525);
  nand n25588(x25588, x16846, x25501);
  nand n25589(x25589, x25588, x25587);
  nand n25590(x25590, x16758, x25528);
  nand n25591(x25591, x16846, x25504);
  nand n25592(x25592, x25591, x25590);
  nand n25593(x25593, x16758, x25531);
  nand n25594(x25594, x16846, x25507);
  nand n25595(x25595, x25594, x25593);
  nand n25596(x25596, x16758, x25534);
  nand n25597(x25597, x16846, x25510);
  nand n25598(x25598, x25597, x25596);
  nand n25599(x25599, x16758, x25537);
  nand n25600(x25600, x16846, x25513);
  nand n25601(x25601, x25600, x25599);
  nand n25602(x25602, x16758, x25540);
  nand n25603(x25603, x16846, x25516);
  nand n25604(x25604, x25603, x25602);
  nand n25605(x25605, x16758, x25543);
  nand n25606(x25606, x16846, x25519);
  nand n25607(x25607, x25606, x25605);
  nand n25608(x25608, x16758, x25546);
  nand n25609(x25609, x16846, x25522);
  nand n25610(x25610, x25609, x25608);
  nand n25611(x25611, x16758, x25549);
  nand n25612(x25612, x16846, x25525);
  nand n25613(x25613, x25612, x25611);
  nand n25614(x25614, x16758, x25552);
  nand n25615(x25615, x16846, x25528);
  nand n25616(x25616, x25615, x25614);
  nand n25617(x25617, x16758, x25555);
  nand n25618(x25618, x16846, x25531);
  nand n25619(x25619, x25618, x25617);
  nand n25620(x25620, x16758, x25558);
  nand n25621(x25621, x16846, x25534);
  nand n25622(x25622, x25621, x25620);
  nand n25623(x25623, x16758, x25561);
  nand n25624(x25624, x16846, x25537);
  nand n25625(x25625, x25624, x25623);
  nand n25626(x25626, x16758, x25564);
  nand n25627(x25627, x16846, x25540);
  nand n25628(x25628, x25627, x25626);
  nand n25629(x25629, x16758, x25567);
  nand n25630(x25630, x16846, x25543);
  nand n25631(x25631, x25630, x25629);
  nand n25632(x25632, x16758, x25570);
  nand n25633(x25633, x16846, x25546);
  nand n25634(x25634, x25633, x25632);
  nand n25635(x25635, x16758, x25573);
  nand n25636(x25636, x16846, x25549);
  nand n25637(x25637, x25636, x25635);
  nand n25638(x25638, x16758, x25576);
  nand n25639(x25639, x16846, x25552);
  nand n25640(x25640, x25639, x25638);
  nand n25641(x25641, x16758, x25579);
  nand n25642(x25642, x16846, x25555);
  nand n25643(x25643, x25642, x25641);
  nand n25644(x25644, x16758, x25582);
  nand n25645(x25645, x16846, x25558);
  nand n25646(x25646, x25645, x25644);
  nand n25647(x25647, x16758, x83909);
  nand n25648(x25648, x16846, x25561);
  nand n25649(x25649, x25648, x25647);
  nand n25650(x25650, x16758, x83910);
  nand n25651(x25651, x16846, x25564);
  nand n25652(x25652, x25651, x25650);
  nand n25653(x25653, x16758, x83911);
  nand n25654(x25654, x16846, x25567);
  nand n25655(x25655, x25654, x25653);
  nand n25656(x25656, x16758, x83912);
  nand n25657(x25657, x16846, x25570);
  nand n25658(x25658, x25657, x25656);
  nand n25659(x25659, x16846, x25573);
  nand n25660(x25660, x16846, x25576);
  nand n25661(x25661, x16846, x25579);
  nand n25662(x25662, x16846, x25582);
  nand n25663(x25663, x16846, x83909);
  nand n25664(x25664, x16846, x83910);
  nand n25665(x25665, x16846, x83911);
  nand n25666(x25666, x16846, x83912);
  nand n25667(x25667, x16761, x25637);
  nand n25668(x25668, x16847, x25589);
  nand n25669(x25669, x25668, x25667);
  nand n25670(x25670, x16761, x25640);
  nand n25671(x25671, x16847, x25592);
  nand n25672(x25672, x25671, x25670);
  nand n25673(x25673, x16761, x25643);
  nand n25674(x25674, x16847, x25595);
  nand n25675(x25675, x25674, x25673);
  nand n25676(x25676, x16761, x25646);
  nand n25677(x25677, x16847, x25598);
  nand n25678(x25678, x25677, x25676);
  nand n25679(x25679, x16761, x25649);
  nand n25680(x25680, x16847, x25601);
  nand n25681(x25681, x25680, x25679);
  nand n25682(x25682, x16761, x25652);
  nand n25683(x25683, x16847, x25604);
  nand n25684(x25684, x25683, x25682);
  nand n25685(x25685, x16761, x25655);
  nand n25686(x25686, x16847, x25607);
  nand n25687(x25687, x25686, x25685);
  nand n25688(x25688, x16761, x25658);
  nand n25689(x25689, x16847, x25610);
  nand n25690(x25690, x25689, x25688);
  nand n25691(x25691, x16761, x83913);
  nand n25692(x25692, x16847, x25613);
  nand n25693(x25693, x25692, x25691);
  nand n25694(x25694, x16761, x83914);
  nand n25695(x25695, x16847, x25616);
  nand n25696(x25696, x25695, x25694);
  nand n25697(x25697, x16761, x83915);
  nand n25698(x25698, x16847, x25619);
  nand n25699(x25699, x25698, x25697);
  nand n25700(x25700, x16761, x83916);
  nand n25701(x25701, x16847, x25622);
  nand n25702(x25702, x25701, x25700);
  nand n25703(x25703, x16761, x83917);
  nand n25704(x25704, x16847, x25625);
  nand n25705(x25705, x25704, x25703);
  nand n25706(x25706, x16761, x83918);
  nand n25707(x25707, x16847, x25628);
  nand n25708(x25708, x25707, x25706);
  nand n25709(x25709, x16761, x83919);
  nand n25710(x25710, x16847, x25631);
  nand n25711(x25711, x25710, x25709);
  nand n25712(x25712, x16761, x83920);
  nand n25713(x25713, x16847, x25634);
  nand n25714(x25714, x25713, x25712);
  nand n25715(x25715, x16847, x25637);
  nand n25716(x25716, x16847, x25640);
  nand n25717(x25717, x16847, x25643);
  nand n25718(x25718, x16847, x25646);
  nand n25719(x25719, x16847, x25649);
  nand n25720(x25720, x16847, x25652);
  nand n25721(x25721, x16847, x25655);
  nand n25722(x25722, x16847, x25658);
  nand n25723(x25723, x16847, x83913);
  nand n25724(x25724, x16847, x83914);
  nand n25725(x25725, x16847, x83915);
  nand n25726(x25726, x16847, x83916);
  nand n25727(x25727, x16847, x83917);
  nand n25728(x25728, x16847, x83918);
  nand n25729(x25729, x16847, x83919);
  nand n25730(x25730, x16847, x83920);
  nand n25731(x25731, x71977, x16749);
  nand n25732(x25732, x16876, x71642);
  nand n25733(x25733, x71977, x71642);
  nand n25734(x25734, x16876, x25669);
  nand n25735(x25735, x25734, x25733);
  nand n25736(x25736, x71977, x83890);
  nand n25737(x25737, x16876, x24860);
  nand n25738(x25738, x71977, x17748);
  nand n25739(x25739, x16876, x17748);
  nand n25740(x25740, x25739, x25738);
  nand n25741(x25741, x71977, x24926);
  nand n25742(x25742, x16876, x24893);
  nand n25743(x25743, x25742, x25741);
  nand n25744(x25744, x71977, x24860);
  nand n25745(x25745, x25734, x25744);
  nand n25746(x25746, x16876, x16974);
  nand n25747(x25747, x25746, x25744);
  nand n25748(x25748, x71977, x72047);
  nand n25750(x25750, x25749, x83937);
  nand n25751(x25751, x25749, x83938);
  nand n25752(x25752, x71982, x25735);
  nand n25753(x25753, x25749, x83939);
  nand n25754(x25754, x25753, x25752);
  nand n25755(x25755, x71982, x83940);
  nand n25756(x25756, x25749, x25740);
  nand n25757(x25757, x25756, x25755);
  nand n25758(x25758, x71982, x25743);
  nand n25759(x25759, x25749, x25745);
  nand n25760(x25760, x25759, x25758);
  nand n25761(x25761, x71982, x83939);
  nand n25762(x25762, x25749, x83940);
  nand n25763(x25763, x25762, x25761);
  nand n25764(x25764, x71982, x25740);
  nand n25765(x25765, x25749, x25743);
  nand n25766(x25766, x25765, x25764);
  nand n25767(x25767, x71982, x25747);
  nand n25768(x25768, x25749, x83941);
  nand n25769(x25769, x25768, x25767);
  nand n25770(x25770, x71987, x83942);
  nand n25771(x25771, x71987, x83943);
  nand n25773(x25773, x25772, x25754);
  nand n25774(x25774, x25773, x25771);
  nand n25775(x25775, x71987, x25757);
  nand n25776(x25776, x25772, x25760);
  nand n25777(x25777, x25776, x25775);
  nand n25778(x25778, x71987, x25763);
  nand n25779(x25779, x25772, x25766);
  nand n25780(x25780, x25779, x25778);
  nand n25781(x25781, x71987, x25769);
  nand n25783(x25783, x25782, x83944);
  nand n25784(x25784, x71992, x25774);
  nand n25785(x25785, x25782, x25777);
  nand n25786(x25786, x25785, x25784);
  nand n25787(x25787, x71992, x25780);
  nand n25788(x25788, x25782, x83945);
  nand n25789(x25789, x25788, x25787);
  nand n25791(x25791, x25790, x83946);
  nand n25792(x25792, x71997, x25786);
  nand n25793(x25793, x25790, x25789);
  nand n25794(x25794, x25793, x25792);
  nand n25795(x25795, x72002, x83947);
  nand n25797(x25797, x25796, x25794);
  nand n25798(x25798, x25797, x25795);
  nand n25799(x25799, x71977, x16752);
  nand n25800(x25800, x16876, x71647);
  nand n25801(x25801, x71977, x71647);
  nand n25802(x25802, x16876, x25672);
  nand n25803(x25803, x25802, x25801);
  nand n25804(x25804, x71977, x83891);
  nand n25805(x25805, x16876, x83843);
  nand n25806(x25806, x71977, x17753);
  nand n25807(x25807, x16876, x17753);
  nand n25808(x25808, x25807, x25806);
  nand n25809(x25809, x71977, x24928);
  nand n25810(x25810, x16876, x24894);
  nand n25811(x25811, x25810, x25809);
  nand n25812(x25812, x71977, x17912);
  nand n25813(x25813, x25802, x25812);
  nand n25814(x25814, x16876, x16980);
  nand n25815(x25815, x25814, x25812);
  nand n25816(x25816, x71977, x24739);
  nand n25817(x25817, x25749, x83948);
  nand n25818(x25818, x25749, x83949);
  nand n25819(x25819, x71982, x25803);
  nand n25820(x25820, x25749, x83950);
  nand n25821(x25821, x25820, x25819);
  nand n25822(x25822, x71982, x83951);
  nand n25823(x25823, x25749, x25808);
  nand n25824(x25824, x25823, x25822);
  nand n25825(x25825, x71982, x25811);
  nand n25826(x25826, x25749, x25813);
  nand n25827(x25827, x25826, x25825);
  nand n25828(x25828, x71982, x83950);
  nand n25829(x25829, x25749, x83951);
  nand n25830(x25830, x25829, x25828);
  nand n25831(x25831, x71982, x25808);
  nand n25832(x25832, x25749, x25811);
  nand n25833(x25833, x25832, x25831);
  nand n25834(x25834, x71982, x25815);
  nand n25835(x25835, x25749, x83952);
  nand n25836(x25836, x25835, x25834);
  nand n25837(x25837, x71987, x83953);
  nand n25838(x25838, x71987, x83954);
  nand n25839(x25839, x25772, x25821);
  nand n25840(x25840, x25839, x25838);
  nand n25841(x25841, x71987, x25824);
  nand n25842(x25842, x25772, x25827);
  nand n25843(x25843, x25842, x25841);
  nand n25844(x25844, x71987, x25830);
  nand n25845(x25845, x25772, x25833);
  nand n25846(x25846, x25845, x25844);
  nand n25847(x25847, x71987, x25836);
  nand n25848(x25848, x25782, x83955);
  nand n25849(x25849, x71992, x25840);
  nand n25850(x25850, x25782, x25843);
  nand n25851(x25851, x25850, x25849);
  nand n25852(x25852, x71992, x25846);
  nand n25853(x25853, x25782, x83956);
  nand n25854(x25854, x25853, x25852);
  nand n25855(x25855, x25790, x83957);
  nand n25856(x25856, x71997, x25851);
  nand n25857(x25857, x25790, x25854);
  nand n25858(x25858, x25857, x25856);
  nand n25859(x25859, x72002, x83958);
  nand n25860(x25860, x25796, x25858);
  nand n25861(x25861, x25860, x25859);
  nand n25862(x25862, x71977, x16755);
  nand n25863(x25863, x16876, x71652);
  nand n25864(x25864, x71977, x71652);
  nand n25865(x25865, x16876, x25675);
  nand n25866(x25866, x25865, x25864);
  nand n25867(x25867, x71977, x83892);
  nand n25868(x25868, x16876, x83844);
  nand n25869(x25869, x71977, x17758);
  nand n25870(x25870, x16876, x17758);
  nand n25871(x25871, x25870, x25869);
  nand n25872(x25872, x71977, x24930);
  nand n25873(x25873, x16876, x24895);
  nand n25874(x25874, x25873, x25872);
  nand n25875(x25875, x71977, x17927);
  nand n25876(x25876, x25865, x25875);
  nand n25877(x25877, x16876, x16986);
  nand n25878(x25878, x25877, x25875);
  nand n25879(x25879, x71977, x24743);
  nand n25880(x25880, x25749, x83959);
  nand n25881(x25881, x25749, x83960);
  nand n25882(x25882, x71982, x25866);
  nand n25883(x25883, x25749, x83961);
  nand n25884(x25884, x25883, x25882);
  nand n25885(x25885, x71982, x83962);
  nand n25886(x25886, x25749, x25871);
  nand n25887(x25887, x25886, x25885);
  nand n25888(x25888, x71982, x25874);
  nand n25889(x25889, x25749, x25876);
  nand n25890(x25890, x25889, x25888);
  nand n25891(x25891, x71982, x83961);
  nand n25892(x25892, x25749, x83962);
  nand n25893(x25893, x25892, x25891);
  nand n25894(x25894, x71982, x25871);
  nand n25895(x25895, x25749, x25874);
  nand n25896(x25896, x25895, x25894);
  nand n25897(x25897, x71982, x25878);
  nand n25898(x25898, x25749, x83963);
  nand n25899(x25899, x25898, x25897);
  nand n25900(x25900, x71987, x83964);
  nand n25901(x25901, x71987, x83965);
  nand n25902(x25902, x25772, x25884);
  nand n25903(x25903, x25902, x25901);
  nand n25904(x25904, x71987, x25887);
  nand n25905(x25905, x25772, x25890);
  nand n25906(x25906, x25905, x25904);
  nand n25907(x25907, x71987, x25893);
  nand n25908(x25908, x25772, x25896);
  nand n25909(x25909, x25908, x25907);
  nand n25910(x25910, x71987, x25899);
  nand n25911(x25911, x25782, x83966);
  nand n25912(x25912, x71992, x25903);
  nand n25913(x25913, x25782, x25906);
  nand n25914(x25914, x25913, x25912);
  nand n25915(x25915, x71992, x25909);
  nand n25916(x25916, x25782, x83967);
  nand n25917(x25917, x25916, x25915);
  nand n25918(x25918, x25790, x83968);
  nand n25919(x25919, x71997, x25914);
  nand n25920(x25920, x25790, x25917);
  nand n25921(x25921, x25920, x25919);
  nand n25922(x25922, x72002, x83969);
  nand n25923(x25923, x25796, x25921);
  nand n25924(x25924, x25923, x25922);
  nand n25925(x25925, x71977, x16758);
  nand n25926(x25926, x16876, x71657);
  nand n25927(x25927, x71977, x71657);
  nand n25928(x25928, x16876, x25678);
  nand n25929(x25929, x25928, x25927);
  nand n25930(x25930, x71977, x83893);
  nand n25931(x25931, x16876, x83845);
  nand n25932(x25932, x71977, x17763);
  nand n25933(x25933, x16876, x17763);
  nand n25934(x25934, x25933, x25932);
  nand n25935(x25935, x71977, x24932);
  nand n25936(x25936, x16876, x24896);
  nand n25937(x25937, x25936, x25935);
  nand n25938(x25938, x71977, x17951);
  nand n25939(x25939, x25928, x25938);
  nand n25940(x25940, x16876, x16992);
  nand n25941(x25941, x25940, x25938);
  nand n25942(x25942, x71977, x24747);
  nand n25943(x25943, x25749, x83970);
  nand n25944(x25944, x25749, x83971);
  nand n25945(x25945, x71982, x25929);
  nand n25946(x25946, x25749, x83972);
  nand n25947(x25947, x25946, x25945);
  nand n25948(x25948, x71982, x83973);
  nand n25949(x25949, x25749, x25934);
  nand n25950(x25950, x25949, x25948);
  nand n25951(x25951, x71982, x25937);
  nand n25952(x25952, x25749, x25939);
  nand n25953(x25953, x25952, x25951);
  nand n25954(x25954, x71982, x83972);
  nand n25955(x25955, x25749, x83973);
  nand n25956(x25956, x25955, x25954);
  nand n25957(x25957, x71982, x25934);
  nand n25958(x25958, x25749, x25937);
  nand n25959(x25959, x25958, x25957);
  nand n25960(x25960, x71982, x25941);
  nand n25961(x25961, x25749, x83974);
  nand n25962(x25962, x25961, x25960);
  nand n25963(x25963, x71987, x83975);
  nand n25964(x25964, x71987, x83976);
  nand n25965(x25965, x25772, x25947);
  nand n25966(x25966, x25965, x25964);
  nand n25967(x25967, x71987, x25950);
  nand n25968(x25968, x25772, x25953);
  nand n25969(x25969, x25968, x25967);
  nand n25970(x25970, x71987, x25956);
  nand n25971(x25971, x25772, x25959);
  nand n25972(x25972, x25971, x25970);
  nand n25973(x25973, x71987, x25962);
  nand n25974(x25974, x25782, x83977);
  nand n25975(x25975, x71992, x25966);
  nand n25976(x25976, x25782, x25969);
  nand n25977(x25977, x25976, x25975);
  nand n25978(x25978, x71992, x25972);
  nand n25979(x25979, x25782, x83978);
  nand n25980(x25980, x25979, x25978);
  nand n25981(x25981, x25790, x83979);
  nand n25982(x25982, x71997, x25977);
  nand n25983(x25983, x25790, x25980);
  nand n25984(x25984, x25983, x25982);
  nand n25985(x25985, x72002, x83980);
  nand n25986(x25986, x25796, x25984);
  nand n25987(x25987, x25986, x25985);
  nand n25988(x25988, x71977, x16761);
  nand n25989(x25989, x16876, x71662);
  nand n25990(x25990, x71977, x71662);
  nand n25991(x25991, x16876, x25681);
  nand n25992(x25992, x25991, x25990);
  nand n25993(x25993, x71977, x83894);
  nand n25994(x25994, x16876, x83846);
  nand n25995(x25995, x71977, x17768);
  nand n25996(x25996, x16876, x17768);
  nand n25997(x25997, x25996, x25995);
  nand n25998(x25998, x71977, x24934);
  nand n25999(x25999, x16876, x24897);
  nand n26000(x26000, x25999, x25998);
  nand n26001(x26001, x71977, x17982);
  nand n26002(x26002, x25991, x26001);
  nand n26003(x26003, x16876, x16998);
  nand n26004(x26004, x26003, x26001);
  nand n26005(x26005, x71977, x24751);
  nand n26006(x26006, x25749, x83981);
  nand n26007(x26007, x25749, x83982);
  nand n26008(x26008, x71982, x25992);
  nand n26009(x26009, x25749, x83983);
  nand n26010(x26010, x26009, x26008);
  nand n26011(x26011, x71982, x83984);
  nand n26012(x26012, x25749, x25997);
  nand n26013(x26013, x26012, x26011);
  nand n26014(x26014, x71982, x26000);
  nand n26015(x26015, x25749, x26002);
  nand n26016(x26016, x26015, x26014);
  nand n26017(x26017, x71982, x83983);
  nand n26018(x26018, x25749, x83984);
  nand n26019(x26019, x26018, x26017);
  nand n26020(x26020, x71982, x25997);
  nand n26021(x26021, x25749, x26000);
  nand n26022(x26022, x26021, x26020);
  nand n26023(x26023, x71982, x26004);
  nand n26024(x26024, x25749, x83985);
  nand n26025(x26025, x26024, x26023);
  nand n26026(x26026, x71987, x83986);
  nand n26027(x26027, x71987, x83987);
  nand n26028(x26028, x25772, x26010);
  nand n26029(x26029, x26028, x26027);
  nand n26030(x26030, x71987, x26013);
  nand n26031(x26031, x25772, x26016);
  nand n26032(x26032, x26031, x26030);
  nand n26033(x26033, x71987, x26019);
  nand n26034(x26034, x25772, x26022);
  nand n26035(x26035, x26034, x26033);
  nand n26036(x26036, x71987, x26025);
  nand n26037(x26037, x25782, x83988);
  nand n26038(x26038, x71992, x26029);
  nand n26039(x26039, x25782, x26032);
  nand n26040(x26040, x26039, x26038);
  nand n26041(x26041, x71992, x26035);
  nand n26042(x26042, x25782, x83989);
  nand n26043(x26043, x26042, x26041);
  nand n26044(x26044, x25790, x83990);
  nand n26045(x26045, x71997, x26040);
  nand n26046(x26046, x25790, x26043);
  nand n26047(x26047, x26046, x26045);
  nand n26048(x26048, x72002, x83991);
  nand n26049(x26049, x25796, x26047);
  nand n26050(x26050, x26049, x26048);
  nand n26051(x26051, x71977, x16764);
  nand n26052(x26052, x16876, x71667);
  nand n26053(x26053, x71977, x71667);
  nand n26054(x26054, x16876, x25684);
  nand n26055(x26055, x26054, x26053);
  nand n26056(x26056, x71977, x83895);
  nand n26057(x26057, x16876, x83847);
  nand n26058(x26058, x71977, x17773);
  nand n26059(x26059, x16876, x17773);
  nand n26060(x26060, x26059, x26058);
  nand n26061(x26061, x71977, x24936);
  nand n26062(x26062, x16876, x24898);
  nand n26063(x26063, x26062, x26061);
  nand n26064(x26064, x71977, x18021);
  nand n26065(x26065, x26054, x26064);
  nand n26066(x26066, x16876, x17004);
  nand n26067(x26067, x26066, x26064);
  nand n26068(x26068, x71977, x24755);
  nand n26069(x26069, x25749, x83992);
  nand n26070(x26070, x25749, x83993);
  nand n26071(x26071, x71982, x26055);
  nand n26072(x26072, x25749, x83994);
  nand n26073(x26073, x26072, x26071);
  nand n26074(x26074, x71982, x83995);
  nand n26075(x26075, x25749, x26060);
  nand n26076(x26076, x26075, x26074);
  nand n26077(x26077, x71982, x26063);
  nand n26078(x26078, x25749, x26065);
  nand n26079(x26079, x26078, x26077);
  nand n26080(x26080, x71982, x83994);
  nand n26081(x26081, x25749, x83995);
  nand n26082(x26082, x26081, x26080);
  nand n26083(x26083, x71982, x26060);
  nand n26084(x26084, x25749, x26063);
  nand n26085(x26085, x26084, x26083);
  nand n26086(x26086, x71982, x26067);
  nand n26087(x26087, x25749, x83996);
  nand n26088(x26088, x26087, x26086);
  nand n26089(x26089, x71987, x83997);
  nand n26090(x26090, x71987, x83998);
  nand n26091(x26091, x25772, x26073);
  nand n26092(x26092, x26091, x26090);
  nand n26093(x26093, x71987, x26076);
  nand n26094(x26094, x25772, x26079);
  nand n26095(x26095, x26094, x26093);
  nand n26096(x26096, x71987, x26082);
  nand n26097(x26097, x25772, x26085);
  nand n26098(x26098, x26097, x26096);
  nand n26099(x26099, x71987, x26088);
  nand n26100(x26100, x25782, x83999);
  nand n26101(x26101, x71992, x26092);
  nand n26102(x26102, x25782, x26095);
  nand n26103(x26103, x26102, x26101);
  nand n26104(x26104, x71992, x26098);
  nand n26105(x26105, x25782, x84000);
  nand n26106(x26106, x26105, x26104);
  nand n26107(x26107, x25790, x84001);
  nand n26108(x26108, x71997, x26103);
  nand n26109(x26109, x25790, x26106);
  nand n26110(x26110, x26109, x26108);
  nand n26111(x26111, x72002, x84002);
  nand n26112(x26112, x25796, x26110);
  nand n26113(x26113, x26112, x26111);
  nand n26114(x26114, x71977, x16767);
  nand n26115(x26115, x16876, x71672);
  nand n26116(x26116, x71977, x71672);
  nand n26117(x26117, x16876, x25687);
  nand n26118(x26118, x26117, x26116);
  nand n26119(x26119, x71977, x83896);
  nand n26120(x26120, x16876, x24403);
  nand n26121(x26121, x71977, x17778);
  nand n26122(x26122, x16876, x17778);
  nand n26123(x26123, x26122, x26121);
  nand n26124(x26124, x71977, x24938);
  nand n26125(x26125, x16876, x24899);
  nand n26126(x26126, x26125, x26124);
  nand n26127(x26127, x71977, x18069);
  nand n26128(x26128, x26117, x26127);
  nand n26129(x26129, x16876, x17010);
  nand n26130(x26130, x26129, x26127);
  nand n26131(x26131, x71977, x24759);
  nand n26132(x26132, x25749, x84003);
  nand n26133(x26133, x25749, x84004);
  nand n26134(x26134, x71982, x26118);
  nand n26135(x26135, x25749, x84005);
  nand n26136(x26136, x26135, x26134);
  nand n26137(x26137, x71982, x84006);
  nand n26138(x26138, x25749, x26123);
  nand n26139(x26139, x26138, x26137);
  nand n26140(x26140, x71982, x26126);
  nand n26141(x26141, x25749, x26128);
  nand n26142(x26142, x26141, x26140);
  nand n26143(x26143, x71982, x84005);
  nand n26144(x26144, x25749, x84006);
  nand n26145(x26145, x26144, x26143);
  nand n26146(x26146, x71982, x26123);
  nand n26147(x26147, x25749, x26126);
  nand n26148(x26148, x26147, x26146);
  nand n26149(x26149, x71982, x26130);
  nand n26150(x26150, x25749, x84007);
  nand n26151(x26151, x26150, x26149);
  nand n26152(x26152, x71987, x84008);
  nand n26153(x26153, x71987, x84009);
  nand n26154(x26154, x25772, x26136);
  nand n26155(x26155, x26154, x26153);
  nand n26156(x26156, x71987, x26139);
  nand n26157(x26157, x25772, x26142);
  nand n26158(x26158, x26157, x26156);
  nand n26159(x26159, x71987, x26145);
  nand n26160(x26160, x25772, x26148);
  nand n26161(x26161, x26160, x26159);
  nand n26162(x26162, x71987, x26151);
  nand n26163(x26163, x25782, x84010);
  nand n26164(x26164, x71992, x26155);
  nand n26165(x26165, x25782, x26158);
  nand n26166(x26166, x26165, x26164);
  nand n26167(x26167, x71992, x26161);
  nand n26168(x26168, x25782, x84011);
  nand n26169(x26169, x26168, x26167);
  nand n26170(x26170, x25790, x84012);
  nand n26171(x26171, x71997, x26166);
  nand n26172(x26172, x25790, x26169);
  nand n26173(x26173, x26172, x26171);
  nand n26174(x26174, x72002, x84013);
  nand n26175(x26175, x25796, x26173);
  nand n26176(x26176, x26175, x26174);
  nand n26177(x26177, x71977, x16770);
  nand n26178(x26178, x16876, x71677);
  nand n26179(x26179, x71977, x71677);
  nand n26180(x26180, x16876, x25690);
  nand n26181(x26181, x26180, x26179);
  nand n26182(x26182, x71977, x83897);
  nand n26183(x26183, x16876, x24407);
  nand n26184(x26184, x71977, x17783);
  nand n26185(x26185, x16876, x17783);
  nand n26186(x26186, x26185, x26184);
  nand n26187(x26187, x71977, x24940);
  nand n26188(x26188, x16876, x24900);
  nand n26189(x26189, x26188, x26187);
  nand n26190(x26190, x71977, x18124);
  nand n26191(x26191, x26180, x26190);
  nand n26192(x26192, x16876, x17016);
  nand n26193(x26193, x26192, x26190);
  nand n26194(x26194, x71977, x24763);
  nand n26195(x26195, x25749, x84014);
  nand n26196(x26196, x25749, x84015);
  nand n26197(x26197, x71982, x26181);
  nand n26198(x26198, x25749, x84016);
  nand n26199(x26199, x26198, x26197);
  nand n26200(x26200, x71982, x84017);
  nand n26201(x26201, x25749, x26186);
  nand n26202(x26202, x26201, x26200);
  nand n26203(x26203, x71982, x26189);
  nand n26204(x26204, x25749, x26191);
  nand n26205(x26205, x26204, x26203);
  nand n26206(x26206, x71982, x84016);
  nand n26207(x26207, x25749, x84017);
  nand n26208(x26208, x26207, x26206);
  nand n26209(x26209, x71982, x26186);
  nand n26210(x26210, x25749, x26189);
  nand n26211(x26211, x26210, x26209);
  nand n26212(x26212, x71982, x26193);
  nand n26213(x26213, x25749, x84018);
  nand n26214(x26214, x26213, x26212);
  nand n26215(x26215, x71987, x84019);
  nand n26216(x26216, x71987, x84020);
  nand n26217(x26217, x25772, x26199);
  nand n26218(x26218, x26217, x26216);
  nand n26219(x26219, x71987, x26202);
  nand n26220(x26220, x25772, x26205);
  nand n26221(x26221, x26220, x26219);
  nand n26222(x26222, x71987, x26208);
  nand n26223(x26223, x25772, x26211);
  nand n26224(x26224, x26223, x26222);
  nand n26225(x26225, x71987, x26214);
  nand n26226(x26226, x25782, x84021);
  nand n26227(x26227, x71992, x26218);
  nand n26228(x26228, x25782, x26221);
  nand n26229(x26229, x26228, x26227);
  nand n26230(x26230, x71992, x26224);
  nand n26231(x26231, x25782, x84022);
  nand n26232(x26232, x26231, x26230);
  nand n26233(x26233, x25790, x84023);
  nand n26234(x26234, x71997, x26229);
  nand n26235(x26235, x25790, x26232);
  nand n26236(x26236, x26235, x26234);
  nand n26237(x26237, x72002, x84024);
  nand n26238(x26238, x25796, x26236);
  nand n26239(x26239, x26238, x26237);
  nand n26240(x26240, x71977, x16773);
  nand n26241(x26241, x16876, x71682);
  nand n26242(x26242, x71977, x71682);
  nand n26243(x26243, x16876, x25693);
  nand n26244(x26244, x26243, x26242);
  nand n26245(x26245, x71977, x83898);
  nand n26246(x26246, x16876, x24411);
  nand n26247(x26247, x71977, x17788);
  nand n26248(x26248, x16876, x17788);
  nand n26249(x26249, x26248, x26247);
  nand n26250(x26250, x71977, x24942);
  nand n26251(x26251, x16876, x24901);
  nand n26252(x26252, x26251, x26250);
  nand n26253(x26253, x71977, x18187);
  nand n26254(x26254, x26243, x26253);
  nand n26255(x26255, x16876, x17022);
  nand n26256(x26256, x26255, x26253);
  nand n26257(x26257, x71977, x24767);
  nand n26258(x26258, x25749, x84025);
  nand n26259(x26259, x25749, x84026);
  nand n26260(x26260, x71982, x26244);
  nand n26261(x26261, x25749, x84027);
  nand n26262(x26262, x26261, x26260);
  nand n26263(x26263, x71982, x84028);
  nand n26264(x26264, x25749, x26249);
  nand n26265(x26265, x26264, x26263);
  nand n26266(x26266, x71982, x26252);
  nand n26267(x26267, x25749, x26254);
  nand n26268(x26268, x26267, x26266);
  nand n26269(x26269, x71982, x84027);
  nand n26270(x26270, x25749, x84028);
  nand n26271(x26271, x26270, x26269);
  nand n26272(x26272, x71982, x26249);
  nand n26273(x26273, x25749, x26252);
  nand n26274(x26274, x26273, x26272);
  nand n26275(x26275, x71982, x26256);
  nand n26276(x26276, x25749, x84029);
  nand n26277(x26277, x26276, x26275);
  nand n26278(x26278, x71987, x84030);
  nand n26279(x26279, x71987, x84031);
  nand n26280(x26280, x25772, x26262);
  nand n26281(x26281, x26280, x26279);
  nand n26282(x26282, x71987, x26265);
  nand n26283(x26283, x25772, x26268);
  nand n26284(x26284, x26283, x26282);
  nand n26285(x26285, x71987, x26271);
  nand n26286(x26286, x25772, x26274);
  nand n26287(x26287, x26286, x26285);
  nand n26288(x26288, x71987, x26277);
  nand n26289(x26289, x25782, x84032);
  nand n26290(x26290, x71992, x26281);
  nand n26291(x26291, x25782, x26284);
  nand n26292(x26292, x26291, x26290);
  nand n26293(x26293, x71992, x26287);
  nand n26294(x26294, x25782, x84033);
  nand n26295(x26295, x26294, x26293);
  nand n26296(x26296, x25790, x84034);
  nand n26297(x26297, x71997, x26292);
  nand n26298(x26298, x25790, x26295);
  nand n26299(x26299, x26298, x26297);
  nand n26300(x26300, x72002, x84035);
  nand n26301(x26301, x25796, x26299);
  nand n26302(x26302, x26301, x26300);
  nand n26303(x26303, x71977, x16776);
  nand n26304(x26304, x16876, x71687);
  nand n26305(x26305, x71977, x71687);
  nand n26306(x26306, x16876, x25696);
  nand n26307(x26307, x26306, x26305);
  nand n26308(x26308, x71977, x83899);
  nand n26309(x26309, x16876, x24415);
  nand n26310(x26310, x71977, x17793);
  nand n26311(x26311, x16876, x17793);
  nand n26312(x26312, x26311, x26310);
  nand n26313(x26313, x71977, x24944);
  nand n26314(x26314, x16876, x24902);
  nand n26315(x26315, x26314, x26313);
  nand n26316(x26316, x71977, x18259);
  nand n26317(x26317, x26306, x26316);
  nand n26318(x26318, x16876, x17028);
  nand n26319(x26319, x26318, x26316);
  nand n26320(x26320, x71977, x24771);
  nand n26321(x26321, x25749, x84036);
  nand n26322(x26322, x25749, x84037);
  nand n26323(x26323, x71982, x26307);
  nand n26324(x26324, x25749, x84038);
  nand n26325(x26325, x26324, x26323);
  nand n26326(x26326, x71982, x84039);
  nand n26327(x26327, x25749, x26312);
  nand n26328(x26328, x26327, x26326);
  nand n26329(x26329, x71982, x26315);
  nand n26330(x26330, x25749, x26317);
  nand n26331(x26331, x26330, x26329);
  nand n26332(x26332, x71982, x84038);
  nand n26333(x26333, x25749, x84039);
  nand n26334(x26334, x26333, x26332);
  nand n26335(x26335, x71982, x26312);
  nand n26336(x26336, x25749, x26315);
  nand n26337(x26337, x26336, x26335);
  nand n26338(x26338, x71982, x26319);
  nand n26339(x26339, x25749, x84040);
  nand n26340(x26340, x26339, x26338);
  nand n26341(x26341, x71987, x84041);
  nand n26342(x26342, x71987, x84042);
  nand n26343(x26343, x25772, x26325);
  nand n26344(x26344, x26343, x26342);
  nand n26345(x26345, x71987, x26328);
  nand n26346(x26346, x25772, x26331);
  nand n26347(x26347, x26346, x26345);
  nand n26348(x26348, x71987, x26334);
  nand n26349(x26349, x25772, x26337);
  nand n26350(x26350, x26349, x26348);
  nand n26351(x26351, x71987, x26340);
  nand n26352(x26352, x25782, x84043);
  nand n26353(x26353, x71992, x26344);
  nand n26354(x26354, x25782, x26347);
  nand n26355(x26355, x26354, x26353);
  nand n26356(x26356, x71992, x26350);
  nand n26357(x26357, x25782, x84044);
  nand n26358(x26358, x26357, x26356);
  nand n26359(x26359, x25790, x84045);
  nand n26360(x26360, x71997, x26355);
  nand n26361(x26361, x25790, x26358);
  nand n26362(x26362, x26361, x26360);
  nand n26363(x26363, x72002, x84046);
  nand n26364(x26364, x25796, x26362);
  nand n26365(x26365, x26364, x26363);
  nand n26366(x26366, x71977, x16779);
  nand n26367(x26367, x16876, x71692);
  nand n26368(x26368, x71977, x71692);
  nand n26369(x26369, x16876, x25699);
  nand n26370(x26370, x26369, x26368);
  nand n26371(x26371, x71977, x83900);
  nand n26372(x26372, x16876, x24419);
  nand n26373(x26373, x71977, x17798);
  nand n26374(x26374, x16876, x17798);
  nand n26375(x26375, x26374, x26373);
  nand n26376(x26376, x71977, x24946);
  nand n26377(x26377, x16876, x24903);
  nand n26378(x26378, x26377, x26376);
  nand n26379(x26379, x71977, x18338);
  nand n26380(x26380, x26369, x26379);
  nand n26381(x26381, x16876, x17034);
  nand n26382(x26382, x26381, x26379);
  nand n26383(x26383, x71977, x24775);
  nand n26384(x26384, x25749, x84047);
  nand n26385(x26385, x25749, x84048);
  nand n26386(x26386, x71982, x26370);
  nand n26387(x26387, x25749, x84049);
  nand n26388(x26388, x26387, x26386);
  nand n26389(x26389, x71982, x84050);
  nand n26390(x26390, x25749, x26375);
  nand n26391(x26391, x26390, x26389);
  nand n26392(x26392, x71982, x26378);
  nand n26393(x26393, x25749, x26380);
  nand n26394(x26394, x26393, x26392);
  nand n26395(x26395, x71982, x84049);
  nand n26396(x26396, x25749, x84050);
  nand n26397(x26397, x26396, x26395);
  nand n26398(x26398, x71982, x26375);
  nand n26399(x26399, x25749, x26378);
  nand n26400(x26400, x26399, x26398);
  nand n26401(x26401, x71982, x26382);
  nand n26402(x26402, x25749, x84051);
  nand n26403(x26403, x26402, x26401);
  nand n26404(x26404, x71987, x84052);
  nand n26405(x26405, x71987, x84053);
  nand n26406(x26406, x25772, x26388);
  nand n26407(x26407, x26406, x26405);
  nand n26408(x26408, x71987, x26391);
  nand n26409(x26409, x25772, x26394);
  nand n26410(x26410, x26409, x26408);
  nand n26411(x26411, x71987, x26397);
  nand n26412(x26412, x25772, x26400);
  nand n26413(x26413, x26412, x26411);
  nand n26414(x26414, x71987, x26403);
  nand n26415(x26415, x25782, x84054);
  nand n26416(x26416, x71992, x26407);
  nand n26417(x26417, x25782, x26410);
  nand n26418(x26418, x26417, x26416);
  nand n26419(x26419, x71992, x26413);
  nand n26420(x26420, x25782, x84055);
  nand n26421(x26421, x26420, x26419);
  nand n26422(x26422, x25790, x84056);
  nand n26423(x26423, x71997, x26418);
  nand n26424(x26424, x25790, x26421);
  nand n26425(x26425, x26424, x26423);
  nand n26426(x26426, x72002, x84057);
  nand n26427(x26427, x25796, x26425);
  nand n26428(x26428, x26427, x26426);
  nand n26429(x26429, x71977, x16782);
  nand n26430(x26430, x16876, x71697);
  nand n26431(x26431, x71977, x71697);
  nand n26432(x26432, x16876, x25702);
  nand n26433(x26433, x26432, x26431);
  nand n26434(x26434, x71977, x83901);
  nand n26435(x26435, x16876, x24423);
  nand n26436(x26436, x71977, x17803);
  nand n26437(x26437, x16876, x17803);
  nand n26438(x26438, x26437, x26436);
  nand n26439(x26439, x71977, x24948);
  nand n26440(x26440, x16876, x24904);
  nand n26441(x26441, x26440, x26439);
  nand n26442(x26442, x71977, x18425);
  nand n26443(x26443, x26432, x26442);
  nand n26444(x26444, x16876, x17040);
  nand n26445(x26445, x26444, x26442);
  nand n26446(x26446, x71977, x24779);
  nand n26447(x26447, x25749, x84058);
  nand n26448(x26448, x25749, x84059);
  nand n26449(x26449, x71982, x26433);
  nand n26450(x26450, x25749, x84060);
  nand n26451(x26451, x26450, x26449);
  nand n26452(x26452, x71982, x84061);
  nand n26453(x26453, x25749, x26438);
  nand n26454(x26454, x26453, x26452);
  nand n26455(x26455, x71982, x26441);
  nand n26456(x26456, x25749, x26443);
  nand n26457(x26457, x26456, x26455);
  nand n26458(x26458, x71982, x84060);
  nand n26459(x26459, x25749, x84061);
  nand n26460(x26460, x26459, x26458);
  nand n26461(x26461, x71982, x26438);
  nand n26462(x26462, x25749, x26441);
  nand n26463(x26463, x26462, x26461);
  nand n26464(x26464, x71982, x26445);
  nand n26465(x26465, x25749, x84062);
  nand n26466(x26466, x26465, x26464);
  nand n26467(x26467, x71987, x84063);
  nand n26468(x26468, x71987, x84064);
  nand n26469(x26469, x25772, x26451);
  nand n26470(x26470, x26469, x26468);
  nand n26471(x26471, x71987, x26454);
  nand n26472(x26472, x25772, x26457);
  nand n26473(x26473, x26472, x26471);
  nand n26474(x26474, x71987, x26460);
  nand n26475(x26475, x25772, x26463);
  nand n26476(x26476, x26475, x26474);
  nand n26477(x26477, x71987, x26466);
  nand n26478(x26478, x25782, x84065);
  nand n26479(x26479, x71992, x26470);
  nand n26480(x26480, x25782, x26473);
  nand n26481(x26481, x26480, x26479);
  nand n26482(x26482, x71992, x26476);
  nand n26483(x26483, x25782, x84066);
  nand n26484(x26484, x26483, x26482);
  nand n26485(x26485, x25790, x84067);
  nand n26486(x26486, x71997, x26481);
  nand n26487(x26487, x25790, x26484);
  nand n26488(x26488, x26487, x26486);
  nand n26489(x26489, x72002, x84068);
  nand n26490(x26490, x25796, x26488);
  nand n26491(x26491, x26490, x26489);
  nand n26492(x26492, x71977, x16785);
  nand n26493(x26493, x16876, x71702);
  nand n26494(x26494, x71977, x71702);
  nand n26495(x26495, x16876, x25705);
  nand n26496(x26496, x26495, x26494);
  nand n26497(x26497, x71977, x83902);
  nand n26498(x26498, x16876, x24427);
  nand n26499(x26499, x71977, x17808);
  nand n26500(x26500, x16876, x17808);
  nand n26501(x26501, x26500, x26499);
  nand n26502(x26502, x71977, x24950);
  nand n26503(x26503, x16876, x24905);
  nand n26504(x26504, x26503, x26502);
  nand n26505(x26505, x71977, x18521);
  nand n26506(x26506, x26495, x26505);
  nand n26507(x26507, x16876, x17046);
  nand n26508(x26508, x26507, x26505);
  nand n26509(x26509, x71977, x24783);
  nand n26510(x26510, x25749, x84069);
  nand n26511(x26511, x25749, x84070);
  nand n26512(x26512, x71982, x26496);
  nand n26513(x26513, x25749, x84071);
  nand n26514(x26514, x26513, x26512);
  nand n26515(x26515, x71982, x84072);
  nand n26516(x26516, x25749, x26501);
  nand n26517(x26517, x26516, x26515);
  nand n26518(x26518, x71982, x26504);
  nand n26519(x26519, x25749, x26506);
  nand n26520(x26520, x26519, x26518);
  nand n26521(x26521, x71982, x84071);
  nand n26522(x26522, x25749, x84072);
  nand n26523(x26523, x26522, x26521);
  nand n26524(x26524, x71982, x26501);
  nand n26525(x26525, x25749, x26504);
  nand n26526(x26526, x26525, x26524);
  nand n26527(x26527, x71982, x26508);
  nand n26528(x26528, x25749, x84073);
  nand n26529(x26529, x26528, x26527);
  nand n26530(x26530, x71987, x84074);
  nand n26531(x26531, x71987, x84075);
  nand n26532(x26532, x25772, x26514);
  nand n26533(x26533, x26532, x26531);
  nand n26534(x26534, x71987, x26517);
  nand n26535(x26535, x25772, x26520);
  nand n26536(x26536, x26535, x26534);
  nand n26537(x26537, x71987, x26523);
  nand n26538(x26538, x25772, x26526);
  nand n26539(x26539, x26538, x26537);
  nand n26540(x26540, x71987, x26529);
  nand n26541(x26541, x25782, x84076);
  nand n26542(x26542, x71992, x26533);
  nand n26543(x26543, x25782, x26536);
  nand n26544(x26544, x26543, x26542);
  nand n26545(x26545, x71992, x26539);
  nand n26546(x26546, x25782, x84077);
  nand n26547(x26547, x26546, x26545);
  nand n26548(x26548, x25790, x84078);
  nand n26549(x26549, x71997, x26544);
  nand n26550(x26550, x25790, x26547);
  nand n26551(x26551, x26550, x26549);
  nand n26552(x26552, x72002, x84079);
  nand n26553(x26553, x25796, x26551);
  nand n26554(x26554, x26553, x26552);
  nand n26555(x26555, x71977, x16788);
  nand n26556(x26556, x16876, x71707);
  nand n26557(x26557, x71977, x71707);
  nand n26558(x26558, x16876, x25708);
  nand n26559(x26559, x26558, x26557);
  nand n26560(x26560, x71977, x83903);
  nand n26561(x26561, x16876, x24431);
  nand n26562(x26562, x71977, x17813);
  nand n26563(x26563, x16876, x17813);
  nand n26564(x26564, x26563, x26562);
  nand n26565(x26565, x71977, x24952);
  nand n26566(x26566, x16876, x24906);
  nand n26567(x26567, x26566, x26565);
  nand n26568(x26568, x71977, x18624);
  nand n26569(x26569, x26558, x26568);
  nand n26570(x26570, x16876, x17052);
  nand n26571(x26571, x26570, x26568);
  nand n26572(x26572, x71977, x24787);
  nand n26573(x26573, x25749, x84080);
  nand n26574(x26574, x25749, x84081);
  nand n26575(x26575, x71982, x26559);
  nand n26576(x26576, x25749, x84082);
  nand n26577(x26577, x26576, x26575);
  nand n26578(x26578, x71982, x84083);
  nand n26579(x26579, x25749, x26564);
  nand n26580(x26580, x26579, x26578);
  nand n26581(x26581, x71982, x26567);
  nand n26582(x26582, x25749, x26569);
  nand n26583(x26583, x26582, x26581);
  nand n26584(x26584, x71982, x84082);
  nand n26585(x26585, x25749, x84083);
  nand n26586(x26586, x26585, x26584);
  nand n26587(x26587, x71982, x26564);
  nand n26588(x26588, x25749, x26567);
  nand n26589(x26589, x26588, x26587);
  nand n26590(x26590, x71982, x26571);
  nand n26591(x26591, x25749, x84084);
  nand n26592(x26592, x26591, x26590);
  nand n26593(x26593, x71987, x84085);
  nand n26594(x26594, x71987, x84086);
  nand n26595(x26595, x25772, x26577);
  nand n26596(x26596, x26595, x26594);
  nand n26597(x26597, x71987, x26580);
  nand n26598(x26598, x25772, x26583);
  nand n26599(x26599, x26598, x26597);
  nand n26600(x26600, x71987, x26586);
  nand n26601(x26601, x25772, x26589);
  nand n26602(x26602, x26601, x26600);
  nand n26603(x26603, x71987, x26592);
  nand n26604(x26604, x25782, x84087);
  nand n26605(x26605, x71992, x26596);
  nand n26606(x26606, x25782, x26599);
  nand n26607(x26607, x26606, x26605);
  nand n26608(x26608, x71992, x26602);
  nand n26609(x26609, x25782, x84088);
  nand n26610(x26610, x26609, x26608);
  nand n26611(x26611, x25790, x84089);
  nand n26612(x26612, x71997, x26607);
  nand n26613(x26613, x25790, x26610);
  nand n26614(x26614, x26613, x26612);
  nand n26615(x26615, x72002, x84090);
  nand n26616(x26616, x25796, x26614);
  nand n26617(x26617, x26616, x26615);
  nand n26618(x26618, x71977, x16791);
  nand n26619(x26619, x16876, x71712);
  nand n26620(x26620, x71977, x71712);
  nand n26621(x26621, x16876, x25711);
  nand n26622(x26622, x26621, x26620);
  nand n26623(x26623, x71977, x83904);
  nand n26624(x26624, x16876, x24436);
  nand n26625(x26625, x71977, x17818);
  nand n26626(x26626, x16876, x17818);
  nand n26627(x26627, x26626, x26625);
  nand n26628(x26628, x71977, x24954);
  nand n26629(x26629, x16876, x24907);
  nand n26630(x26630, x26629, x26628);
  nand n26631(x26631, x71977, x18735);
  nand n26632(x26632, x26621, x26631);
  nand n26633(x26633, x16876, x17058);
  nand n26634(x26634, x26633, x26631);
  nand n26635(x26635, x71977, x24791);
  nand n26636(x26636, x25749, x84091);
  nand n26637(x26637, x25749, x84092);
  nand n26638(x26638, x71982, x26622);
  nand n26639(x26639, x25749, x84093);
  nand n26640(x26640, x26639, x26638);
  nand n26641(x26641, x71982, x84094);
  nand n26642(x26642, x25749, x26627);
  nand n26643(x26643, x26642, x26641);
  nand n26644(x26644, x71982, x26630);
  nand n26645(x26645, x25749, x26632);
  nand n26646(x26646, x26645, x26644);
  nand n26647(x26647, x71982, x84093);
  nand n26648(x26648, x25749, x84094);
  nand n26649(x26649, x26648, x26647);
  nand n26650(x26650, x71982, x26627);
  nand n26651(x26651, x25749, x26630);
  nand n26652(x26652, x26651, x26650);
  nand n26653(x26653, x71982, x26634);
  nand n26654(x26654, x25749, x84095);
  nand n26655(x26655, x26654, x26653);
  nand n26656(x26656, x71987, x84096);
  nand n26657(x26657, x71987, x84097);
  nand n26658(x26658, x25772, x26640);
  nand n26659(x26659, x26658, x26657);
  nand n26660(x26660, x71987, x26643);
  nand n26661(x26661, x25772, x26646);
  nand n26662(x26662, x26661, x26660);
  nand n26663(x26663, x71987, x26649);
  nand n26664(x26664, x25772, x26652);
  nand n26665(x26665, x26664, x26663);
  nand n26666(x26666, x71987, x26655);
  nand n26667(x26667, x25782, x84098);
  nand n26668(x26668, x71992, x26659);
  nand n26669(x26669, x25782, x26662);
  nand n26670(x26670, x26669, x26668);
  nand n26671(x26671, x71992, x26665);
  nand n26672(x26672, x25782, x84099);
  nand n26673(x26673, x26672, x26671);
  nand n26674(x26674, x25790, x84100);
  nand n26675(x26675, x71997, x26670);
  nand n26676(x26676, x25790, x26673);
  nand n26677(x26677, x26676, x26675);
  nand n26678(x26678, x72002, x84101);
  nand n26679(x26679, x25796, x26677);
  nand n26680(x26680, x26679, x26678);
  nand n26681(x26681, x71977, x16794);
  nand n26682(x26682, x16876, x71717);
  nand n26683(x26683, x71977, x71717);
  nand n26684(x26684, x16876, x25714);
  nand n26685(x26685, x26684, x26683);
  nand n26686(x26686, x71977, x83905);
  nand n26687(x26687, x16876, x24441);
  nand n26688(x26688, x71977, x17823);
  nand n26689(x26689, x16876, x17823);
  nand n26690(x26690, x26689, x26688);
  nand n26691(x26691, x71977, x24956);
  nand n26692(x26692, x16876, x24908);
  nand n26693(x26693, x26692, x26691);
  nand n26694(x26694, x71977, x18855);
  nand n26695(x26695, x26684, x26694);
  nand n26696(x26696, x16876, x17064);
  nand n26697(x26697, x26696, x26694);
  nand n26698(x26698, x71977, x24795);
  nand n26699(x26699, x25749, x84102);
  nand n26700(x26700, x25749, x84103);
  nand n26701(x26701, x71982, x26685);
  nand n26702(x26702, x25749, x84104);
  nand n26703(x26703, x26702, x26701);
  nand n26704(x26704, x71982, x84105);
  nand n26705(x26705, x25749, x26690);
  nand n26706(x26706, x26705, x26704);
  nand n26707(x26707, x71982, x26693);
  nand n26708(x26708, x25749, x26695);
  nand n26709(x26709, x26708, x26707);
  nand n26710(x26710, x71982, x84104);
  nand n26711(x26711, x25749, x84105);
  nand n26712(x26712, x26711, x26710);
  nand n26713(x26713, x71982, x26690);
  nand n26714(x26714, x25749, x26693);
  nand n26715(x26715, x26714, x26713);
  nand n26716(x26716, x71982, x26697);
  nand n26717(x26717, x25749, x84106);
  nand n26718(x26718, x26717, x26716);
  nand n26719(x26719, x71987, x84107);
  nand n26720(x26720, x71987, x84108);
  nand n26721(x26721, x25772, x26703);
  nand n26722(x26722, x26721, x26720);
  nand n26723(x26723, x71987, x26706);
  nand n26724(x26724, x25772, x26709);
  nand n26725(x26725, x26724, x26723);
  nand n26726(x26726, x71987, x26712);
  nand n26727(x26727, x25772, x26715);
  nand n26728(x26728, x26727, x26726);
  nand n26729(x26729, x71987, x26718);
  nand n26730(x26730, x25782, x84109);
  nand n26731(x26731, x71992, x26722);
  nand n26732(x26732, x25782, x26725);
  nand n26733(x26733, x26732, x26731);
  nand n26734(x26734, x71992, x26728);
  nand n26735(x26735, x25782, x84110);
  nand n26736(x26736, x26735, x26734);
  nand n26737(x26737, x25790, x84111);
  nand n26738(x26738, x71997, x26733);
  nand n26739(x26739, x25790, x26736);
  nand n26740(x26740, x26739, x26738);
  nand n26741(x26741, x72002, x84112);
  nand n26742(x26742, x25796, x26740);
  nand n26743(x26743, x26742, x26741);
  nand n26744(x26744, x71977, x16797);
  nand n26745(x26745, x16876, x71722);
  nand n26746(x26746, x71977, x71722);
  nand n26747(x26747, x16876, x83921);
  nand n26748(x26748, x26747, x26746);
  nand n26749(x26749, x71977, x25330);
  nand n26750(x26750, x16876, x24445);
  nand n26751(x26751, x71977, x17828);
  nand n26752(x26752, x16876, x17828);
  nand n26753(x26753, x26752, x26751);
  nand n26754(x26754, x71977, x24958);
  nand n26755(x26755, x16876, x24909);
  nand n26756(x26756, x26755, x26754);
  nand n26757(x26757, x71977, x24862);
  nand n26758(x26758, x26747, x26757);
  nand n26759(x26759, x16876, x17070);
  nand n26760(x26760, x26759, x26757);
  nand n26761(x26761, x71977, x24799);
  nand n26762(x26762, x25749, x84113);
  nand n26763(x26763, x25749, x84114);
  nand n26764(x26764, x71982, x26748);
  nand n26765(x26765, x25749, x84115);
  nand n26766(x26766, x26765, x26764);
  nand n26767(x26767, x71982, x84116);
  nand n26768(x26768, x25749, x26753);
  nand n26769(x26769, x26768, x26767);
  nand n26770(x26770, x71982, x26756);
  nand n26771(x26771, x25749, x26758);
  nand n26772(x26772, x26771, x26770);
  nand n26773(x26773, x71982, x84115);
  nand n26774(x26774, x25749, x84116);
  nand n26775(x26775, x26774, x26773);
  nand n26776(x26776, x71982, x26753);
  nand n26777(x26777, x25749, x26756);
  nand n26778(x26778, x26777, x26776);
  nand n26779(x26779, x71982, x26760);
  nand n26780(x26780, x25749, x84117);
  nand n26781(x26781, x26780, x26779);
  nand n26782(x26782, x71987, x84118);
  nand n26783(x26783, x71987, x84119);
  nand n26784(x26784, x25772, x26766);
  nand n26785(x26785, x26784, x26783);
  nand n26786(x26786, x71987, x26769);
  nand n26787(x26787, x25772, x26772);
  nand n26788(x26788, x26787, x26786);
  nand n26789(x26789, x71987, x26775);
  nand n26790(x26790, x25772, x26778);
  nand n26791(x26791, x26790, x26789);
  nand n26792(x26792, x71987, x26781);
  nand n26793(x26793, x25782, x84120);
  nand n26794(x26794, x71992, x26785);
  nand n26795(x26795, x25782, x26788);
  nand n26796(x26796, x26795, x26794);
  nand n26797(x26797, x71992, x26791);
  nand n26798(x26798, x25782, x84121);
  nand n26799(x26799, x26798, x26797);
  nand n26800(x26800, x25790, x84122);
  nand n26801(x26801, x71997, x26796);
  nand n26802(x26802, x25790, x26799);
  nand n26803(x26803, x26802, x26801);
  nand n26804(x26804, x72002, x84123);
  nand n26805(x26805, x25796, x26803);
  nand n26806(x26806, x26805, x26804);
  nand n26807(x26807, x71977, x16800);
  nand n26808(x26808, x16876, x71727);
  nand n26809(x26809, x71977, x71727);
  nand n26810(x26810, x16876, x83922);
  nand n26811(x26811, x26810, x26809);
  nand n26812(x26812, x71977, x25333);
  nand n26813(x26813, x16876, x24449);
  nand n26814(x26814, x71977, x17833);
  nand n26815(x26815, x16876, x17833);
  nand n26816(x26816, x26815, x26814);
  nand n26817(x26817, x71977, x24960);
  nand n26818(x26818, x16876, x24910);
  nand n26819(x26819, x26818, x26817);
  nand n26820(x26820, x71977, x24864);
  nand n26821(x26821, x26810, x26820);
  nand n26822(x26822, x16876, x17076);
  nand n26823(x26823, x26822, x26820);
  nand n26824(x26824, x71977, x24803);
  nand n26825(x26825, x25749, x84124);
  nand n26826(x26826, x25749, x84125);
  nand n26827(x26827, x71982, x26811);
  nand n26828(x26828, x25749, x84126);
  nand n26829(x26829, x26828, x26827);
  nand n26830(x26830, x71982, x84127);
  nand n26831(x26831, x25749, x26816);
  nand n26832(x26832, x26831, x26830);
  nand n26833(x26833, x71982, x26819);
  nand n26834(x26834, x25749, x26821);
  nand n26835(x26835, x26834, x26833);
  nand n26836(x26836, x71982, x84126);
  nand n26837(x26837, x25749, x84127);
  nand n26838(x26838, x26837, x26836);
  nand n26839(x26839, x71982, x26816);
  nand n26840(x26840, x25749, x26819);
  nand n26841(x26841, x26840, x26839);
  nand n26842(x26842, x71982, x26823);
  nand n26843(x26843, x25749, x84128);
  nand n26844(x26844, x26843, x26842);
  nand n26845(x26845, x71987, x84129);
  nand n26846(x26846, x71987, x84130);
  nand n26847(x26847, x25772, x26829);
  nand n26848(x26848, x26847, x26846);
  nand n26849(x26849, x71987, x26832);
  nand n26850(x26850, x25772, x26835);
  nand n26851(x26851, x26850, x26849);
  nand n26852(x26852, x71987, x26838);
  nand n26853(x26853, x25772, x26841);
  nand n26854(x26854, x26853, x26852);
  nand n26855(x26855, x71987, x26844);
  nand n26856(x26856, x25782, x84131);
  nand n26857(x26857, x71992, x26848);
  nand n26858(x26858, x25782, x26851);
  nand n26859(x26859, x26858, x26857);
  nand n26860(x26860, x71992, x26854);
  nand n26861(x26861, x25782, x84132);
  nand n26862(x26862, x26861, x26860);
  nand n26863(x26863, x25790, x84133);
  nand n26864(x26864, x71997, x26859);
  nand n26865(x26865, x25790, x26862);
  nand n26866(x26866, x26865, x26864);
  nand n26867(x26867, x72002, x84134);
  nand n26868(x26868, x25796, x26866);
  nand n26869(x26869, x26868, x26867);
  nand n26870(x26870, x71977, x16803);
  nand n26871(x26871, x16876, x71732);
  nand n26872(x26872, x71977, x71732);
  nand n26873(x26873, x16876, x83923);
  nand n26874(x26874, x26873, x26872);
  nand n26875(x26875, x71977, x25336);
  nand n26876(x26876, x16876, x24453);
  nand n26877(x26877, x71977, x17838);
  nand n26878(x26878, x16876, x17838);
  nand n26879(x26879, x26878, x26877);
  nand n26880(x26880, x71977, x24962);
  nand n26881(x26881, x16876, x24911);
  nand n26882(x26882, x26881, x26880);
  nand n26883(x26883, x71977, x24866);
  nand n26884(x26884, x26873, x26883);
  nand n26885(x26885, x16876, x17082);
  nand n26886(x26886, x26885, x26883);
  nand n26887(x26887, x71977, x24807);
  nand n26888(x26888, x25749, x84135);
  nand n26889(x26889, x25749, x84136);
  nand n26890(x26890, x71982, x26874);
  nand n26891(x26891, x25749, x84137);
  nand n26892(x26892, x26891, x26890);
  nand n26893(x26893, x71982, x84138);
  nand n26894(x26894, x25749, x26879);
  nand n26895(x26895, x26894, x26893);
  nand n26896(x26896, x71982, x26882);
  nand n26897(x26897, x25749, x26884);
  nand n26898(x26898, x26897, x26896);
  nand n26899(x26899, x71982, x84137);
  nand n26900(x26900, x25749, x84138);
  nand n26901(x26901, x26900, x26899);
  nand n26902(x26902, x71982, x26879);
  nand n26903(x26903, x25749, x26882);
  nand n26904(x26904, x26903, x26902);
  nand n26905(x26905, x71982, x26886);
  nand n26906(x26906, x25749, x84139);
  nand n26907(x26907, x26906, x26905);
  nand n26908(x26908, x71987, x84140);
  nand n26909(x26909, x71987, x84141);
  nand n26910(x26910, x25772, x26892);
  nand n26911(x26911, x26910, x26909);
  nand n26912(x26912, x71987, x26895);
  nand n26913(x26913, x25772, x26898);
  nand n26914(x26914, x26913, x26912);
  nand n26915(x26915, x71987, x26901);
  nand n26916(x26916, x25772, x26904);
  nand n26917(x26917, x26916, x26915);
  nand n26918(x26918, x71987, x26907);
  nand n26919(x26919, x25782, x84142);
  nand n26920(x26920, x71992, x26911);
  nand n26921(x26921, x25782, x26914);
  nand n26922(x26922, x26921, x26920);
  nand n26923(x26923, x71992, x26917);
  nand n26924(x26924, x25782, x84143);
  nand n26925(x26925, x26924, x26923);
  nand n26926(x26926, x25790, x84144);
  nand n26927(x26927, x71997, x26922);
  nand n26928(x26928, x25790, x26925);
  nand n26929(x26929, x26928, x26927);
  nand n26930(x26930, x72002, x84145);
  nand n26931(x26931, x25796, x26929);
  nand n26932(x26932, x26931, x26930);
  nand n26933(x26933, x71977, x16806);
  nand n26934(x26934, x16876, x71737);
  nand n26935(x26935, x71977, x71737);
  nand n26936(x26936, x16876, x83924);
  nand n26937(x26937, x26936, x26935);
  nand n26938(x26938, x71977, x25339);
  nand n26939(x26939, x16876, x24457);
  nand n26940(x26940, x71977, x17843);
  nand n26941(x26941, x16876, x17843);
  nand n26942(x26942, x26941, x26940);
  nand n26943(x26943, x71977, x24964);
  nand n26944(x26944, x16876, x24912);
  nand n26945(x26945, x26944, x26943);
  nand n26946(x26946, x71977, x24868);
  nand n26947(x26947, x26936, x26946);
  nand n26948(x26948, x16876, x17088);
  nand n26949(x26949, x26948, x26946);
  nand n26950(x26950, x71977, x24811);
  nand n26951(x26951, x25749, x84146);
  nand n26952(x26952, x25749, x84147);
  nand n26953(x26953, x71982, x26937);
  nand n26954(x26954, x25749, x84148);
  nand n26955(x26955, x26954, x26953);
  nand n26956(x26956, x71982, x84149);
  nand n26957(x26957, x25749, x26942);
  nand n26958(x26958, x26957, x26956);
  nand n26959(x26959, x71982, x26945);
  nand n26960(x26960, x25749, x26947);
  nand n26961(x26961, x26960, x26959);
  nand n26962(x26962, x71982, x84148);
  nand n26963(x26963, x25749, x84149);
  nand n26964(x26964, x26963, x26962);
  nand n26965(x26965, x71982, x26942);
  nand n26966(x26966, x25749, x26945);
  nand n26967(x26967, x26966, x26965);
  nand n26968(x26968, x71982, x26949);
  nand n26969(x26969, x25749, x84150);
  nand n26970(x26970, x26969, x26968);
  nand n26971(x26971, x71987, x84151);
  nand n26972(x26972, x71987, x84152);
  nand n26973(x26973, x25772, x26955);
  nand n26974(x26974, x26973, x26972);
  nand n26975(x26975, x71987, x26958);
  nand n26976(x26976, x25772, x26961);
  nand n26977(x26977, x26976, x26975);
  nand n26978(x26978, x71987, x26964);
  nand n26979(x26979, x25772, x26967);
  nand n26980(x26980, x26979, x26978);
  nand n26981(x26981, x71987, x26970);
  nand n26982(x26982, x25782, x84153);
  nand n26983(x26983, x71992, x26974);
  nand n26984(x26984, x25782, x26977);
  nand n26985(x26985, x26984, x26983);
  nand n26986(x26986, x71992, x26980);
  nand n26987(x26987, x25782, x84154);
  nand n26988(x26988, x26987, x26986);
  nand n26989(x26989, x25790, x84155);
  nand n26990(x26990, x71997, x26985);
  nand n26991(x26991, x25790, x26988);
  nand n26992(x26992, x26991, x26990);
  nand n26993(x26993, x72002, x84156);
  nand n26994(x26994, x25796, x26992);
  nand n26995(x26995, x26994, x26993);
  nand n26996(x26996, x71977, x16809);
  nand n26997(x26997, x16876, x71742);
  nand n26998(x26998, x71977, x71742);
  nand n26999(x26999, x16876, x83925);
  nand n27000(x27000, x26999, x26998);
  nand n27001(x27001, x71977, x25342);
  nand n27002(x27002, x16876, x24461);
  nand n27003(x27003, x71977, x17848);
  nand n27004(x27004, x16876, x17848);
  nand n27005(x27005, x27004, x27003);
  nand n27006(x27006, x71977, x24966);
  nand n27007(x27007, x16876, x24913);
  nand n27008(x27008, x27007, x27006);
  nand n27009(x27009, x71977, x24870);
  nand n27010(x27010, x26999, x27009);
  nand n27011(x27011, x16876, x17094);
  nand n27012(x27012, x27011, x27009);
  nand n27013(x27013, x71977, x24815);
  nand n27014(x27014, x25749, x84157);
  nand n27015(x27015, x25749, x84158);
  nand n27016(x27016, x71982, x27000);
  nand n27017(x27017, x25749, x84159);
  nand n27018(x27018, x27017, x27016);
  nand n27019(x27019, x71982, x84160);
  nand n27020(x27020, x25749, x27005);
  nand n27021(x27021, x27020, x27019);
  nand n27022(x27022, x71982, x27008);
  nand n27023(x27023, x25749, x27010);
  nand n27024(x27024, x27023, x27022);
  nand n27025(x27025, x71982, x84159);
  nand n27026(x27026, x25749, x84160);
  nand n27027(x27027, x27026, x27025);
  nand n27028(x27028, x71982, x27005);
  nand n27029(x27029, x25749, x27008);
  nand n27030(x27030, x27029, x27028);
  nand n27031(x27031, x71982, x27012);
  nand n27032(x27032, x25749, x84161);
  nand n27033(x27033, x27032, x27031);
  nand n27034(x27034, x71987, x84162);
  nand n27035(x27035, x71987, x84163);
  nand n27036(x27036, x25772, x27018);
  nand n27037(x27037, x27036, x27035);
  nand n27038(x27038, x71987, x27021);
  nand n27039(x27039, x25772, x27024);
  nand n27040(x27040, x27039, x27038);
  nand n27041(x27041, x71987, x27027);
  nand n27042(x27042, x25772, x27030);
  nand n27043(x27043, x27042, x27041);
  nand n27044(x27044, x71987, x27033);
  nand n27045(x27045, x25782, x84164);
  nand n27046(x27046, x71992, x27037);
  nand n27047(x27047, x25782, x27040);
  nand n27048(x27048, x27047, x27046);
  nand n27049(x27049, x71992, x27043);
  nand n27050(x27050, x25782, x84165);
  nand n27051(x27051, x27050, x27049);
  nand n27052(x27052, x25790, x84166);
  nand n27053(x27053, x71997, x27048);
  nand n27054(x27054, x25790, x27051);
  nand n27055(x27055, x27054, x27053);
  nand n27056(x27056, x72002, x84167);
  nand n27057(x27057, x25796, x27055);
  nand n27058(x27058, x27057, x27056);
  nand n27059(x27059, x71977, x16812);
  nand n27060(x27060, x16876, x71747);
  nand n27061(x27061, x71977, x71747);
  nand n27062(x27062, x16876, x83926);
  nand n27063(x27063, x27062, x27061);
  nand n27064(x27064, x71977, x25345);
  nand n27065(x27065, x16876, x24465);
  nand n27066(x27066, x71977, x17853);
  nand n27067(x27067, x16876, x17853);
  nand n27068(x27068, x27067, x27066);
  nand n27069(x27069, x71977, x24968);
  nand n27070(x27070, x16876, x24914);
  nand n27071(x27071, x27070, x27069);
  nand n27072(x27072, x71977, x24872);
  nand n27073(x27073, x27062, x27072);
  nand n27074(x27074, x16876, x17100);
  nand n27075(x27075, x27074, x27072);
  nand n27076(x27076, x71977, x24819);
  nand n27077(x27077, x25749, x84168);
  nand n27078(x27078, x25749, x84169);
  nand n27079(x27079, x71982, x27063);
  nand n27080(x27080, x25749, x84170);
  nand n27081(x27081, x27080, x27079);
  nand n27082(x27082, x71982, x84171);
  nand n27083(x27083, x25749, x27068);
  nand n27084(x27084, x27083, x27082);
  nand n27085(x27085, x71982, x27071);
  nand n27086(x27086, x25749, x27073);
  nand n27087(x27087, x27086, x27085);
  nand n27088(x27088, x71982, x84170);
  nand n27089(x27089, x25749, x84171);
  nand n27090(x27090, x27089, x27088);
  nand n27091(x27091, x71982, x27068);
  nand n27092(x27092, x25749, x27071);
  nand n27093(x27093, x27092, x27091);
  nand n27094(x27094, x71982, x27075);
  nand n27095(x27095, x25749, x84172);
  nand n27096(x27096, x27095, x27094);
  nand n27097(x27097, x71987, x84173);
  nand n27098(x27098, x71987, x84174);
  nand n27099(x27099, x25772, x27081);
  nand n27100(x27100, x27099, x27098);
  nand n27101(x27101, x71987, x27084);
  nand n27102(x27102, x25772, x27087);
  nand n27103(x27103, x27102, x27101);
  nand n27104(x27104, x71987, x27090);
  nand n27105(x27105, x25772, x27093);
  nand n27106(x27106, x27105, x27104);
  nand n27107(x27107, x71987, x27096);
  nand n27108(x27108, x25782, x84175);
  nand n27109(x27109, x71992, x27100);
  nand n27110(x27110, x25782, x27103);
  nand n27111(x27111, x27110, x27109);
  nand n27112(x27112, x71992, x27106);
  nand n27113(x27113, x25782, x84176);
  nand n27114(x27114, x27113, x27112);
  nand n27115(x27115, x25790, x84177);
  nand n27116(x27116, x71997, x27111);
  nand n27117(x27117, x25790, x27114);
  nand n27118(x27118, x27117, x27116);
  nand n27119(x27119, x72002, x84178);
  nand n27120(x27120, x25796, x27118);
  nand n27121(x27121, x27120, x27119);
  nand n27122(x27122, x71977, x16815);
  nand n27123(x27123, x16876, x71752);
  nand n27124(x27124, x71977, x71752);
  nand n27125(x27125, x16876, x83927);
  nand n27126(x27126, x27125, x27124);
  nand n27127(x27127, x71977, x25348);
  nand n27128(x27128, x16876, x24470);
  nand n27129(x27129, x71977, x17858);
  nand n27130(x27130, x16876, x17858);
  nand n27131(x27131, x27130, x27129);
  nand n27132(x27132, x71977, x24970);
  nand n27133(x27133, x16876, x24915);
  nand n27134(x27134, x27133, x27132);
  nand n27135(x27135, x71977, x24874);
  nand n27136(x27136, x27125, x27135);
  nand n27137(x27137, x16876, x17106);
  nand n27138(x27138, x27137, x27135);
  nand n27139(x27139, x71977, x24823);
  nand n27140(x27140, x25749, x84179);
  nand n27141(x27141, x25749, x84180);
  nand n27142(x27142, x71982, x27126);
  nand n27143(x27143, x25749, x84181);
  nand n27144(x27144, x27143, x27142);
  nand n27145(x27145, x71982, x84182);
  nand n27146(x27146, x25749, x27131);
  nand n27147(x27147, x27146, x27145);
  nand n27148(x27148, x71982, x27134);
  nand n27149(x27149, x25749, x27136);
  nand n27150(x27150, x27149, x27148);
  nand n27151(x27151, x71982, x84181);
  nand n27152(x27152, x25749, x84182);
  nand n27153(x27153, x27152, x27151);
  nand n27154(x27154, x71982, x27131);
  nand n27155(x27155, x25749, x27134);
  nand n27156(x27156, x27155, x27154);
  nand n27157(x27157, x71982, x27138);
  nand n27158(x27158, x25749, x84183);
  nand n27159(x27159, x27158, x27157);
  nand n27160(x27160, x71987, x84184);
  nand n27161(x27161, x71987, x84185);
  nand n27162(x27162, x25772, x27144);
  nand n27163(x27163, x27162, x27161);
  nand n27164(x27164, x71987, x27147);
  nand n27165(x27165, x25772, x27150);
  nand n27166(x27166, x27165, x27164);
  nand n27167(x27167, x71987, x27153);
  nand n27168(x27168, x25772, x27156);
  nand n27169(x27169, x27168, x27167);
  nand n27170(x27170, x71987, x27159);
  nand n27171(x27171, x25782, x84186);
  nand n27172(x27172, x71992, x27163);
  nand n27173(x27173, x25782, x27166);
  nand n27174(x27174, x27173, x27172);
  nand n27175(x27175, x71992, x27169);
  nand n27176(x27176, x25782, x84187);
  nand n27177(x27177, x27176, x27175);
  nand n27178(x27178, x25790, x84188);
  nand n27179(x27179, x71997, x27174);
  nand n27180(x27180, x25790, x27177);
  nand n27181(x27181, x27180, x27179);
  nand n27182(x27182, x72002, x84189);
  nand n27183(x27183, x25796, x27181);
  nand n27184(x27184, x27183, x27182);
  nand n27185(x27185, x71977, x16818);
  nand n27186(x27186, x16876, x71757);
  nand n27187(x27187, x71977, x71757);
  nand n27188(x27188, x16876, x83928);
  nand n27189(x27189, x27188, x27187);
  nand n27190(x27190, x71977, x25351);
  nand n27191(x27191, x16876, x24475);
  nand n27192(x27192, x71977, x17863);
  nand n27193(x27193, x16876, x17863);
  nand n27194(x27194, x27193, x27192);
  nand n27195(x27195, x71977, x24972);
  nand n27196(x27196, x16876, x24916);
  nand n27197(x27197, x27196, x27195);
  nand n27198(x27198, x71977, x24876);
  nand n27199(x27199, x27188, x27198);
  nand n27200(x27200, x16876, x17112);
  nand n27201(x27201, x27200, x27198);
  nand n27202(x27202, x71977, x24827);
  nand n27203(x27203, x25749, x84190);
  nand n27204(x27204, x25749, x84191);
  nand n27205(x27205, x71982, x27189);
  nand n27206(x27206, x25749, x84192);
  nand n27207(x27207, x27206, x27205);
  nand n27208(x27208, x71982, x84193);
  nand n27209(x27209, x25749, x27194);
  nand n27210(x27210, x27209, x27208);
  nand n27211(x27211, x71982, x27197);
  nand n27212(x27212, x25749, x27199);
  nand n27213(x27213, x27212, x27211);
  nand n27214(x27214, x71982, x84192);
  nand n27215(x27215, x25749, x84193);
  nand n27216(x27216, x27215, x27214);
  nand n27217(x27217, x71982, x27194);
  nand n27218(x27218, x25749, x27197);
  nand n27219(x27219, x27218, x27217);
  nand n27220(x27220, x71982, x27201);
  nand n27221(x27221, x25749, x84194);
  nand n27222(x27222, x27221, x27220);
  nand n27223(x27223, x71987, x84195);
  nand n27224(x27224, x71987, x84196);
  nand n27225(x27225, x25772, x27207);
  nand n27226(x27226, x27225, x27224);
  nand n27227(x27227, x71987, x27210);
  nand n27228(x27228, x25772, x27213);
  nand n27229(x27229, x27228, x27227);
  nand n27230(x27230, x71987, x27216);
  nand n27231(x27231, x25772, x27219);
  nand n27232(x27232, x27231, x27230);
  nand n27233(x27233, x71987, x27222);
  nand n27234(x27234, x25782, x84197);
  nand n27235(x27235, x71992, x27226);
  nand n27236(x27236, x25782, x27229);
  nand n27237(x27237, x27236, x27235);
  nand n27238(x27238, x71992, x27232);
  nand n27239(x27239, x25782, x84198);
  nand n27240(x27240, x27239, x27238);
  nand n27241(x27241, x25790, x84199);
  nand n27242(x27242, x71997, x27237);
  nand n27243(x27243, x25790, x27240);
  nand n27244(x27244, x27243, x27242);
  nand n27245(x27245, x72002, x84200);
  nand n27246(x27246, x25796, x27244);
  nand n27247(x27247, x27246, x27245);
  nand n27248(x27248, x71977, x16821);
  nand n27249(x27249, x16876, x71762);
  nand n27250(x27250, x71977, x71762);
  nand n27251(x27251, x16876, x83929);
  nand n27252(x27252, x27251, x27250);
  nand n27253(x27253, x71977, x25354);
  nand n27254(x27254, x16876, x24480);
  nand n27255(x27255, x71977, x17868);
  nand n27256(x27256, x16876, x17868);
  nand n27257(x27257, x27256, x27255);
  nand n27258(x27258, x71977, x24974);
  nand n27259(x27259, x16876, x24917);
  nand n27260(x27260, x27259, x27258);
  nand n27261(x27261, x71977, x24878);
  nand n27262(x27262, x27251, x27261);
  nand n27263(x27263, x16876, x17118);
  nand n27264(x27264, x27263, x27261);
  nand n27265(x27265, x71977, x24831);
  nand n27266(x27266, x25749, x84201);
  nand n27267(x27267, x25749, x84202);
  nand n27268(x27268, x71982, x27252);
  nand n27269(x27269, x25749, x84203);
  nand n27270(x27270, x27269, x27268);
  nand n27271(x27271, x71982, x84204);
  nand n27272(x27272, x25749, x27257);
  nand n27273(x27273, x27272, x27271);
  nand n27274(x27274, x71982, x27260);
  nand n27275(x27275, x25749, x27262);
  nand n27276(x27276, x27275, x27274);
  nand n27277(x27277, x71982, x84203);
  nand n27278(x27278, x25749, x84204);
  nand n27279(x27279, x27278, x27277);
  nand n27280(x27280, x71982, x27257);
  nand n27281(x27281, x25749, x27260);
  nand n27282(x27282, x27281, x27280);
  nand n27283(x27283, x71982, x27264);
  nand n27284(x27284, x25749, x84205);
  nand n27285(x27285, x27284, x27283);
  nand n27286(x27286, x71987, x84206);
  nand n27287(x27287, x71987, x84207);
  nand n27288(x27288, x25772, x27270);
  nand n27289(x27289, x27288, x27287);
  nand n27290(x27290, x71987, x27273);
  nand n27291(x27291, x25772, x27276);
  nand n27292(x27292, x27291, x27290);
  nand n27293(x27293, x71987, x27279);
  nand n27294(x27294, x25772, x27282);
  nand n27295(x27295, x27294, x27293);
  nand n27296(x27296, x71987, x27285);
  nand n27297(x27297, x25782, x84208);
  nand n27298(x27298, x71992, x27289);
  nand n27299(x27299, x25782, x27292);
  nand n27300(x27300, x27299, x27298);
  nand n27301(x27301, x71992, x27295);
  nand n27302(x27302, x25782, x84209);
  nand n27303(x27303, x27302, x27301);
  nand n27304(x27304, x25790, x84210);
  nand n27305(x27305, x71997, x27300);
  nand n27306(x27306, x25790, x27303);
  nand n27307(x27307, x27306, x27305);
  nand n27308(x27308, x72002, x84211);
  nand n27309(x27309, x25796, x27307);
  nand n27310(x27310, x27309, x27308);
  nand n27311(x27311, x71977, x16824);
  nand n27312(x27312, x16876, x71767);
  nand n27313(x27313, x71977, x71767);
  nand n27314(x27314, x16876, x83930);
  nand n27315(x27315, x27314, x27313);
  nand n27316(x27316, x71977, x25357);
  nand n27317(x27317, x16876, x24485);
  nand n27318(x27318, x71977, x17873);
  nand n27319(x27319, x16876, x17873);
  nand n27320(x27320, x27319, x27318);
  nand n27321(x27321, x71977, x24976);
  nand n27322(x27322, x16876, x24918);
  nand n27323(x27323, x27322, x27321);
  nand n27324(x27324, x71977, x24880);
  nand n27325(x27325, x27314, x27324);
  nand n27326(x27326, x16876, x17124);
  nand n27327(x27327, x27326, x27324);
  nand n27328(x27328, x71977, x24835);
  nand n27329(x27329, x25749, x84212);
  nand n27330(x27330, x25749, x84213);
  nand n27331(x27331, x71982, x27315);
  nand n27332(x27332, x25749, x84214);
  nand n27333(x27333, x27332, x27331);
  nand n27334(x27334, x71982, x84215);
  nand n27335(x27335, x25749, x27320);
  nand n27336(x27336, x27335, x27334);
  nand n27337(x27337, x71982, x27323);
  nand n27338(x27338, x25749, x27325);
  nand n27339(x27339, x27338, x27337);
  nand n27340(x27340, x71982, x84214);
  nand n27341(x27341, x25749, x84215);
  nand n27342(x27342, x27341, x27340);
  nand n27343(x27343, x71982, x27320);
  nand n27344(x27344, x25749, x27323);
  nand n27345(x27345, x27344, x27343);
  nand n27346(x27346, x71982, x27327);
  nand n27347(x27347, x25749, x84216);
  nand n27348(x27348, x27347, x27346);
  nand n27349(x27349, x71987, x84217);
  nand n27350(x27350, x71987, x84218);
  nand n27351(x27351, x25772, x27333);
  nand n27352(x27352, x27351, x27350);
  nand n27353(x27353, x71987, x27336);
  nand n27354(x27354, x25772, x27339);
  nand n27355(x27355, x27354, x27353);
  nand n27356(x27356, x71987, x27342);
  nand n27357(x27357, x25772, x27345);
  nand n27358(x27358, x27357, x27356);
  nand n27359(x27359, x71987, x27348);
  nand n27360(x27360, x25782, x84219);
  nand n27361(x27361, x71992, x27352);
  nand n27362(x27362, x25782, x27355);
  nand n27363(x27363, x27362, x27361);
  nand n27364(x27364, x71992, x27358);
  nand n27365(x27365, x25782, x84220);
  nand n27366(x27366, x27365, x27364);
  nand n27367(x27367, x25790, x84221);
  nand n27368(x27368, x71997, x27363);
  nand n27369(x27369, x25790, x27366);
  nand n27370(x27370, x27369, x27368);
  nand n27371(x27371, x72002, x84222);
  nand n27372(x27372, x25796, x27370);
  nand n27373(x27373, x27372, x27371);
  nand n27374(x27374, x71977, x16827);
  nand n27375(x27375, x16876, x71772);
  nand n27376(x27376, x71977, x71772);
  nand n27377(x27377, x16876, x83931);
  nand n27378(x27378, x27377, x27376);
  nand n27379(x27379, x71977, x25360);
  nand n27380(x27380, x16876, x24490);
  nand n27381(x27381, x71977, x17878);
  nand n27382(x27382, x16876, x17878);
  nand n27383(x27383, x27382, x27381);
  nand n27384(x27384, x71977, x24978);
  nand n27385(x27385, x16876, x24919);
  nand n27386(x27386, x27385, x27384);
  nand n27387(x27387, x71977, x24882);
  nand n27388(x27388, x27377, x27387);
  nand n27389(x27389, x16876, x17130);
  nand n27390(x27390, x27389, x27387);
  nand n27391(x27391, x71977, x24839);
  nand n27392(x27392, x25749, x84223);
  nand n27393(x27393, x25749, x84224);
  nand n27394(x27394, x71982, x27378);
  nand n27395(x27395, x25749, x84225);
  nand n27396(x27396, x27395, x27394);
  nand n27397(x27397, x71982, x84226);
  nand n27398(x27398, x25749, x27383);
  nand n27399(x27399, x27398, x27397);
  nand n27400(x27400, x71982, x27386);
  nand n27401(x27401, x25749, x27388);
  nand n27402(x27402, x27401, x27400);
  nand n27403(x27403, x71982, x84225);
  nand n27404(x27404, x25749, x84226);
  nand n27405(x27405, x27404, x27403);
  nand n27406(x27406, x71982, x27383);
  nand n27407(x27407, x25749, x27386);
  nand n27408(x27408, x27407, x27406);
  nand n27409(x27409, x71982, x27390);
  nand n27410(x27410, x25749, x84227);
  nand n27411(x27411, x27410, x27409);
  nand n27412(x27412, x71987, x84228);
  nand n27413(x27413, x71987, x84229);
  nand n27414(x27414, x25772, x27396);
  nand n27415(x27415, x27414, x27413);
  nand n27416(x27416, x71987, x27399);
  nand n27417(x27417, x25772, x27402);
  nand n27418(x27418, x27417, x27416);
  nand n27419(x27419, x71987, x27405);
  nand n27420(x27420, x25772, x27408);
  nand n27421(x27421, x27420, x27419);
  nand n27422(x27422, x71987, x27411);
  nand n27423(x27423, x25782, x84230);
  nand n27424(x27424, x71992, x27415);
  nand n27425(x27425, x25782, x27418);
  nand n27426(x27426, x27425, x27424);
  nand n27427(x27427, x71992, x27421);
  nand n27428(x27428, x25782, x84231);
  nand n27429(x27429, x27428, x27427);
  nand n27430(x27430, x25790, x84232);
  nand n27431(x27431, x71997, x27426);
  nand n27432(x27432, x25790, x27429);
  nand n27433(x27433, x27432, x27431);
  nand n27434(x27434, x72002, x84233);
  nand n27435(x27435, x25796, x27433);
  nand n27436(x27436, x27435, x27434);
  nand n27437(x27437, x71977, x16830);
  nand n27438(x27438, x16876, x71777);
  nand n27439(x27439, x71977, x71777);
  nand n27440(x27440, x16876, x83932);
  nand n27441(x27441, x27440, x27439);
  nand n27442(x27442, x71977, x25363);
  nand n27443(x27443, x16876, x24495);
  nand n27444(x27444, x71977, x17883);
  nand n27445(x27445, x16876, x17883);
  nand n27446(x27446, x27445, x27444);
  nand n27447(x27447, x71977, x24980);
  nand n27448(x27448, x16876, x24920);
  nand n27449(x27449, x27448, x27447);
  nand n27450(x27450, x71977, x24884);
  nand n27451(x27451, x27440, x27450);
  nand n27452(x27452, x16876, x17136);
  nand n27453(x27453, x27452, x27450);
  nand n27454(x27454, x71977, x24843);
  nand n27455(x27455, x25749, x84234);
  nand n27456(x27456, x25749, x84235);
  nand n27457(x27457, x71982, x27441);
  nand n27458(x27458, x25749, x84236);
  nand n27459(x27459, x27458, x27457);
  nand n27460(x27460, x71982, x84237);
  nand n27461(x27461, x25749, x27446);
  nand n27462(x27462, x27461, x27460);
  nand n27463(x27463, x71982, x27449);
  nand n27464(x27464, x25749, x27451);
  nand n27465(x27465, x27464, x27463);
  nand n27466(x27466, x71982, x84236);
  nand n27467(x27467, x25749, x84237);
  nand n27468(x27468, x27467, x27466);
  nand n27469(x27469, x71982, x27446);
  nand n27470(x27470, x25749, x27449);
  nand n27471(x27471, x27470, x27469);
  nand n27472(x27472, x71982, x27453);
  nand n27473(x27473, x25749, x84238);
  nand n27474(x27474, x27473, x27472);
  nand n27475(x27475, x71987, x84239);
  nand n27476(x27476, x71987, x84240);
  nand n27477(x27477, x25772, x27459);
  nand n27478(x27478, x27477, x27476);
  nand n27479(x27479, x71987, x27462);
  nand n27480(x27480, x25772, x27465);
  nand n27481(x27481, x27480, x27479);
  nand n27482(x27482, x71987, x27468);
  nand n27483(x27483, x25772, x27471);
  nand n27484(x27484, x27483, x27482);
  nand n27485(x27485, x71987, x27474);
  nand n27486(x27486, x25782, x84241);
  nand n27487(x27487, x71992, x27478);
  nand n27488(x27488, x25782, x27481);
  nand n27489(x27489, x27488, x27487);
  nand n27490(x27490, x71992, x27484);
  nand n27491(x27491, x25782, x84242);
  nand n27492(x27492, x27491, x27490);
  nand n27493(x27493, x25790, x84243);
  nand n27494(x27494, x71997, x27489);
  nand n27495(x27495, x25790, x27492);
  nand n27496(x27496, x27495, x27494);
  nand n27497(x27497, x72002, x84244);
  nand n27498(x27498, x25796, x27496);
  nand n27499(x27499, x27498, x27497);
  nand n27500(x27500, x71977, x16833);
  nand n27501(x27501, x16876, x71782);
  nand n27502(x27502, x71977, x71782);
  nand n27503(x27503, x16876, x83933);
  nand n27504(x27504, x27503, x27502);
  nand n27505(x27505, x71977, x25366);
  nand n27506(x27506, x16876, x24500);
  nand n27507(x27507, x71977, x17888);
  nand n27508(x27508, x16876, x17888);
  nand n27509(x27509, x27508, x27507);
  nand n27510(x27510, x71977, x24982);
  nand n27511(x27511, x16876, x24921);
  nand n27512(x27512, x27511, x27510);
  nand n27513(x27513, x71977, x24886);
  nand n27514(x27514, x27503, x27513);
  nand n27515(x27515, x16876, x17142);
  nand n27516(x27516, x27515, x27513);
  nand n27517(x27517, x71977, x24847);
  nand n27518(x27518, x25749, x84245);
  nand n27519(x27519, x25749, x84246);
  nand n27520(x27520, x71982, x27504);
  nand n27521(x27521, x25749, x84247);
  nand n27522(x27522, x27521, x27520);
  nand n27523(x27523, x71982, x84248);
  nand n27524(x27524, x25749, x27509);
  nand n27525(x27525, x27524, x27523);
  nand n27526(x27526, x71982, x27512);
  nand n27527(x27527, x25749, x27514);
  nand n27528(x27528, x27527, x27526);
  nand n27529(x27529, x71982, x84247);
  nand n27530(x27530, x25749, x84248);
  nand n27531(x27531, x27530, x27529);
  nand n27532(x27532, x71982, x27509);
  nand n27533(x27533, x25749, x27512);
  nand n27534(x27534, x27533, x27532);
  nand n27535(x27535, x71982, x27516);
  nand n27536(x27536, x25749, x84249);
  nand n27537(x27537, x27536, x27535);
  nand n27538(x27538, x71987, x84250);
  nand n27539(x27539, x71987, x84251);
  nand n27540(x27540, x25772, x27522);
  nand n27541(x27541, x27540, x27539);
  nand n27542(x27542, x71987, x27525);
  nand n27543(x27543, x25772, x27528);
  nand n27544(x27544, x27543, x27542);
  nand n27545(x27545, x71987, x27531);
  nand n27546(x27546, x25772, x27534);
  nand n27547(x27547, x27546, x27545);
  nand n27548(x27548, x71987, x27537);
  nand n27549(x27549, x25782, x84252);
  nand n27550(x27550, x71992, x27541);
  nand n27551(x27551, x25782, x27544);
  nand n27552(x27552, x27551, x27550);
  nand n27553(x27553, x71992, x27547);
  nand n27554(x27554, x25782, x84253);
  nand n27555(x27555, x27554, x27553);
  nand n27556(x27556, x25790, x84254);
  nand n27557(x27557, x71997, x27552);
  nand n27558(x27558, x25790, x27555);
  nand n27559(x27559, x27558, x27557);
  nand n27560(x27560, x72002, x84255);
  nand n27561(x27561, x25796, x27559);
  nand n27562(x27562, x27561, x27560);
  nand n27563(x27563, x71977, x16836);
  nand n27564(x27564, x16876, x71787);
  nand n27565(x27565, x71977, x71787);
  nand n27566(x27566, x16876, x83934);
  nand n27567(x27567, x27566, x27565);
  nand n27568(x27568, x71977, x25369);
  nand n27569(x27569, x16876, x24505);
  nand n27570(x27570, x71977, x17893);
  nand n27571(x27571, x16876, x17893);
  nand n27572(x27572, x27571, x27570);
  nand n27573(x27573, x71977, x24984);
  nand n27574(x27574, x16876, x24922);
  nand n27575(x27575, x27574, x27573);
  nand n27576(x27576, x71977, x24888);
  nand n27577(x27577, x27566, x27576);
  nand n27578(x27578, x16876, x17148);
  nand n27579(x27579, x27578, x27576);
  nand n27580(x27580, x71977, x24851);
  nand n27581(x27581, x25749, x84256);
  nand n27582(x27582, x25749, x84257);
  nand n27583(x27583, x71982, x27567);
  nand n27584(x27584, x25749, x84258);
  nand n27585(x27585, x27584, x27583);
  nand n27586(x27586, x71982, x84259);
  nand n27587(x27587, x25749, x27572);
  nand n27588(x27588, x27587, x27586);
  nand n27589(x27589, x71982, x27575);
  nand n27590(x27590, x25749, x27577);
  nand n27591(x27591, x27590, x27589);
  nand n27592(x27592, x71982, x84258);
  nand n27593(x27593, x25749, x84259);
  nand n27594(x27594, x27593, x27592);
  nand n27595(x27595, x71982, x27572);
  nand n27596(x27596, x25749, x27575);
  nand n27597(x27597, x27596, x27595);
  nand n27598(x27598, x71982, x27579);
  nand n27599(x27599, x25749, x84260);
  nand n27600(x27600, x27599, x27598);
  nand n27601(x27601, x71987, x84261);
  nand n27602(x27602, x71987, x84262);
  nand n27603(x27603, x25772, x27585);
  nand n27604(x27604, x27603, x27602);
  nand n27605(x27605, x71987, x27588);
  nand n27606(x27606, x25772, x27591);
  nand n27607(x27607, x27606, x27605);
  nand n27608(x27608, x71987, x27594);
  nand n27609(x27609, x25772, x27597);
  nand n27610(x27610, x27609, x27608);
  nand n27611(x27611, x71987, x27600);
  nand n27612(x27612, x25782, x84263);
  nand n27613(x27613, x71992, x27604);
  nand n27614(x27614, x25782, x27607);
  nand n27615(x27615, x27614, x27613);
  nand n27616(x27616, x71992, x27610);
  nand n27617(x27617, x25782, x84264);
  nand n27618(x27618, x27617, x27616);
  nand n27619(x27619, x25790, x84265);
  nand n27620(x27620, x71997, x27615);
  nand n27621(x27621, x25790, x27618);
  nand n27622(x27622, x27621, x27620);
  nand n27623(x27623, x72002, x84266);
  nand n27624(x27624, x25796, x27622);
  nand n27625(x27625, x27624, x27623);
  nand n27626(x27626, x71977, x16839);
  nand n27627(x27627, x16876, x71792);
  nand n27628(x27628, x71977, x71792);
  nand n27629(x27629, x16876, x83935);
  nand n27630(x27630, x27629, x27628);
  nand n27631(x27631, x71977, x25372);
  nand n27632(x27632, x16876, x24510);
  nand n27633(x27633, x71977, x17898);
  nand n27634(x27634, x16876, x17898);
  nand n27635(x27635, x27634, x27633);
  nand n27636(x27636, x71977, x24986);
  nand n27637(x27637, x16876, x24923);
  nand n27638(x27638, x27637, x27636);
  nand n27639(x27639, x71977, x24890);
  nand n27640(x27640, x27629, x27639);
  nand n27641(x27641, x16876, x17154);
  nand n27642(x27642, x27641, x27639);
  nand n27643(x27643, x71977, x24855);
  nand n27644(x27644, x25749, x84267);
  nand n27645(x27645, x25749, x84268);
  nand n27646(x27646, x71982, x27630);
  nand n27647(x27647, x25749, x84269);
  nand n27648(x27648, x27647, x27646);
  nand n27649(x27649, x71982, x84270);
  nand n27650(x27650, x25749, x27635);
  nand n27651(x27651, x27650, x27649);
  nand n27652(x27652, x71982, x27638);
  nand n27653(x27653, x25749, x27640);
  nand n27654(x27654, x27653, x27652);
  nand n27655(x27655, x71982, x84269);
  nand n27656(x27656, x25749, x84270);
  nand n27657(x27657, x27656, x27655);
  nand n27658(x27658, x71982, x27635);
  nand n27659(x27659, x25749, x27638);
  nand n27660(x27660, x27659, x27658);
  nand n27661(x27661, x71982, x27642);
  nand n27662(x27662, x25749, x84271);
  nand n27663(x27663, x27662, x27661);
  nand n27664(x27664, x71987, x84272);
  nand n27665(x27665, x71987, x84273);
  nand n27666(x27666, x25772, x27648);
  nand n27667(x27667, x27666, x27665);
  nand n27668(x27668, x71987, x27651);
  nand n27669(x27669, x25772, x27654);
  nand n27670(x27670, x27669, x27668);
  nand n27671(x27671, x71987, x27657);
  nand n27672(x27672, x25772, x27660);
  nand n27673(x27673, x27672, x27671);
  nand n27674(x27674, x71987, x27663);
  nand n27675(x27675, x25782, x84274);
  nand n27676(x27676, x71992, x27667);
  nand n27677(x27677, x25782, x27670);
  nand n27678(x27678, x27677, x27676);
  nand n27679(x27679, x71992, x27673);
  nand n27680(x27680, x25782, x84275);
  nand n27681(x27681, x27680, x27679);
  nand n27682(x27682, x25790, x84276);
  nand n27683(x27683, x71997, x27678);
  nand n27684(x27684, x25790, x27681);
  nand n27685(x27685, x27684, x27683);
  nand n27686(x27686, x72002, x84277);
  nand n27687(x27687, x25796, x27685);
  nand n27688(x27688, x27687, x27686);
  nand n27689(x27689, x71977, x16842);
  nand n27690(x27690, x16876, x71797);
  nand n27691(x27691, x71977, x71797);
  nand n27692(x27692, x16876, x83936);
  nand n27693(x27693, x27692, x27691);
  nand n27694(x27694, x71977, x25375);
  nand n27695(x27695, x16876, x24515);
  nand n27696(x27696, x71977, x17903);
  nand n27697(x27697, x16876, x17903);
  nand n27698(x27698, x27697, x27696);
  nand n27699(x27699, x71977, x24988);
  nand n27700(x27700, x16876, x24924);
  nand n27701(x27701, x27700, x27699);
  nand n27702(x27702, x71977, x24892);
  nand n27703(x27703, x27692, x27702);
  nand n27704(x27704, x16876, x17160);
  nand n27705(x27705, x27704, x27702);
  nand n27706(x27706, x71977, x24859);
  nand n27707(x27707, x25749, x84278);
  nand n27708(x27708, x25749, x84279);
  nand n27709(x27709, x71982, x27693);
  nand n27710(x27710, x25749, x84280);
  nand n27711(x27711, x27710, x27709);
  nand n27712(x27712, x71982, x84281);
  nand n27713(x27713, x25749, x27698);
  nand n27714(x27714, x27713, x27712);
  nand n27715(x27715, x71982, x27701);
  nand n27716(x27716, x25749, x27703);
  nand n27717(x27717, x27716, x27715);
  nand n27718(x27718, x71982, x84280);
  nand n27719(x27719, x25749, x84281);
  nand n27720(x27720, x27719, x27718);
  nand n27721(x27721, x71982, x27698);
  nand n27722(x27722, x25749, x27701);
  nand n27723(x27723, x27722, x27721);
  nand n27724(x27724, x71982, x27705);
  nand n27725(x27725, x25749, x84282);
  nand n27726(x27726, x27725, x27724);
  nand n27727(x27727, x71987, x84283);
  nand n27728(x27728, x71987, x84284);
  nand n27729(x27729, x25772, x27711);
  nand n27730(x27730, x27729, x27728);
  nand n27731(x27731, x71987, x27714);
  nand n27732(x27732, x25772, x27717);
  nand n27733(x27733, x27732, x27731);
  nand n27734(x27734, x71987, x27720);
  nand n27735(x27735, x25772, x27723);
  nand n27736(x27736, x27735, x27734);
  nand n27737(x27737, x71987, x27726);
  nand n27738(x27738, x25782, x84285);
  nand n27739(x27739, x71992, x27730);
  nand n27740(x27740, x25782, x27733);
  nand n27741(x27741, x27740, x27739);
  nand n27742(x27742, x71992, x27736);
  nand n27743(x27743, x25782, x84286);
  nand n27744(x27744, x27743, x27742);
  nand n27745(x27745, x25790, x84287);
  nand n27746(x27746, x71997, x27741);
  nand n27747(x27747, x25790, x27744);
  nand n27748(x27748, x27747, x27746);
  nand n27749(x27749, x72002, x84288);
  nand n27750(x27750, x25796, x27748);
  nand n27751(x27751, x27750, x27749);
  nand n27752(x27752, x16745, x25798);
  nand n27753(x27753, x68738, x27755);
  nand n27754(x27754, x27753, x27752);
  nand n27756(x27756, x16745, x25861);
  nand n27757(x27757, x68738, x27759);
  nand n27758(x27758, x27757, x27756);
  nand n27760(x27760, x16745, x25924);
  nand n27761(x27761, x68738, x27763);
  nand n27762(x27762, x27761, x27760);
  nand n27764(x27764, x16745, x25987);
  nand n27765(x27765, x68738, x27767);
  nand n27766(x27766, x27765, x27764);
  nand n27768(x27768, x16745, x26050);
  nand n27769(x27769, x68738, x27771);
  nand n27770(x27770, x27769, x27768);
  nand n27772(x27772, x16745, x26113);
  nand n27773(x27773, x68738, x27775);
  nand n27774(x27774, x27773, x27772);
  nand n27776(x27776, x16745, x26176);
  nand n27777(x27777, x68738, x27779);
  nand n27778(x27778, x27777, x27776);
  nand n27780(x27780, x16745, x26239);
  nand n27781(x27781, x68738, x27783);
  nand n27782(x27782, x27781, x27780);
  nand n27784(x27784, x16745, x26302);
  nand n27785(x27785, x68738, x27787);
  nand n27786(x27786, x27785, x27784);
  nand n27788(x27788, x16745, x26365);
  nand n27789(x27789, x68738, x27791);
  nand n27790(x27790, x27789, x27788);
  nand n27792(x27792, x16745, x26428);
  nand n27793(x27793, x68738, x27795);
  nand n27794(x27794, x27793, x27792);
  nand n27796(x27796, x16745, x26491);
  nand n27797(x27797, x68738, x27799);
  nand n27798(x27798, x27797, x27796);
  nand n27800(x27800, x16745, x26554);
  nand n27801(x27801, x68738, x27803);
  nand n27802(x27802, x27801, x27800);
  nand n27804(x27804, x16745, x26617);
  nand n27805(x27805, x68738, x27807);
  nand n27806(x27806, x27805, x27804);
  nand n27808(x27808, x16745, x26680);
  nand n27809(x27809, x68738, x27811);
  nand n27810(x27810, x27809, x27808);
  nand n27812(x27812, x16745, x26743);
  nand n27813(x27813, x68738, x27815);
  nand n27814(x27814, x27813, x27812);
  nand n27816(x27816, x16745, x26806);
  nand n27817(x27817, x68738, x27819);
  nand n27818(x27818, x27817, x27816);
  nand n27820(x27820, x16745, x26869);
  nand n27821(x27821, x68738, x27823);
  nand n27822(x27822, x27821, x27820);
  nand n27824(x27824, x16745, x26932);
  nand n27825(x27825, x68738, x27827);
  nand n27826(x27826, x27825, x27824);
  nand n27828(x27828, x16745, x26995);
  nand n27829(x27829, x68738, x27831);
  nand n27830(x27830, x27829, x27828);
  nand n27832(x27832, x16745, x27058);
  nand n27833(x27833, x68738, x27835);
  nand n27834(x27834, x27833, x27832);
  nand n27836(x27836, x16745, x27121);
  nand n27837(x27837, x68738, x27839);
  nand n27838(x27838, x27837, x27836);
  nand n27840(x27840, x16745, x27184);
  nand n27841(x27841, x68738, x27843);
  nand n27842(x27842, x27841, x27840);
  nand n27844(x27844, x16745, x27247);
  nand n27845(x27845, x68738, x27847);
  nand n27846(x27846, x27845, x27844);
  nand n27848(x27848, x16745, x27310);
  nand n27849(x27849, x68738, x27851);
  nand n27850(x27850, x27849, x27848);
  nand n27852(x27852, x16745, x27373);
  nand n27853(x27853, x68738, x27855);
  nand n27854(x27854, x27853, x27852);
  nand n27856(x27856, x16745, x27436);
  nand n27857(x27857, x68738, x27859);
  nand n27858(x27858, x27857, x27856);
  nand n27860(x27860, x16745, x27499);
  nand n27861(x27861, x68738, x27863);
  nand n27862(x27862, x27861, x27860);
  nand n27864(x27864, x16745, x27562);
  nand n27865(x27865, x68738, x27867);
  nand n27866(x27866, x27865, x27864);
  nand n27868(x27868, x16745, x27625);
  nand n27869(x27869, x68738, x27871);
  nand n27870(x27870, x27869, x27868);
  nand n27872(x27872, x16745, x27688);
  nand n27873(x27873, x68738, x27875);
  nand n27874(x27874, x27873, x27872);
  nand n27876(x27876, x16745, x27751);
  nand n27877(x27877, x68738, x27879);
  nand n27878(x27878, x27877, x27876);
  nand n27880(x27880, x16747, x72697);
  nand n27881(x27881, x27880, x16746);
  nand n27882(x27882, x16747, x72702);
  nand n27883(x27883, x27882, x16750);
  nand n27884(x27884, x16747, x72707);
  nand n27885(x27885, x27884, x16753);
  nand n27886(x27886, x16747, x72712);
  nand n27887(x27887, x27886, x16756);
  nand n27888(x27888, x16747, x72717);
  nand n27889(x27889, x27888, x16759);
  nand n27890(x27890, x16747, x72722);
  nand n27891(x27891, x27890, x16762);
  nand n27892(x27892, x16747, x72727);
  nand n27893(x27893, x27892, x16765);
  nand n27894(x27894, x16747, x72732);
  nand n27895(x27895, x27894, x16768);
  nand n27896(x27896, x16747, x72737);
  nand n27897(x27897, x27896, x16771);
  nand n27898(x27898, x16747, x72742);
  nand n27899(x27899, x27898, x16774);
  nand n27900(x27900, x16747, x72747);
  nand n27901(x27901, x27900, x16777);
  nand n27902(x27902, x16747, x72752);
  nand n27903(x27903, x27902, x16780);
  nand n27904(x27904, x16747, x72757);
  nand n27905(x27905, x27904, x16783);
  nand n27906(x27906, x16747, x72762);
  nand n27907(x27907, x27906, x16786);
  nand n27908(x27908, x16747, x72767);
  nand n27909(x27909, x27908, x16789);
  nand n27910(x27910, x16747, x72772);
  nand n27911(x27911, x27910, x16792);
  nand n27912(x27912, x16747, x72777);
  nand n27913(x27913, x27912, x16795);
  nand n27914(x27914, x16747, x72782);
  nand n27915(x27915, x27914, x16798);
  nand n27916(x27916, x16747, x72787);
  nand n27917(x27917, x27916, x16801);
  nand n27918(x27918, x16747, x72792);
  nand n27919(x27919, x27918, x16804);
  nand n27920(x27920, x16747, x72797);
  nand n27921(x27921, x27920, x16807);
  nand n27922(x27922, x16747, x72802);
  nand n27923(x27923, x27922, x16810);
  nand n27924(x27924, x16747, x72807);
  nand n27925(x27925, x27924, x16813);
  nand n27926(x27926, x16747, x72812);
  nand n27927(x27927, x27926, x16816);
  nand n27928(x27928, x16747, x72817);
  nand n27929(x27929, x27928, x16819);
  nand n27930(x27930, x16747, x72822);
  nand n27931(x27931, x27930, x16822);
  nand n27932(x27932, x16747, x72827);
  nand n27933(x27933, x27932, x16825);
  nand n27934(x27934, x16747, x72832);
  nand n27935(x27935, x27934, x16828);
  nand n27936(x27936, x16747, x72837);
  nand n27937(x27937, x27936, x16831);
  nand n27938(x27938, x16747, x72842);
  nand n27939(x27939, x27938, x16834);
  nand n27940(x27940, x16747, x72847);
  nand n27941(x27941, x27940, x16837);
  nand n27942(x27942, x16747, x72852);
  nand n27943(x27943, x27942, x16840);
  nand n27976(x27976, x71977, x27944);
  nand n27977(x27977, x16876, x27881);
  nand n27978(x27978, x27977, x27976);
  nand n27979(x27979, x71977, x27945);
  nand n27980(x27980, x16876, x27883);
  nand n27981(x27981, x27980, x27979);
  nand n27982(x27982, x71977, x27946);
  nand n27983(x27983, x16876, x27885);
  nand n27984(x27984, x27983, x27982);
  nand n27985(x27985, x71977, x27947);
  nand n27986(x27986, x16876, x27887);
  nand n27987(x27987, x27986, x27985);
  nand n27988(x27988, x71977, x27948);
  nand n27989(x27989, x16876, x27889);
  nand n27990(x27990, x27989, x27988);
  nand n27991(x27991, x71977, x27949);
  nand n27992(x27992, x16876, x27891);
  nand n27993(x27993, x27992, x27991);
  nand n27994(x27994, x71977, x27950);
  nand n27995(x27995, x16876, x27893);
  nand n27996(x27996, x27995, x27994);
  nand n27997(x27997, x71977, x27951);
  nand n27998(x27998, x16876, x27895);
  nand n27999(x27999, x27998, x27997);
  nand n28000(x28000, x71977, x27952);
  nand n28001(x28001, x16876, x27897);
  nand n28002(x28002, x28001, x28000);
  nand n28003(x28003, x71977, x27953);
  nand n28004(x28004, x16876, x27899);
  nand n28005(x28005, x28004, x28003);
  nand n28006(x28006, x71977, x27954);
  nand n28007(x28007, x16876, x27901);
  nand n28008(x28008, x28007, x28006);
  nand n28009(x28009, x71977, x27955);
  nand n28010(x28010, x16876, x27903);
  nand n28011(x28011, x28010, x28009);
  nand n28012(x28012, x71977, x27956);
  nand n28013(x28013, x16876, x27905);
  nand n28014(x28014, x28013, x28012);
  nand n28015(x28015, x71977, x27957);
  nand n28016(x28016, x16876, x27907);
  nand n28017(x28017, x28016, x28015);
  nand n28018(x28018, x71977, x27958);
  nand n28019(x28019, x16876, x27909);
  nand n28020(x28020, x28019, x28018);
  nand n28021(x28021, x71977, x27959);
  nand n28022(x28022, x16876, x27911);
  nand n28023(x28023, x28022, x28021);
  nand n28024(x28024, x71977, x27960);
  nand n28025(x28025, x16876, x27913);
  nand n28026(x28026, x28025, x28024);
  nand n28027(x28027, x71977, x27961);
  nand n28028(x28028, x16876, x27915);
  nand n28029(x28029, x28028, x28027);
  nand n28030(x28030, x71977, x27962);
  nand n28031(x28031, x16876, x27917);
  nand n28032(x28032, x28031, x28030);
  nand n28033(x28033, x71977, x27963);
  nand n28034(x28034, x16876, x27919);
  nand n28035(x28035, x28034, x28033);
  nand n28036(x28036, x71977, x27964);
  nand n28037(x28037, x16876, x27921);
  nand n28038(x28038, x28037, x28036);
  nand n28039(x28039, x71977, x27965);
  nand n28040(x28040, x16876, x27923);
  nand n28041(x28041, x28040, x28039);
  nand n28042(x28042, x71977, x27966);
  nand n28043(x28043, x16876, x27925);
  nand n28044(x28044, x28043, x28042);
  nand n28045(x28045, x71977, x27967);
  nand n28046(x28046, x16876, x27927);
  nand n28047(x28047, x28046, x28045);
  nand n28048(x28048, x71977, x27968);
  nand n28049(x28049, x16876, x27929);
  nand n28050(x28050, x28049, x28048);
  nand n28051(x28051, x71977, x27969);
  nand n28052(x28052, x16876, x27931);
  nand n28053(x28053, x28052, x28051);
  nand n28054(x28054, x71977, x27970);
  nand n28055(x28055, x16876, x27933);
  nand n28056(x28056, x28055, x28054);
  nand n28057(x28057, x71977, x27971);
  nand n28058(x28058, x16876, x27935);
  nand n28059(x28059, x28058, x28057);
  nand n28060(x28060, x71977, x27972);
  nand n28061(x28061, x16876, x27937);
  nand n28062(x28062, x28061, x28060);
  nand n28063(x28063, x71977, x27973);
  nand n28064(x28064, x16876, x27939);
  nand n28065(x28065, x28064, x28063);
  nand n28066(x28066, x71977, x27974);
  nand n28067(x28067, x16876, x27941);
  nand n28068(x28068, x28067, x28066);
  nand n28069(x28069, x71977, x27975);
  nand n28070(x28070, x16876, x27943);
  nand n28071(x28071, x28070, x28069);
  nand n28072(x28072, x72537, x27978);
  nand n28075(x28075, x28074, x28073);
  nand n28076(x28076, x28075, x28072);
  nand n28078(x28078, x72542, x27981);
  nand n28081(x28081, x28080, x28079);
  nand n28082(x28082, x28081, x28078);
  nand n28084(x28084, x72547, x27984);
  nand n28087(x28087, x28086, x28085);
  nand n28088(x28088, x28087, x28084);
  nand n28090(x28090, x72552, x27987);
  nand n28093(x28093, x28092, x28091);
  nand n28094(x28094, x28093, x28090);
  nand n28096(x28096, x72557, x27990);
  nand n28099(x28099, x28098, x28097);
  nand n28100(x28100, x28099, x28096);
  nand n28102(x28102, x72562, x27993);
  nand n28105(x28105, x28104, x28103);
  nand n28106(x28106, x28105, x28102);
  nand n28108(x28108, x72567, x27996);
  nand n28111(x28111, x28110, x28109);
  nand n28112(x28112, x28111, x28108);
  nand n28114(x28114, x72572, x27999);
  nand n28117(x28117, x28116, x28115);
  nand n28118(x28118, x28117, x28114);
  nand n28120(x28120, x72577, x28002);
  nand n28123(x28123, x28122, x28121);
  nand n28124(x28124, x28123, x28120);
  nand n28126(x28126, x72582, x28005);
  nand n28129(x28129, x28128, x28127);
  nand n28130(x28130, x28129, x28126);
  nand n28132(x28132, x72587, x28008);
  nand n28135(x28135, x28134, x28133);
  nand n28136(x28136, x28135, x28132);
  nand n28138(x28138, x72592, x28011);
  nand n28141(x28141, x28140, x28139);
  nand n28142(x28142, x28141, x28138);
  nand n28144(x28144, x72597, x28014);
  nand n28147(x28147, x28146, x28145);
  nand n28148(x28148, x28147, x28144);
  nand n28150(x28150, x72602, x28017);
  nand n28153(x28153, x28152, x28151);
  nand n28154(x28154, x28153, x28150);
  nand n28156(x28156, x72607, x28020);
  nand n28159(x28159, x28158, x28157);
  nand n28160(x28160, x28159, x28156);
  nand n28162(x28162, x72612, x28023);
  nand n28165(x28165, x28164, x28163);
  nand n28166(x28166, x28165, x28162);
  nand n28168(x28168, x72617, x28026);
  nand n28171(x28171, x28170, x28169);
  nand n28172(x28172, x28171, x28168);
  nand n28174(x28174, x72622, x28029);
  nand n28177(x28177, x28176, x28175);
  nand n28178(x28178, x28177, x28174);
  nand n28180(x28180, x72627, x28032);
  nand n28183(x28183, x28182, x28181);
  nand n28184(x28184, x28183, x28180);
  nand n28186(x28186, x72632, x28035);
  nand n28189(x28189, x28188, x28187);
  nand n28190(x28190, x28189, x28186);
  nand n28192(x28192, x72637, x28038);
  nand n28195(x28195, x28194, x28193);
  nand n28196(x28196, x28195, x28192);
  nand n28198(x28198, x72642, x28041);
  nand n28201(x28201, x28200, x28199);
  nand n28202(x28202, x28201, x28198);
  nand n28204(x28204, x72647, x28044);
  nand n28207(x28207, x28206, x28205);
  nand n28208(x28208, x28207, x28204);
  nand n28210(x28210, x72652, x28047);
  nand n28213(x28213, x28212, x28211);
  nand n28214(x28214, x28213, x28210);
  nand n28216(x28216, x72657, x28050);
  nand n28219(x28219, x28218, x28217);
  nand n28220(x28220, x28219, x28216);
  nand n28222(x28222, x72662, x28053);
  nand n28225(x28225, x28224, x28223);
  nand n28226(x28226, x28225, x28222);
  nand n28228(x28228, x72667, x28056);
  nand n28231(x28231, x28230, x28229);
  nand n28232(x28232, x28231, x28228);
  nand n28234(x28234, x72672, x28059);
  nand n28237(x28237, x28236, x28235);
  nand n28238(x28238, x28237, x28234);
  nand n28240(x28240, x72677, x28062);
  nand n28243(x28243, x28242, x28241);
  nand n28244(x28244, x28243, x28240);
  nand n28246(x28246, x72682, x28065);
  nand n28249(x28249, x28248, x28247);
  nand n28250(x28250, x28249, x28246);
  nand n28252(x28252, x72687, x28068);
  nand n28255(x28255, x28254, x28253);
  nand n28256(x28256, x28255, x28252);
  nand n28258(x28258, x72692, x28071);
  nand n28261(x28261, x28260, x28259);
  nand n28262(x28262, x28261, x28258);
  nand n28294(x28294, x28077, x71977);
  nand n28295(x28295, x28294, x28072);
  nand n28296(x28296, x28083, x28264);
  nand n28297(x28297, x28296, x28078);
  nand n28298(x28298, x28083, x28077);
  nand n28300(x28300, x28089, x28265);
  nand n28301(x28301, x28300, x28084);
  nand n28302(x28302, x28089, x28083);
  nand n28304(x28304, x28095, x28266);
  nand n28305(x28305, x28304, x28090);
  nand n28306(x28306, x28095, x28089);
  nand n28308(x28308, x28101, x28267);
  nand n28309(x28309, x28308, x28096);
  nand n28310(x28310, x28101, x28095);
  nand n28312(x28312, x28107, x28268);
  nand n28313(x28313, x28312, x28102);
  nand n28314(x28314, x28107, x28101);
  nand n28316(x28316, x28113, x28269);
  nand n28317(x28317, x28316, x28108);
  nand n28318(x28318, x28113, x28107);
  nand n28320(x28320, x28119, x28270);
  nand n28321(x28321, x28320, x28114);
  nand n28322(x28322, x28119, x28113);
  nand n28324(x28324, x28125, x28271);
  nand n28325(x28325, x28324, x28120);
  nand n28326(x28326, x28125, x28119);
  nand n28328(x28328, x28131, x28272);
  nand n28329(x28329, x28328, x28126);
  nand n28330(x28330, x28131, x28125);
  nand n28332(x28332, x28137, x28273);
  nand n28333(x28333, x28332, x28132);
  nand n28334(x28334, x28137, x28131);
  nand n28336(x28336, x28143, x28274);
  nand n28337(x28337, x28336, x28138);
  nand n28338(x28338, x28143, x28137);
  nand n28340(x28340, x28149, x28275);
  nand n28341(x28341, x28340, x28144);
  nand n28342(x28342, x28149, x28143);
  nand n28344(x28344, x28155, x28276);
  nand n28345(x28345, x28344, x28150);
  nand n28346(x28346, x28155, x28149);
  nand n28348(x28348, x28161, x28277);
  nand n28349(x28349, x28348, x28156);
  nand n28350(x28350, x28161, x28155);
  nand n28352(x28352, x28167, x28278);
  nand n28353(x28353, x28352, x28162);
  nand n28354(x28354, x28167, x28161);
  nand n28356(x28356, x28173, x28279);
  nand n28357(x28357, x28356, x28168);
  nand n28358(x28358, x28173, x28167);
  nand n28360(x28360, x28179, x28280);
  nand n28361(x28361, x28360, x28174);
  nand n28362(x28362, x28179, x28173);
  nand n28364(x28364, x28185, x28281);
  nand n28365(x28365, x28364, x28180);
  nand n28366(x28366, x28185, x28179);
  nand n28368(x28368, x28191, x28282);
  nand n28369(x28369, x28368, x28186);
  nand n28370(x28370, x28191, x28185);
  nand n28372(x28372, x28197, x28283);
  nand n28373(x28373, x28372, x28192);
  nand n28374(x28374, x28197, x28191);
  nand n28376(x28376, x28203, x28284);
  nand n28377(x28377, x28376, x28198);
  nand n28378(x28378, x28203, x28197);
  nand n28380(x28380, x28209, x28285);
  nand n28381(x28381, x28380, x28204);
  nand n28382(x28382, x28209, x28203);
  nand n28384(x28384, x28215, x28286);
  nand n28385(x28385, x28384, x28210);
  nand n28386(x28386, x28215, x28209);
  nand n28388(x28388, x28221, x28287);
  nand n28389(x28389, x28388, x28216);
  nand n28390(x28390, x28221, x28215);
  nand n28392(x28392, x28227, x28288);
  nand n28393(x28393, x28392, x28222);
  nand n28394(x28394, x28227, x28221);
  nand n28396(x28396, x28233, x28289);
  nand n28397(x28397, x28396, x28228);
  nand n28398(x28398, x28233, x28227);
  nand n28400(x28400, x28239, x28290);
  nand n28401(x28401, x28400, x28234);
  nand n28402(x28402, x28239, x28233);
  nand n28404(x28404, x28245, x28291);
  nand n28405(x28405, x28404, x28240);
  nand n28406(x28406, x28245, x28239);
  nand n28408(x28408, x28251, x28292);
  nand n28409(x28409, x28408, x28246);
  nand n28410(x28410, x28251, x28245);
  nand n28412(x28412, x28257, x28293);
  nand n28413(x28413, x28412, x28252);
  nand n28414(x28414, x28257, x28251);
  nand n28416(x28416, x28299, x71977);
  nand n28418(x28418, x28416, x28417);
  nand n28419(x28419, x28303, x28295);
  nand n28421(x28421, x28419, x28420);
  nand n28422(x28422, x28307, x28297);
  nand n28424(x28424, x28422, x28423);
  nand n28425(x28425, x28307, x28299);
  nand n28427(x28427, x28311, x28301);
  nand n28429(x28429, x28427, x28428);
  nand n28430(x28430, x28311, x28303);
  nand n28432(x28432, x28315, x28305);
  nand n28434(x28434, x28432, x28433);
  nand n28435(x28435, x28315, x28307);
  nand n28437(x28437, x28319, x28309);
  nand n28439(x28439, x28437, x28438);
  nand n28440(x28440, x28319, x28311);
  nand n28442(x28442, x28323, x28313);
  nand n28444(x28444, x28442, x28443);
  nand n28445(x28445, x28323, x28315);
  nand n28447(x28447, x28327, x28317);
  nand n28449(x28449, x28447, x28448);
  nand n28450(x28450, x28327, x28319);
  nand n28452(x28452, x28331, x28321);
  nand n28454(x28454, x28452, x28453);
  nand n28455(x28455, x28331, x28323);
  nand n28457(x28457, x28335, x28325);
  nand n28459(x28459, x28457, x28458);
  nand n28460(x28460, x28335, x28327);
  nand n28462(x28462, x28339, x28329);
  nand n28464(x28464, x28462, x28463);
  nand n28465(x28465, x28339, x28331);
  nand n28467(x28467, x28343, x28333);
  nand n28469(x28469, x28467, x28468);
  nand n28470(x28470, x28343, x28335);
  nand n28472(x28472, x28347, x28337);
  nand n28474(x28474, x28472, x28473);
  nand n28475(x28475, x28347, x28339);
  nand n28477(x28477, x28351, x28341);
  nand n28479(x28479, x28477, x28478);
  nand n28480(x28480, x28351, x28343);
  nand n28482(x28482, x28355, x28345);
  nand n28484(x28484, x28482, x28483);
  nand n28485(x28485, x28355, x28347);
  nand n28487(x28487, x28359, x28349);
  nand n28489(x28489, x28487, x28488);
  nand n28490(x28490, x28359, x28351);
  nand n28492(x28492, x28363, x28353);
  nand n28494(x28494, x28492, x28493);
  nand n28495(x28495, x28363, x28355);
  nand n28497(x28497, x28367, x28357);
  nand n28499(x28499, x28497, x28498);
  nand n28500(x28500, x28367, x28359);
  nand n28502(x28502, x28371, x28361);
  nand n28504(x28504, x28502, x28503);
  nand n28505(x28505, x28371, x28363);
  nand n28507(x28507, x28375, x28365);
  nand n28509(x28509, x28507, x28508);
  nand n28510(x28510, x28375, x28367);
  nand n28512(x28512, x28379, x28369);
  nand n28514(x28514, x28512, x28513);
  nand n28515(x28515, x28379, x28371);
  nand n28517(x28517, x28383, x28373);
  nand n28519(x28519, x28517, x28518);
  nand n28520(x28520, x28383, x28375);
  nand n28522(x28522, x28387, x28377);
  nand n28524(x28524, x28522, x28523);
  nand n28525(x28525, x28387, x28379);
  nand n28527(x28527, x28391, x28381);
  nand n28529(x28529, x28527, x28528);
  nand n28530(x28530, x28391, x28383);
  nand n28532(x28532, x28395, x28385);
  nand n28534(x28534, x28532, x28533);
  nand n28535(x28535, x28395, x28387);
  nand n28537(x28537, x28399, x28389);
  nand n28539(x28539, x28537, x28538);
  nand n28540(x28540, x28399, x28391);
  nand n28542(x28542, x28403, x28393);
  nand n28544(x28544, x28542, x28543);
  nand n28545(x28545, x28403, x28395);
  nand n28547(x28547, x28407, x28397);
  nand n28549(x28549, x28547, x28548);
  nand n28550(x28550, x28407, x28399);
  nand n28552(x28552, x28411, x28401);
  nand n28554(x28554, x28552, x28553);
  nand n28555(x28555, x28411, x28403);
  nand n28557(x28557, x28415, x28405);
  nand n28559(x28559, x28557, x28558);
  nand n28560(x28560, x28415, x28407);
  nand n28562(x28562, x28426, x71977);
  nand n28564(x28564, x28562, x28563);
  nand n28565(x28565, x28431, x28295);
  nand n28567(x28567, x28565, x28566);
  nand n28568(x28568, x28436, x28418);
  nand n28570(x28570, x28568, x28569);
  nand n28571(x28571, x28441, x28421);
  nand n28573(x28573, x28571, x28572);
  nand n28574(x28574, x28446, x28424);
  nand n28576(x28576, x28574, x28575);
  nand n28577(x28577, x28446, x28426);
  nand n28579(x28579, x28451, x28429);
  nand n28581(x28581, x28579, x28580);
  nand n28582(x28582, x28451, x28431);
  nand n28584(x28584, x28456, x28434);
  nand n28586(x28586, x28584, x28585);
  nand n28587(x28587, x28456, x28436);
  nand n28589(x28589, x28461, x28439);
  nand n28591(x28591, x28589, x28590);
  nand n28592(x28592, x28461, x28441);
  nand n28594(x28594, x28466, x28444);
  nand n28596(x28596, x28594, x28595);
  nand n28597(x28597, x28466, x28446);
  nand n28599(x28599, x28471, x28449);
  nand n28601(x28601, x28599, x28600);
  nand n28602(x28602, x28471, x28451);
  nand n28604(x28604, x28476, x28454);
  nand n28606(x28606, x28604, x28605);
  nand n28607(x28607, x28476, x28456);
  nand n28609(x28609, x28481, x28459);
  nand n28611(x28611, x28609, x28610);
  nand n28612(x28612, x28481, x28461);
  nand n28614(x28614, x28486, x28464);
  nand n28616(x28616, x28614, x28615);
  nand n28617(x28617, x28486, x28466);
  nand n28619(x28619, x28491, x28469);
  nand n28621(x28621, x28619, x28620);
  nand n28622(x28622, x28491, x28471);
  nand n28624(x28624, x28496, x28474);
  nand n28626(x28626, x28624, x28625);
  nand n28627(x28627, x28496, x28476);
  nand n28629(x28629, x28501, x28479);
  nand n28631(x28631, x28629, x28630);
  nand n28632(x28632, x28501, x28481);
  nand n28634(x28634, x28506, x28484);
  nand n28636(x28636, x28634, x28635);
  nand n28637(x28637, x28506, x28486);
  nand n28639(x28639, x28511, x28489);
  nand n28641(x28641, x28639, x28640);
  nand n28642(x28642, x28511, x28491);
  nand n28644(x28644, x28516, x28494);
  nand n28646(x28646, x28644, x28645);
  nand n28647(x28647, x28516, x28496);
  nand n28649(x28649, x28521, x28499);
  nand n28651(x28651, x28649, x28650);
  nand n28652(x28652, x28521, x28501);
  nand n28654(x28654, x28526, x28504);
  nand n28656(x28656, x28654, x28655);
  nand n28657(x28657, x28526, x28506);
  nand n28659(x28659, x28531, x28509);
  nand n28661(x28661, x28659, x28660);
  nand n28662(x28662, x28531, x28511);
  nand n28664(x28664, x28536, x28514);
  nand n28666(x28666, x28664, x28665);
  nand n28667(x28667, x28536, x28516);
  nand n28669(x28669, x28541, x28519);
  nand n28671(x28671, x28669, x28670);
  nand n28672(x28672, x28541, x28521);
  nand n28674(x28674, x28546, x28524);
  nand n28676(x28676, x28674, x28675);
  nand n28677(x28677, x28546, x28526);
  nand n28679(x28679, x28551, x28529);
  nand n28681(x28681, x28679, x28680);
  nand n28682(x28682, x28551, x28531);
  nand n28684(x28684, x28556, x28534);
  nand n28686(x28686, x28684, x28685);
  nand n28687(x28687, x28556, x28536);
  nand n28689(x28689, x28561, x28539);
  nand n28691(x28691, x28689, x28690);
  nand n28692(x28692, x28561, x28541);
  nand n28694(x28694, x28578, x71977);
  nand n28696(x28696, x28694, x28695);
  nand n28697(x28697, x28583, x28295);
  nand n28699(x28699, x28697, x28698);
  nand n28700(x28700, x28588, x28418);
  nand n28702(x28702, x28700, x28701);
  nand n28703(x28703, x28593, x28421);
  nand n28705(x28705, x28703, x28704);
  nand n28706(x28706, x28598, x28564);
  nand n28708(x28708, x28706, x28707);
  nand n28709(x28709, x28603, x28567);
  nand n28711(x28711, x28709, x28710);
  nand n28712(x28712, x28608, x28570);
  nand n28714(x28714, x28712, x28713);
  nand n28715(x28715, x28613, x28573);
  nand n28717(x28717, x28715, x28716);
  nand n28718(x28718, x28618, x28576);
  nand n28720(x28720, x28718, x28719);
  nand n28721(x28721, x28618, x28578);
  nand n28723(x28723, x28623, x28581);
  nand n28725(x28725, x28723, x28724);
  nand n28726(x28726, x28623, x28583);
  nand n28728(x28728, x28628, x28586);
  nand n28730(x28730, x28728, x28729);
  nand n28731(x28731, x28628, x28588);
  nand n28733(x28733, x28633, x28591);
  nand n28735(x28735, x28733, x28734);
  nand n28736(x28736, x28633, x28593);
  nand n28738(x28738, x28638, x28596);
  nand n28740(x28740, x28738, x28739);
  nand n28741(x28741, x28638, x28598);
  nand n28743(x28743, x28643, x28601);
  nand n28745(x28745, x28743, x28744);
  nand n28746(x28746, x28643, x28603);
  nand n28748(x28748, x28648, x28606);
  nand n28750(x28750, x28748, x28749);
  nand n28751(x28751, x28648, x28608);
  nand n28753(x28753, x28653, x28611);
  nand n28755(x28755, x28753, x28754);
  nand n28756(x28756, x28653, x28613);
  nand n28758(x28758, x28658, x28616);
  nand n28760(x28760, x28758, x28759);
  nand n28761(x28761, x28658, x28618);
  nand n28763(x28763, x28663, x28621);
  nand n28765(x28765, x28763, x28764);
  nand n28766(x28766, x28663, x28623);
  nand n28768(x28768, x28668, x28626);
  nand n28770(x28770, x28768, x28769);
  nand n28771(x28771, x28668, x28628);
  nand n28773(x28773, x28673, x28631);
  nand n28775(x28775, x28773, x28774);
  nand n28776(x28776, x28673, x28633);
  nand n28778(x28778, x28678, x28636);
  nand n28780(x28780, x28778, x28779);
  nand n28781(x28781, x28678, x28638);
  nand n28783(x28783, x28683, x28641);
  nand n28785(x28785, x28783, x28784);
  nand n28786(x28786, x28683, x28643);
  nand n28788(x28788, x28688, x28646);
  nand n28790(x28790, x28788, x28789);
  nand n28791(x28791, x28688, x28648);
  nand n28793(x28793, x28693, x28651);
  nand n28795(x28795, x28793, x28794);
  nand n28796(x28796, x28693, x28653);
  nand n28798(x28798, x28722, x71977);
  nand n28800(x28800, x28798, x28799);
  nand n28801(x28801, x28727, x28295);
  nand n28803(x28803, x28801, x28802);
  nand n28804(x28804, x28732, x28418);
  nand n28806(x28806, x28804, x28805);
  nand n28807(x28807, x28737, x28421);
  nand n28809(x28809, x28807, x28808);
  nand n28810(x28810, x28742, x28564);
  nand n28812(x28812, x28810, x28811);
  nand n28813(x28813, x28747, x28567);
  nand n28815(x28815, x28813, x28814);
  nand n28816(x28816, x28752, x28570);
  nand n28818(x28818, x28816, x28817);
  nand n28819(x28819, x28757, x28573);
  nand n28821(x28821, x28819, x28820);
  nand n28822(x28822, x28762, x28696);
  nand n28824(x28824, x28822, x28823);
  nand n28825(x28825, x28767, x28699);
  nand n28827(x28827, x28825, x28826);
  nand n28828(x28828, x28772, x28702);
  nand n28830(x28830, x28828, x28829);
  nand n28831(x28831, x28777, x28705);
  nand n28833(x28833, x28831, x28832);
  nand n28834(x28834, x28782, x28708);
  nand n28836(x28836, x28834, x28835);
  nand n28837(x28837, x28787, x28711);
  nand n28839(x28839, x28837, x28838);
  nand n28840(x28840, x28792, x28714);
  nand n28842(x28842, x28840, x28841);
  nand n28843(x28843, x28797, x28717);
  nand n28845(x28845, x28843, x28844);
  nand n28846(x28846, x28076, x16876);
  nand n28847(x28847, x28846, x28294);
  nand n28849(x28849, x28083, x28295);
  nand n28851(x28851, x28082, x28850);
  nand n28852(x28852, x28851, x28849);
  nand n28854(x28854, x28089, x28418);
  nand n28856(x28856, x28088, x28855);
  nand n28857(x28857, x28856, x28854);
  nand n28859(x28859, x28095, x28421);
  nand n28861(x28861, x28094, x28860);
  nand n28862(x28862, x28861, x28859);
  nand n28864(x28864, x28101, x28564);
  nand n28866(x28866, x28100, x28865);
  nand n28867(x28867, x28866, x28864);
  nand n28869(x28869, x28107, x28567);
  nand n28871(x28871, x28106, x28870);
  nand n28872(x28872, x28871, x28869);
  nand n28874(x28874, x28113, x28570);
  nand n28876(x28876, x28112, x28875);
  nand n28877(x28877, x28876, x28874);
  nand n28879(x28879, x28119, x28573);
  nand n28881(x28881, x28118, x28880);
  nand n28882(x28882, x28881, x28879);
  nand n28884(x28884, x28125, x28696);
  nand n28886(x28886, x28124, x28885);
  nand n28887(x28887, x28886, x28884);
  nand n28889(x28889, x28131, x28699);
  nand n28891(x28891, x28130, x28890);
  nand n28892(x28892, x28891, x28889);
  nand n28894(x28894, x28137, x28702);
  nand n28896(x28896, x28136, x28895);
  nand n28897(x28897, x28896, x28894);
  nand n28899(x28899, x28143, x28705);
  nand n28901(x28901, x28142, x28900);
  nand n28902(x28902, x28901, x28899);
  nand n28904(x28904, x28149, x28708);
  nand n28906(x28906, x28148, x28905);
  nand n28907(x28907, x28906, x28904);
  nand n28909(x28909, x28155, x28711);
  nand n28911(x28911, x28154, x28910);
  nand n28912(x28912, x28911, x28909);
  nand n28914(x28914, x28161, x28714);
  nand n28916(x28916, x28160, x28915);
  nand n28917(x28917, x28916, x28914);
  nand n28919(x28919, x28167, x28717);
  nand n28921(x28921, x28166, x28920);
  nand n28922(x28922, x28921, x28919);
  nand n28924(x28924, x28173, x28800);
  nand n28926(x28926, x28172, x28925);
  nand n28927(x28927, x28926, x28924);
  nand n28929(x28929, x28179, x28803);
  nand n28931(x28931, x28178, x28930);
  nand n28932(x28932, x28931, x28929);
  nand n28934(x28934, x28185, x28806);
  nand n28936(x28936, x28184, x28935);
  nand n28937(x28937, x28936, x28934);
  nand n28939(x28939, x28191, x28809);
  nand n28941(x28941, x28190, x28940);
  nand n28942(x28942, x28941, x28939);
  nand n28944(x28944, x28197, x28812);
  nand n28946(x28946, x28196, x28945);
  nand n28947(x28947, x28946, x28944);
  nand n28949(x28949, x28203, x28815);
  nand n28951(x28951, x28202, x28950);
  nand n28952(x28952, x28951, x28949);
  nand n28954(x28954, x28209, x28818);
  nand n28956(x28956, x28208, x28955);
  nand n28957(x28957, x28956, x28954);
  nand n28959(x28959, x28215, x28821);
  nand n28961(x28961, x28214, x28960);
  nand n28962(x28962, x28961, x28959);
  nand n28964(x28964, x28221, x28824);
  nand n28966(x28966, x28220, x28965);
  nand n28967(x28967, x28966, x28964);
  nand n28969(x28969, x28227, x28827);
  nand n28971(x28971, x28226, x28970);
  nand n28972(x28972, x28971, x28969);
  nand n28974(x28974, x28233, x28830);
  nand n28976(x28976, x28232, x28975);
  nand n28977(x28977, x28976, x28974);
  nand n28979(x28979, x28239, x28833);
  nand n28981(x28981, x28238, x28980);
  nand n28982(x28982, x28981, x28979);
  nand n28984(x28984, x28245, x28836);
  nand n28986(x28986, x28244, x28985);
  nand n28987(x28987, x28986, x28984);
  nand n28989(x28989, x28251, x28839);
  nand n28991(x28991, x28250, x28990);
  nand n28992(x28992, x28991, x28989);
  nand n28994(x28994, x28257, x28842);
  nand n28996(x28996, x28256, x28995);
  nand n28997(x28997, x28996, x28994);
  nand n28999(x28999, x28263, x28845);
  nand n29001(x29001, x28262, x29000);
  nand n29002(x29002, x29001, x28999);
  nand n29004(x29004, x72537, x27881);
  nand n29005(x29005, x72542, x27881);
  nand n29007(x29007, x72537, x27883);
  nand n29009(x29009, x72547, x27881);
  nand n29011(x29011, x72542, x27883);
  nand n29013(x29013, x72537, x27885);
  nand n29015(x29015, x72552, x27881);
  nand n29017(x29017, x72547, x27883);
  nand n29019(x29019, x72542, x27885);
  nand n29021(x29021, x72537, x27887);
  nand n29022(x29022, x72557, x27881);
  nand n29024(x29024, x72552, x27883);
  nand n29026(x29026, x72547, x27885);
  nand n29028(x29028, x72542, x27887);
  nand n29030(x29030, x72537, x27889);
  nand n29032(x29032, x72562, x27881);
  nand n29034(x29034, x72557, x27883);
  nand n29036(x29036, x72552, x27885);
  nand n29038(x29038, x72547, x27887);
  nand n29040(x29040, x72542, x27889);
  nand n29042(x29042, x72537, x27891);
  nand n29044(x29044, x72567, x27881);
  nand n29046(x29046, x72562, x27883);
  nand n29048(x29048, x72557, x27885);
  nand n29050(x29050, x72552, x27887);
  nand n29052(x29052, x72547, x27889);
  nand n29054(x29054, x72542, x27891);
  nand n29056(x29056, x72537, x27893);
  nand n29057(x29057, x72572, x27881);
  nand n29059(x29059, x72567, x27883);
  nand n29061(x29061, x72562, x27885);
  nand n29063(x29063, x72557, x27887);
  nand n29065(x29065, x72552, x27889);
  nand n29067(x29067, x72547, x27891);
  nand n29069(x29069, x72542, x27893);
  nand n29071(x29071, x72537, x27895);
  nand n29073(x29073, x72577, x27881);
  nand n29075(x29075, x72572, x27883);
  nand n29077(x29077, x72567, x27885);
  nand n29079(x29079, x72562, x27887);
  nand n29081(x29081, x72557, x27889);
  nand n29083(x29083, x72552, x27891);
  nand n29085(x29085, x72547, x27893);
  nand n29087(x29087, x72542, x27895);
  nand n29089(x29089, x72537, x27897);
  nand n29091(x29091, x72582, x27881);
  nand n29093(x29093, x72577, x27883);
  nand n29095(x29095, x72572, x27885);
  nand n29097(x29097, x72567, x27887);
  nand n29099(x29099, x72562, x27889);
  nand n29101(x29101, x72557, x27891);
  nand n29103(x29103, x72552, x27893);
  nand n29105(x29105, x72547, x27895);
  nand n29107(x29107, x72542, x27897);
  nand n29109(x29109, x72537, x27899);
  nand n29110(x29110, x72587, x27881);
  nand n29112(x29112, x72582, x27883);
  nand n29114(x29114, x72577, x27885);
  nand n29116(x29116, x72572, x27887);
  nand n29118(x29118, x72567, x27889);
  nand n29120(x29120, x72562, x27891);
  nand n29122(x29122, x72557, x27893);
  nand n29124(x29124, x72552, x27895);
  nand n29126(x29126, x72547, x27897);
  nand n29128(x29128, x72542, x27899);
  nand n29130(x29130, x72537, x27901);
  nand n29132(x29132, x72592, x27881);
  nand n29134(x29134, x72587, x27883);
  nand n29136(x29136, x72582, x27885);
  nand n29138(x29138, x72577, x27887);
  nand n29140(x29140, x72572, x27889);
  nand n29142(x29142, x72567, x27891);
  nand n29144(x29144, x72562, x27893);
  nand n29146(x29146, x72557, x27895);
  nand n29148(x29148, x72552, x27897);
  nand n29150(x29150, x72547, x27899);
  nand n29152(x29152, x72542, x27901);
  nand n29154(x29154, x72537, x27903);
  nand n29156(x29156, x72597, x27881);
  nand n29158(x29158, x72592, x27883);
  nand n29160(x29160, x72587, x27885);
  nand n29162(x29162, x72582, x27887);
  nand n29164(x29164, x72577, x27889);
  nand n29166(x29166, x72572, x27891);
  nand n29168(x29168, x72567, x27893);
  nand n29170(x29170, x72562, x27895);
  nand n29172(x29172, x72557, x27897);
  nand n29174(x29174, x72552, x27899);
  nand n29176(x29176, x72547, x27901);
  nand n29178(x29178, x72542, x27903);
  nand n29180(x29180, x72537, x27905);
  nand n29181(x29181, x72602, x27881);
  nand n29183(x29183, x72597, x27883);
  nand n29185(x29185, x72592, x27885);
  nand n29187(x29187, x72587, x27887);
  nand n29189(x29189, x72582, x27889);
  nand n29191(x29191, x72577, x27891);
  nand n29193(x29193, x72572, x27893);
  nand n29195(x29195, x72567, x27895);
  nand n29197(x29197, x72562, x27897);
  nand n29199(x29199, x72557, x27899);
  nand n29201(x29201, x72552, x27901);
  nand n29203(x29203, x72547, x27903);
  nand n29205(x29205, x72542, x27905);
  nand n29207(x29207, x72537, x27907);
  nand n29209(x29209, x72607, x27881);
  nand n29211(x29211, x72602, x27883);
  nand n29213(x29213, x72597, x27885);
  nand n29215(x29215, x72592, x27887);
  nand n29217(x29217, x72587, x27889);
  nand n29219(x29219, x72582, x27891);
  nand n29221(x29221, x72577, x27893);
  nand n29223(x29223, x72572, x27895);
  nand n29225(x29225, x72567, x27897);
  nand n29227(x29227, x72562, x27899);
  nand n29229(x29229, x72557, x27901);
  nand n29231(x29231, x72552, x27903);
  nand n29233(x29233, x72547, x27905);
  nand n29235(x29235, x72542, x27907);
  nand n29237(x29237, x72537, x27909);
  nand n29239(x29239, x72612, x27881);
  nand n29241(x29241, x72607, x27883);
  nand n29243(x29243, x72602, x27885);
  nand n29245(x29245, x72597, x27887);
  nand n29247(x29247, x72592, x27889);
  nand n29249(x29249, x72587, x27891);
  nand n29251(x29251, x72582, x27893);
  nand n29253(x29253, x72577, x27895);
  nand n29255(x29255, x72572, x27897);
  nand n29257(x29257, x72567, x27899);
  nand n29259(x29259, x72562, x27901);
  nand n29261(x29261, x72557, x27903);
  nand n29263(x29263, x72552, x27905);
  nand n29265(x29265, x72547, x27907);
  nand n29267(x29267, x72542, x27909);
  nand n29269(x29269, x72537, x27911);
  nand n29270(x29270, x72617, x27881);
  nand n29272(x29272, x72612, x27883);
  nand n29274(x29274, x72607, x27885);
  nand n29276(x29276, x72602, x27887);
  nand n29278(x29278, x72597, x27889);
  nand n29280(x29280, x72592, x27891);
  nand n29282(x29282, x72587, x27893);
  nand n29284(x29284, x72582, x27895);
  nand n29286(x29286, x72577, x27897);
  nand n29288(x29288, x72572, x27899);
  nand n29290(x29290, x72567, x27901);
  nand n29292(x29292, x72562, x27903);
  nand n29294(x29294, x72557, x27905);
  nand n29296(x29296, x72552, x27907);
  nand n29298(x29298, x72547, x27909);
  nand n29300(x29300, x72542, x27911);
  nand n29302(x29302, x72537, x27913);
  nand n29304(x29304, x72622, x27881);
  nand n29306(x29306, x72617, x27883);
  nand n29308(x29308, x72612, x27885);
  nand n29310(x29310, x72607, x27887);
  nand n29312(x29312, x72602, x27889);
  nand n29314(x29314, x72597, x27891);
  nand n29316(x29316, x72592, x27893);
  nand n29318(x29318, x72587, x27895);
  nand n29320(x29320, x72582, x27897);
  nand n29322(x29322, x72577, x27899);
  nand n29324(x29324, x72572, x27901);
  nand n29326(x29326, x72567, x27903);
  nand n29328(x29328, x72562, x27905);
  nand n29330(x29330, x72557, x27907);
  nand n29332(x29332, x72552, x27909);
  nand n29334(x29334, x72547, x27911);
  nand n29336(x29336, x72542, x27913);
  nand n29338(x29338, x72537, x27915);
  nand n29340(x29340, x72627, x27881);
  nand n29342(x29342, x72622, x27883);
  nand n29344(x29344, x72617, x27885);
  nand n29346(x29346, x72612, x27887);
  nand n29348(x29348, x72607, x27889);
  nand n29350(x29350, x72602, x27891);
  nand n29352(x29352, x72597, x27893);
  nand n29354(x29354, x72592, x27895);
  nand n29356(x29356, x72587, x27897);
  nand n29358(x29358, x72582, x27899);
  nand n29360(x29360, x72577, x27901);
  nand n29362(x29362, x72572, x27903);
  nand n29364(x29364, x72567, x27905);
  nand n29366(x29366, x72562, x27907);
  nand n29368(x29368, x72557, x27909);
  nand n29370(x29370, x72552, x27911);
  nand n29372(x29372, x72547, x27913);
  nand n29374(x29374, x72542, x27915);
  nand n29376(x29376, x72537, x27917);
  nand n29377(x29377, x72632, x27881);
  nand n29379(x29379, x72627, x27883);
  nand n29381(x29381, x72622, x27885);
  nand n29383(x29383, x72617, x27887);
  nand n29385(x29385, x72612, x27889);
  nand n29387(x29387, x72607, x27891);
  nand n29389(x29389, x72602, x27893);
  nand n29391(x29391, x72597, x27895);
  nand n29393(x29393, x72592, x27897);
  nand n29395(x29395, x72587, x27899);
  nand n29397(x29397, x72582, x27901);
  nand n29399(x29399, x72577, x27903);
  nand n29401(x29401, x72572, x27905);
  nand n29403(x29403, x72567, x27907);
  nand n29405(x29405, x72562, x27909);
  nand n29407(x29407, x72557, x27911);
  nand n29409(x29409, x72552, x27913);
  nand n29411(x29411, x72547, x27915);
  nand n29413(x29413, x72542, x27917);
  nand n29415(x29415, x72537, x27919);
  nand n29417(x29417, x72637, x27881);
  nand n29419(x29419, x72632, x27883);
  nand n29421(x29421, x72627, x27885);
  nand n29423(x29423, x72622, x27887);
  nand n29425(x29425, x72617, x27889);
  nand n29427(x29427, x72612, x27891);
  nand n29429(x29429, x72607, x27893);
  nand n29431(x29431, x72602, x27895);
  nand n29433(x29433, x72597, x27897);
  nand n29435(x29435, x72592, x27899);
  nand n29437(x29437, x72587, x27901);
  nand n29439(x29439, x72582, x27903);
  nand n29441(x29441, x72577, x27905);
  nand n29443(x29443, x72572, x27907);
  nand n29445(x29445, x72567, x27909);
  nand n29447(x29447, x72562, x27911);
  nand n29449(x29449, x72557, x27913);
  nand n29451(x29451, x72552, x27915);
  nand n29453(x29453, x72547, x27917);
  nand n29455(x29455, x72542, x27919);
  nand n29457(x29457, x72537, x27921);
  nand n29459(x29459, x72642, x27881);
  nand n29461(x29461, x72637, x27883);
  nand n29463(x29463, x72632, x27885);
  nand n29465(x29465, x72627, x27887);
  nand n29467(x29467, x72622, x27889);
  nand n29469(x29469, x72617, x27891);
  nand n29471(x29471, x72612, x27893);
  nand n29473(x29473, x72607, x27895);
  nand n29475(x29475, x72602, x27897);
  nand n29477(x29477, x72597, x27899);
  nand n29479(x29479, x72592, x27901);
  nand n29481(x29481, x72587, x27903);
  nand n29483(x29483, x72582, x27905);
  nand n29485(x29485, x72577, x27907);
  nand n29487(x29487, x72572, x27909);
  nand n29489(x29489, x72567, x27911);
  nand n29491(x29491, x72562, x27913);
  nand n29493(x29493, x72557, x27915);
  nand n29495(x29495, x72552, x27917);
  nand n29497(x29497, x72547, x27919);
  nand n29499(x29499, x72542, x27921);
  nand n29501(x29501, x72537, x27923);
  nand n29502(x29502, x72647, x27881);
  nand n29504(x29504, x72642, x27883);
  nand n29506(x29506, x72637, x27885);
  nand n29508(x29508, x72632, x27887);
  nand n29510(x29510, x72627, x27889);
  nand n29512(x29512, x72622, x27891);
  nand n29514(x29514, x72617, x27893);
  nand n29516(x29516, x72612, x27895);
  nand n29518(x29518, x72607, x27897);
  nand n29520(x29520, x72602, x27899);
  nand n29522(x29522, x72597, x27901);
  nand n29524(x29524, x72592, x27903);
  nand n29526(x29526, x72587, x27905);
  nand n29528(x29528, x72582, x27907);
  nand n29530(x29530, x72577, x27909);
  nand n29532(x29532, x72572, x27911);
  nand n29534(x29534, x72567, x27913);
  nand n29536(x29536, x72562, x27915);
  nand n29538(x29538, x72557, x27917);
  nand n29540(x29540, x72552, x27919);
  nand n29542(x29542, x72547, x27921);
  nand n29544(x29544, x72542, x27923);
  nand n29546(x29546, x72537, x27925);
  nand n29548(x29548, x72652, x27881);
  nand n29550(x29550, x72647, x27883);
  nand n29552(x29552, x72642, x27885);
  nand n29554(x29554, x72637, x27887);
  nand n29556(x29556, x72632, x27889);
  nand n29558(x29558, x72627, x27891);
  nand n29560(x29560, x72622, x27893);
  nand n29562(x29562, x72617, x27895);
  nand n29564(x29564, x72612, x27897);
  nand n29566(x29566, x72607, x27899);
  nand n29568(x29568, x72602, x27901);
  nand n29570(x29570, x72597, x27903);
  nand n29572(x29572, x72592, x27905);
  nand n29574(x29574, x72587, x27907);
  nand n29576(x29576, x72582, x27909);
  nand n29578(x29578, x72577, x27911);
  nand n29580(x29580, x72572, x27913);
  nand n29582(x29582, x72567, x27915);
  nand n29584(x29584, x72562, x27917);
  nand n29586(x29586, x72557, x27919);
  nand n29588(x29588, x72552, x27921);
  nand n29590(x29590, x72547, x27923);
  nand n29592(x29592, x72542, x27925);
  nand n29594(x29594, x72537, x27927);
  nand n29596(x29596, x72657, x27881);
  nand n29598(x29598, x72652, x27883);
  nand n29600(x29600, x72647, x27885);
  nand n29602(x29602, x72642, x27887);
  nand n29604(x29604, x72637, x27889);
  nand n29606(x29606, x72632, x27891);
  nand n29608(x29608, x72627, x27893);
  nand n29610(x29610, x72622, x27895);
  nand n29612(x29612, x72617, x27897);
  nand n29614(x29614, x72612, x27899);
  nand n29616(x29616, x72607, x27901);
  nand n29618(x29618, x72602, x27903);
  nand n29620(x29620, x72597, x27905);
  nand n29622(x29622, x72592, x27907);
  nand n29624(x29624, x72587, x27909);
  nand n29626(x29626, x72582, x27911);
  nand n29628(x29628, x72577, x27913);
  nand n29630(x29630, x72572, x27915);
  nand n29632(x29632, x72567, x27917);
  nand n29634(x29634, x72562, x27919);
  nand n29636(x29636, x72557, x27921);
  nand n29638(x29638, x72552, x27923);
  nand n29640(x29640, x72547, x27925);
  nand n29642(x29642, x72542, x27927);
  nand n29644(x29644, x72537, x27929);
  nand n29645(x29645, x72662, x27881);
  nand n29647(x29647, x72657, x27883);
  nand n29649(x29649, x72652, x27885);
  nand n29651(x29651, x72647, x27887);
  nand n29653(x29653, x72642, x27889);
  nand n29655(x29655, x72637, x27891);
  nand n29657(x29657, x72632, x27893);
  nand n29659(x29659, x72627, x27895);
  nand n29661(x29661, x72622, x27897);
  nand n29663(x29663, x72617, x27899);
  nand n29665(x29665, x72612, x27901);
  nand n29667(x29667, x72607, x27903);
  nand n29669(x29669, x72602, x27905);
  nand n29671(x29671, x72597, x27907);
  nand n29673(x29673, x72592, x27909);
  nand n29675(x29675, x72587, x27911);
  nand n29677(x29677, x72582, x27913);
  nand n29679(x29679, x72577, x27915);
  nand n29681(x29681, x72572, x27917);
  nand n29683(x29683, x72567, x27919);
  nand n29685(x29685, x72562, x27921);
  nand n29687(x29687, x72557, x27923);
  nand n29689(x29689, x72552, x27925);
  nand n29691(x29691, x72547, x27927);
  nand n29693(x29693, x72542, x27929);
  nand n29695(x29695, x72537, x27931);
  nand n29697(x29697, x72667, x27881);
  nand n29699(x29699, x72662, x27883);
  nand n29701(x29701, x72657, x27885);
  nand n29703(x29703, x72652, x27887);
  nand n29705(x29705, x72647, x27889);
  nand n29707(x29707, x72642, x27891);
  nand n29709(x29709, x72637, x27893);
  nand n29711(x29711, x72632, x27895);
  nand n29713(x29713, x72627, x27897);
  nand n29715(x29715, x72622, x27899);
  nand n29717(x29717, x72617, x27901);
  nand n29719(x29719, x72612, x27903);
  nand n29721(x29721, x72607, x27905);
  nand n29723(x29723, x72602, x27907);
  nand n29725(x29725, x72597, x27909);
  nand n29727(x29727, x72592, x27911);
  nand n29729(x29729, x72587, x27913);
  nand n29731(x29731, x72582, x27915);
  nand n29733(x29733, x72577, x27917);
  nand n29735(x29735, x72572, x27919);
  nand n29737(x29737, x72567, x27921);
  nand n29739(x29739, x72562, x27923);
  nand n29741(x29741, x72557, x27925);
  nand n29743(x29743, x72552, x27927);
  nand n29745(x29745, x72547, x27929);
  nand n29747(x29747, x72542, x27931);
  nand n29749(x29749, x72537, x27933);
  nand n29751(x29751, x72672, x27881);
  nand n29753(x29753, x72667, x27883);
  nand n29755(x29755, x72662, x27885);
  nand n29757(x29757, x72657, x27887);
  nand n29759(x29759, x72652, x27889);
  nand n29761(x29761, x72647, x27891);
  nand n29763(x29763, x72642, x27893);
  nand n29765(x29765, x72637, x27895);
  nand n29767(x29767, x72632, x27897);
  nand n29769(x29769, x72627, x27899);
  nand n29771(x29771, x72622, x27901);
  nand n29773(x29773, x72617, x27903);
  nand n29775(x29775, x72612, x27905);
  nand n29777(x29777, x72607, x27907);
  nand n29779(x29779, x72602, x27909);
  nand n29781(x29781, x72597, x27911);
  nand n29783(x29783, x72592, x27913);
  nand n29785(x29785, x72587, x27915);
  nand n29787(x29787, x72582, x27917);
  nand n29789(x29789, x72577, x27919);
  nand n29791(x29791, x72572, x27921);
  nand n29793(x29793, x72567, x27923);
  nand n29795(x29795, x72562, x27925);
  nand n29797(x29797, x72557, x27927);
  nand n29799(x29799, x72552, x27929);
  nand n29801(x29801, x72547, x27931);
  nand n29803(x29803, x72542, x27933);
  nand n29805(x29805, x72537, x27935);
  nand n29806(x29806, x72677, x27881);
  nand n29808(x29808, x72672, x27883);
  nand n29810(x29810, x72667, x27885);
  nand n29812(x29812, x72662, x27887);
  nand n29814(x29814, x72657, x27889);
  nand n29816(x29816, x72652, x27891);
  nand n29818(x29818, x72647, x27893);
  nand n29820(x29820, x72642, x27895);
  nand n29822(x29822, x72637, x27897);
  nand n29824(x29824, x72632, x27899);
  nand n29826(x29826, x72627, x27901);
  nand n29828(x29828, x72622, x27903);
  nand n29830(x29830, x72617, x27905);
  nand n29832(x29832, x72612, x27907);
  nand n29834(x29834, x72607, x27909);
  nand n29836(x29836, x72602, x27911);
  nand n29838(x29838, x72597, x27913);
  nand n29840(x29840, x72592, x27915);
  nand n29842(x29842, x72587, x27917);
  nand n29844(x29844, x72582, x27919);
  nand n29846(x29846, x72577, x27921);
  nand n29848(x29848, x72572, x27923);
  nand n29850(x29850, x72567, x27925);
  nand n29852(x29852, x72562, x27927);
  nand n29854(x29854, x72557, x27929);
  nand n29856(x29856, x72552, x27931);
  nand n29858(x29858, x72547, x27933);
  nand n29860(x29860, x72542, x27935);
  nand n29862(x29862, x72537, x27937);
  nand n29864(x29864, x72682, x27881);
  nand n29866(x29866, x72677, x27883);
  nand n29868(x29868, x72672, x27885);
  nand n29870(x29870, x72667, x27887);
  nand n29872(x29872, x72662, x27889);
  nand n29874(x29874, x72657, x27891);
  nand n29876(x29876, x72652, x27893);
  nand n29878(x29878, x72647, x27895);
  nand n29880(x29880, x72642, x27897);
  nand n29882(x29882, x72637, x27899);
  nand n29884(x29884, x72632, x27901);
  nand n29886(x29886, x72627, x27903);
  nand n29888(x29888, x72622, x27905);
  nand n29890(x29890, x72617, x27907);
  nand n29892(x29892, x72612, x27909);
  nand n29894(x29894, x72607, x27911);
  nand n29896(x29896, x72602, x27913);
  nand n29898(x29898, x72597, x27915);
  nand n29900(x29900, x72592, x27917);
  nand n29902(x29902, x72587, x27919);
  nand n29904(x29904, x72582, x27921);
  nand n29906(x29906, x72577, x27923);
  nand n29908(x29908, x72572, x27925);
  nand n29910(x29910, x72567, x27927);
  nand n29912(x29912, x72562, x27929);
  nand n29914(x29914, x72557, x27931);
  nand n29916(x29916, x72552, x27933);
  nand n29918(x29918, x72547, x27935);
  nand n29920(x29920, x72542, x27937);
  nand n29922(x29922, x72537, x27939);
  nand n29924(x29924, x72687, x27881);
  nand n29926(x29926, x72682, x27883);
  nand n29928(x29928, x72677, x27885);
  nand n29930(x29930, x72672, x27887);
  nand n29932(x29932, x72667, x27889);
  nand n29934(x29934, x72662, x27891);
  nand n29936(x29936, x72657, x27893);
  nand n29938(x29938, x72652, x27895);
  nand n29940(x29940, x72647, x27897);
  nand n29942(x29942, x72642, x27899);
  nand n29944(x29944, x72637, x27901);
  nand n29946(x29946, x72632, x27903);
  nand n29948(x29948, x72627, x27905);
  nand n29950(x29950, x72622, x27907);
  nand n29952(x29952, x72617, x27909);
  nand n29954(x29954, x72612, x27911);
  nand n29956(x29956, x72607, x27913);
  nand n29958(x29958, x72602, x27915);
  nand n29960(x29960, x72597, x27917);
  nand n29962(x29962, x72592, x27919);
  nand n29964(x29964, x72587, x27921);
  nand n29966(x29966, x72582, x27923);
  nand n29968(x29968, x72577, x27925);
  nand n29970(x29970, x72572, x27927);
  nand n29972(x29972, x72567, x27929);
  nand n29974(x29974, x72562, x27931);
  nand n29976(x29976, x72557, x27933);
  nand n29978(x29978, x72552, x27935);
  nand n29980(x29980, x72547, x27937);
  nand n29982(x29982, x72542, x27939);
  nand n29984(x29984, x72537, x27941);
  nand n29985(x29985, x72692, x27881);
  nand n29987(x29987, x72687, x27883);
  nand n29989(x29989, x72682, x27885);
  nand n29991(x29991, x72677, x27887);
  nand n29993(x29993, x72672, x27889);
  nand n29995(x29995, x72667, x27891);
  nand n29997(x29997, x72662, x27893);
  nand n29999(x29999, x72657, x27895);
  nand n30001(x30001, x72652, x27897);
  nand n30003(x30003, x72647, x27899);
  nand n30005(x30005, x72642, x27901);
  nand n30007(x30007, x72637, x27903);
  nand n30009(x30009, x72632, x27905);
  nand n30011(x30011, x72627, x27907);
  nand n30013(x30013, x72622, x27909);
  nand n30015(x30015, x72617, x27911);
  nand n30017(x30017, x72612, x27913);
  nand n30019(x30019, x72607, x27915);
  nand n30021(x30021, x72602, x27917);
  nand n30023(x30023, x72597, x27919);
  nand n30025(x30025, x72592, x27921);
  nand n30027(x30027, x72587, x27923);
  nand n30029(x30029, x72582, x27925);
  nand n30031(x30031, x72577, x27927);
  nand n30033(x30033, x72572, x27929);
  nand n30035(x30035, x72567, x27931);
  nand n30037(x30037, x72562, x27933);
  nand n30039(x30039, x72557, x27935);
  nand n30041(x30041, x72552, x27937);
  nand n30043(x30043, x72547, x27939);
  nand n30045(x30045, x72542, x27941);
  nand n30047(x30047, x72537, x27943);
  nand n30049(x30049, x29006, x29008);
  nand n30050(x30050, x29005, x29007);
  nand n30051(x30051, x30050, x30049);
  nand n30052(x30052, x29010, x29012);
  nand n30053(x30053, x29009, x29011);
  nand n30054(x30054, x30053, x30052);
  nand n30056(x30056, x29014, x30055);
  nand n30057(x30057, x29013, x30054);
  nand n30058(x30058, x30057, x30056);
  nand n30059(x30059, x30052, x30056);
  nand n30060(x30060, x29016, x29018);
  nand n30061(x30061, x29015, x29017);
  nand n30062(x30062, x30061, x30060);
  nand n30064(x30064, x29020, x30063);
  nand n30065(x30065, x29019, x30062);
  nand n30066(x30066, x30065, x30064);
  nand n30067(x30067, x30060, x30064);
  nand n30068(x30068, x29023, x29025);
  nand n30069(x30069, x29022, x29024);
  nand n30070(x30070, x30069, x30068);
  nand n30072(x30072, x29027, x30071);
  nand n30073(x30073, x29026, x30070);
  nand n30074(x30074, x30073, x30072);
  nand n30075(x30075, x30068, x30072);
  nand n30076(x30076, x29029, x29031);
  nand n30077(x30077, x29028, x29030);
  nand n30078(x30078, x30077, x30076);
  nand n30079(x30079, x29033, x29035);
  nand n30080(x30080, x29032, x29034);
  nand n30081(x30081, x30080, x30079);
  nand n30083(x30083, x29037, x30082);
  nand n30084(x30084, x29036, x30081);
  nand n30085(x30085, x30084, x30083);
  nand n30086(x30086, x30079, x30083);
  nand n30087(x30087, x29039, x29041);
  nand n30088(x30088, x29038, x29040);
  nand n30089(x30089, x30088, x30087);
  nand n30091(x30091, x29043, x30090);
  nand n30092(x30092, x29042, x30089);
  nand n30093(x30093, x30092, x30091);
  nand n30094(x30094, x30087, x30091);
  nand n30095(x30095, x29045, x29047);
  nand n30096(x30096, x29044, x29046);
  nand n30097(x30097, x30096, x30095);
  nand n30099(x30099, x29049, x30098);
  nand n30100(x30100, x29048, x30097);
  nand n30101(x30101, x30100, x30099);
  nand n30102(x30102, x30095, x30099);
  nand n30103(x30103, x29051, x29053);
  nand n30104(x30104, x29050, x29052);
  nand n30105(x30105, x30104, x30103);
  nand n30107(x30107, x29055, x30106);
  nand n30108(x30108, x29054, x30105);
  nand n30109(x30109, x30108, x30107);
  nand n30111(x30111, x30103, x30107);
  nand n30112(x30112, x29058, x29060);
  nand n30113(x30113, x29057, x29059);
  nand n30114(x30114, x30113, x30112);
  nand n30116(x30116, x29062, x30115);
  nand n30117(x30117, x29061, x30114);
  nand n30118(x30118, x30117, x30116);
  nand n30119(x30119, x30112, x30116);
  nand n30120(x30120, x29064, x29066);
  nand n30121(x30121, x29063, x29065);
  nand n30122(x30122, x30121, x30120);
  nand n30124(x30124, x29068, x30123);
  nand n30125(x30125, x29067, x30122);
  nand n30126(x30126, x30125, x30124);
  nand n30128(x30128, x30120, x30124);
  nand n30129(x30129, x29070, x29072);
  nand n30130(x30130, x29069, x29071);
  nand n30131(x30131, x30130, x30129);
  nand n30132(x30132, x29074, x29076);
  nand n30133(x30133, x29073, x29075);
  nand n30134(x30134, x30133, x30132);
  nand n30136(x30136, x29078, x30135);
  nand n30137(x30137, x29077, x30134);
  nand n30138(x30138, x30137, x30136);
  nand n30139(x30139, x30132, x30136);
  nand n30140(x30140, x29080, x29082);
  nand n30141(x30141, x29079, x29081);
  nand n30142(x30142, x30141, x30140);
  nand n30144(x30144, x29084, x30143);
  nand n30145(x30145, x29083, x30142);
  nand n30146(x30146, x30145, x30144);
  nand n30148(x30148, x30140, x30144);
  nand n30149(x30149, x29086, x29088);
  nand n30150(x30150, x29085, x29087);
  nand n30151(x30151, x30150, x30149);
  nand n30153(x30153, x29090, x30152);
  nand n30154(x30154, x29089, x30151);
  nand n30155(x30155, x30154, x30153);
  nand n30157(x30157, x30149, x30153);
  nand n30158(x30158, x29092, x29094);
  nand n30159(x30159, x29091, x29093);
  nand n30160(x30160, x30159, x30158);
  nand n30162(x30162, x29096, x30161);
  nand n30163(x30163, x29095, x30160);
  nand n30164(x30164, x30163, x30162);
  nand n30165(x30165, x30158, x30162);
  nand n30166(x30166, x29098, x29100);
  nand n30167(x30167, x29097, x29099);
  nand n30168(x30168, x30167, x30166);
  nand n30170(x30170, x29102, x30169);
  nand n30171(x30171, x29101, x30168);
  nand n30172(x30172, x30171, x30170);
  nand n30174(x30174, x30166, x30170);
  nand n30175(x30175, x29104, x29106);
  nand n30176(x30176, x29103, x29105);
  nand n30177(x30177, x30176, x30175);
  nand n30179(x30179, x29108, x30178);
  nand n30180(x30180, x29107, x30177);
  nand n30181(x30181, x30180, x30179);
  nand n30183(x30183, x30175, x30179);
  nand n30184(x30184, x29111, x29113);
  nand n30185(x30185, x29110, x29112);
  nand n30186(x30186, x30185, x30184);
  nand n30188(x30188, x29115, x30187);
  nand n30189(x30189, x29114, x30186);
  nand n30190(x30190, x30189, x30188);
  nand n30191(x30191, x30184, x30188);
  nand n30192(x30192, x29117, x29119);
  nand n30193(x30193, x29116, x29118);
  nand n30194(x30194, x30193, x30192);
  nand n30196(x30196, x29121, x30195);
  nand n30197(x30197, x29120, x30194);
  nand n30198(x30198, x30197, x30196);
  nand n30200(x30200, x30192, x30196);
  nand n30201(x30201, x29123, x29125);
  nand n30202(x30202, x29122, x29124);
  nand n30203(x30203, x30202, x30201);
  nand n30205(x30205, x29127, x30204);
  nand n30206(x30206, x29126, x30203);
  nand n30207(x30207, x30206, x30205);
  nand n30209(x30209, x30201, x30205);
  nand n30210(x30210, x29129, x29131);
  nand n30211(x30211, x29128, x29130);
  nand n30212(x30212, x30211, x30210);
  nand n30213(x30213, x29133, x29135);
  nand n30214(x30214, x29132, x29134);
  nand n30215(x30215, x30214, x30213);
  nand n30217(x30217, x29137, x30216);
  nand n30218(x30218, x29136, x30215);
  nand n30219(x30219, x30218, x30217);
  nand n30220(x30220, x30213, x30217);
  nand n30221(x30221, x29139, x29141);
  nand n30222(x30222, x29138, x29140);
  nand n30223(x30223, x30222, x30221);
  nand n30225(x30225, x29143, x30224);
  nand n30226(x30226, x29142, x30223);
  nand n30227(x30227, x30226, x30225);
  nand n30229(x30229, x30221, x30225);
  nand n30230(x30230, x29145, x29147);
  nand n30231(x30231, x29144, x29146);
  nand n30232(x30232, x30231, x30230);
  nand n30234(x30234, x29149, x30233);
  nand n30235(x30235, x29148, x30232);
  nand n30236(x30236, x30235, x30234);
  nand n30238(x30238, x30230, x30234);
  nand n30239(x30239, x29151, x29153);
  nand n30240(x30240, x29150, x29152);
  nand n30241(x30241, x30240, x30239);
  nand n30243(x30243, x29155, x30242);
  nand n30244(x30244, x29154, x30241);
  nand n30245(x30245, x30244, x30243);
  nand n30247(x30247, x30239, x30243);
  nand n30248(x30248, x29157, x29159);
  nand n30249(x30249, x29156, x29158);
  nand n30250(x30250, x30249, x30248);
  nand n30252(x30252, x29161, x30251);
  nand n30253(x30253, x29160, x30250);
  nand n30254(x30254, x30253, x30252);
  nand n30255(x30255, x30248, x30252);
  nand n30256(x30256, x29163, x29165);
  nand n30257(x30257, x29162, x29164);
  nand n30258(x30258, x30257, x30256);
  nand n30260(x30260, x29167, x30259);
  nand n30261(x30261, x29166, x30258);
  nand n30262(x30262, x30261, x30260);
  nand n30264(x30264, x30256, x30260);
  nand n30265(x30265, x29169, x29171);
  nand n30266(x30266, x29168, x29170);
  nand n30267(x30267, x30266, x30265);
  nand n30269(x30269, x29173, x30268);
  nand n30270(x30270, x29172, x30267);
  nand n30271(x30271, x30270, x30269);
  nand n30273(x30273, x30265, x30269);
  nand n30274(x30274, x29175, x29177);
  nand n30275(x30275, x29174, x29176);
  nand n30276(x30276, x30275, x30274);
  nand n30278(x30278, x29179, x30277);
  nand n30279(x30279, x29178, x30276);
  nand n30280(x30280, x30279, x30278);
  nand n30282(x30282, x30274, x30278);
  nand n30283(x30283, x29182, x29184);
  nand n30284(x30284, x29181, x29183);
  nand n30285(x30285, x30284, x30283);
  nand n30287(x30287, x29186, x30286);
  nand n30288(x30288, x29185, x30285);
  nand n30289(x30289, x30288, x30287);
  nand n30290(x30290, x30283, x30287);
  nand n30291(x30291, x29188, x29190);
  nand n30292(x30292, x29187, x29189);
  nand n30293(x30293, x30292, x30291);
  nand n30295(x30295, x29192, x30294);
  nand n30296(x30296, x29191, x30293);
  nand n30297(x30297, x30296, x30295);
  nand n30299(x30299, x30291, x30295);
  nand n30300(x30300, x29194, x29196);
  nand n30301(x30301, x29193, x29195);
  nand n30302(x30302, x30301, x30300);
  nand n30304(x30304, x29198, x30303);
  nand n30305(x30305, x29197, x30302);
  nand n30306(x30306, x30305, x30304);
  nand n30308(x30308, x30300, x30304);
  nand n30309(x30309, x29200, x29202);
  nand n30310(x30310, x29199, x29201);
  nand n30311(x30311, x30310, x30309);
  nand n30313(x30313, x29204, x30312);
  nand n30314(x30314, x29203, x30311);
  nand n30315(x30315, x30314, x30313);
  nand n30317(x30317, x30309, x30313);
  nand n30318(x30318, x29206, x29208);
  nand n30319(x30319, x29205, x29207);
  nand n30320(x30320, x30319, x30318);
  nand n30321(x30321, x29210, x29212);
  nand n30322(x30322, x29209, x29211);
  nand n30323(x30323, x30322, x30321);
  nand n30325(x30325, x29214, x30324);
  nand n30326(x30326, x29213, x30323);
  nand n30327(x30327, x30326, x30325);
  nand n30328(x30328, x30321, x30325);
  nand n30329(x30329, x29216, x29218);
  nand n30330(x30330, x29215, x29217);
  nand n30331(x30331, x30330, x30329);
  nand n30333(x30333, x29220, x30332);
  nand n30334(x30334, x29219, x30331);
  nand n30335(x30335, x30334, x30333);
  nand n30337(x30337, x30329, x30333);
  nand n30338(x30338, x29222, x29224);
  nand n30339(x30339, x29221, x29223);
  nand n30340(x30340, x30339, x30338);
  nand n30342(x30342, x29226, x30341);
  nand n30343(x30343, x29225, x30340);
  nand n30344(x30344, x30343, x30342);
  nand n30346(x30346, x30338, x30342);
  nand n30347(x30347, x29228, x29230);
  nand n30348(x30348, x29227, x29229);
  nand n30349(x30349, x30348, x30347);
  nand n30351(x30351, x29232, x30350);
  nand n30352(x30352, x29231, x30349);
  nand n30353(x30353, x30352, x30351);
  nand n30355(x30355, x30347, x30351);
  nand n30356(x30356, x29234, x29236);
  nand n30357(x30357, x29233, x29235);
  nand n30358(x30358, x30357, x30356);
  nand n30360(x30360, x29238, x30359);
  nand n30361(x30361, x29237, x30358);
  nand n30362(x30362, x30361, x30360);
  nand n30363(x30363, x30356, x30360);
  nand n30364(x30364, x29240, x29242);
  nand n30365(x30365, x29239, x29241);
  nand n30366(x30366, x30365, x30364);
  nand n30368(x30368, x29244, x30367);
  nand n30369(x30369, x29243, x30366);
  nand n30370(x30370, x30369, x30368);
  nand n30371(x30371, x30364, x30368);
  nand n30372(x30372, x29246, x29248);
  nand n30373(x30373, x29245, x29247);
  nand n30374(x30374, x30373, x30372);
  nand n30376(x30376, x29250, x30375);
  nand n30377(x30377, x29249, x30374);
  nand n30378(x30378, x30377, x30376);
  nand n30380(x30380, x30372, x30376);
  nand n30381(x30381, x29252, x29254);
  nand n30382(x30382, x29251, x29253);
  nand n30383(x30383, x30382, x30381);
  nand n30385(x30385, x29256, x30384);
  nand n30386(x30386, x29255, x30383);
  nand n30387(x30387, x30386, x30385);
  nand n30389(x30389, x30381, x30385);
  nand n30390(x30390, x29258, x29260);
  nand n30391(x30391, x29257, x29259);
  nand n30392(x30392, x30391, x30390);
  nand n30394(x30394, x29262, x30393);
  nand n30395(x30395, x29261, x30392);
  nand n30396(x30396, x30395, x30394);
  nand n30398(x30398, x30390, x30394);
  nand n30399(x30399, x29264, x29266);
  nand n30400(x30400, x29263, x29265);
  nand n30401(x30401, x30400, x30399);
  nand n30403(x30403, x29268, x30402);
  nand n30404(x30404, x29267, x30401);
  nand n30405(x30405, x30404, x30403);
  nand n30407(x30407, x30399, x30403);
  nand n30408(x30408, x29271, x29273);
  nand n30409(x30409, x29270, x29272);
  nand n30410(x30410, x30409, x30408);
  nand n30412(x30412, x29275, x30411);
  nand n30413(x30413, x29274, x30410);
  nand n30414(x30414, x30413, x30412);
  nand n30415(x30415, x30408, x30412);
  nand n30416(x30416, x29277, x29279);
  nand n30417(x30417, x29276, x29278);
  nand n30418(x30418, x30417, x30416);
  nand n30420(x30420, x29281, x30419);
  nand n30421(x30421, x29280, x30418);
  nand n30422(x30422, x30421, x30420);
  nand n30424(x30424, x30416, x30420);
  nand n30425(x30425, x29283, x29285);
  nand n30426(x30426, x29282, x29284);
  nand n30427(x30427, x30426, x30425);
  nand n30429(x30429, x29287, x30428);
  nand n30430(x30430, x29286, x30427);
  nand n30431(x30431, x30430, x30429);
  nand n30433(x30433, x30425, x30429);
  nand n30434(x30434, x29289, x29291);
  nand n30435(x30435, x29288, x29290);
  nand n30436(x30436, x30435, x30434);
  nand n30438(x30438, x29293, x30437);
  nand n30439(x30439, x29292, x30436);
  nand n30440(x30440, x30439, x30438);
  nand n30442(x30442, x30434, x30438);
  nand n30443(x30443, x29295, x29297);
  nand n30444(x30444, x29294, x29296);
  nand n30445(x30445, x30444, x30443);
  nand n30447(x30447, x29299, x30446);
  nand n30448(x30448, x29298, x30445);
  nand n30449(x30449, x30448, x30447);
  nand n30451(x30451, x30443, x30447);
  nand n30452(x30452, x29301, x29303);
  nand n30453(x30453, x29300, x29302);
  nand n30454(x30454, x30453, x30452);
  nand n30455(x30455, x29305, x29307);
  nand n30456(x30456, x29304, x29306);
  nand n30457(x30457, x30456, x30455);
  nand n30459(x30459, x29309, x30458);
  nand n30460(x30460, x29308, x30457);
  nand n30461(x30461, x30460, x30459);
  nand n30462(x30462, x30455, x30459);
  nand n30463(x30463, x29311, x29313);
  nand n30464(x30464, x29310, x29312);
  nand n30465(x30465, x30464, x30463);
  nand n30467(x30467, x29315, x30466);
  nand n30468(x30468, x29314, x30465);
  nand n30469(x30469, x30468, x30467);
  nand n30471(x30471, x30463, x30467);
  nand n30472(x30472, x29317, x29319);
  nand n30473(x30473, x29316, x29318);
  nand n30474(x30474, x30473, x30472);
  nand n30476(x30476, x29321, x30475);
  nand n30477(x30477, x29320, x30474);
  nand n30478(x30478, x30477, x30476);
  nand n30480(x30480, x30472, x30476);
  nand n30481(x30481, x29323, x29325);
  nand n30482(x30482, x29322, x29324);
  nand n30483(x30483, x30482, x30481);
  nand n30485(x30485, x29327, x30484);
  nand n30486(x30486, x29326, x30483);
  nand n30487(x30487, x30486, x30485);
  nand n30489(x30489, x30481, x30485);
  nand n30490(x30490, x29329, x29331);
  nand n30491(x30491, x29328, x29330);
  nand n30492(x30492, x30491, x30490);
  nand n30494(x30494, x29333, x30493);
  nand n30495(x30495, x29332, x30492);
  nand n30496(x30496, x30495, x30494);
  nand n30498(x30498, x30490, x30494);
  nand n30499(x30499, x29335, x29337);
  nand n30500(x30500, x29334, x29336);
  nand n30501(x30501, x30500, x30499);
  nand n30503(x30503, x29339, x30502);
  nand n30504(x30504, x29338, x30501);
  nand n30505(x30505, x30504, x30503);
  nand n30507(x30507, x30499, x30503);
  nand n30508(x30508, x29341, x29343);
  nand n30509(x30509, x29340, x29342);
  nand n30510(x30510, x30509, x30508);
  nand n30512(x30512, x29345, x30511);
  nand n30513(x30513, x29344, x30510);
  nand n30514(x30514, x30513, x30512);
  nand n30515(x30515, x30508, x30512);
  nand n30516(x30516, x29347, x29349);
  nand n30517(x30517, x29346, x29348);
  nand n30518(x30518, x30517, x30516);
  nand n30520(x30520, x29351, x30519);
  nand n30521(x30521, x29350, x30518);
  nand n30522(x30522, x30521, x30520);
  nand n30524(x30524, x30516, x30520);
  nand n30525(x30525, x29353, x29355);
  nand n30526(x30526, x29352, x29354);
  nand n30527(x30527, x30526, x30525);
  nand n30529(x30529, x29357, x30528);
  nand n30530(x30530, x29356, x30527);
  nand n30531(x30531, x30530, x30529);
  nand n30533(x30533, x30525, x30529);
  nand n30534(x30534, x29359, x29361);
  nand n30535(x30535, x29358, x29360);
  nand n30536(x30536, x30535, x30534);
  nand n30538(x30538, x29363, x30537);
  nand n30539(x30539, x29362, x30536);
  nand n30540(x30540, x30539, x30538);
  nand n30542(x30542, x30534, x30538);
  nand n30543(x30543, x29365, x29367);
  nand n30544(x30544, x29364, x29366);
  nand n30545(x30545, x30544, x30543);
  nand n30547(x30547, x29369, x30546);
  nand n30548(x30548, x29368, x30545);
  nand n30549(x30549, x30548, x30547);
  nand n30551(x30551, x30543, x30547);
  nand n30552(x30552, x29371, x29373);
  nand n30553(x30553, x29370, x29372);
  nand n30554(x30554, x30553, x30552);
  nand n30556(x30556, x29375, x30555);
  nand n30557(x30557, x29374, x30554);
  nand n30558(x30558, x30557, x30556);
  nand n30560(x30560, x30552, x30556);
  nand n30561(x30561, x29378, x29380);
  nand n30562(x30562, x29377, x29379);
  nand n30563(x30563, x30562, x30561);
  nand n30565(x30565, x29382, x30564);
  nand n30566(x30566, x29381, x30563);
  nand n30567(x30567, x30566, x30565);
  nand n30568(x30568, x30561, x30565);
  nand n30569(x30569, x29384, x29386);
  nand n30570(x30570, x29383, x29385);
  nand n30571(x30571, x30570, x30569);
  nand n30573(x30573, x29388, x30572);
  nand n30574(x30574, x29387, x30571);
  nand n30575(x30575, x30574, x30573);
  nand n30577(x30577, x30569, x30573);
  nand n30578(x30578, x29390, x29392);
  nand n30579(x30579, x29389, x29391);
  nand n30580(x30580, x30579, x30578);
  nand n30582(x30582, x29394, x30581);
  nand n30583(x30583, x29393, x30580);
  nand n30584(x30584, x30583, x30582);
  nand n30586(x30586, x30578, x30582);
  nand n30587(x30587, x29396, x29398);
  nand n30588(x30588, x29395, x29397);
  nand n30589(x30589, x30588, x30587);
  nand n30591(x30591, x29400, x30590);
  nand n30592(x30592, x29399, x30589);
  nand n30593(x30593, x30592, x30591);
  nand n30595(x30595, x30587, x30591);
  nand n30596(x30596, x29402, x29404);
  nand n30597(x30597, x29401, x29403);
  nand n30598(x30598, x30597, x30596);
  nand n30600(x30600, x29406, x30599);
  nand n30601(x30601, x29405, x30598);
  nand n30602(x30602, x30601, x30600);
  nand n30604(x30604, x30596, x30600);
  nand n30605(x30605, x29408, x29410);
  nand n30606(x30606, x29407, x29409);
  nand n30607(x30607, x30606, x30605);
  nand n30609(x30609, x29412, x30608);
  nand n30610(x30610, x29411, x30607);
  nand n30611(x30611, x30610, x30609);
  nand n30613(x30613, x30605, x30609);
  nand n30614(x30614, x29414, x29416);
  nand n30615(x30615, x29413, x29415);
  nand n30616(x30616, x30615, x30614);
  nand n30617(x30617, x29418, x29420);
  nand n30618(x30618, x29417, x29419);
  nand n30619(x30619, x30618, x30617);
  nand n30621(x30621, x29422, x30620);
  nand n30622(x30622, x29421, x30619);
  nand n30623(x30623, x30622, x30621);
  nand n30624(x30624, x30617, x30621);
  nand n30625(x30625, x29424, x29426);
  nand n30626(x30626, x29423, x29425);
  nand n30627(x30627, x30626, x30625);
  nand n30629(x30629, x29428, x30628);
  nand n30630(x30630, x29427, x30627);
  nand n30631(x30631, x30630, x30629);
  nand n30633(x30633, x30625, x30629);
  nand n30634(x30634, x29430, x29432);
  nand n30635(x30635, x29429, x29431);
  nand n30636(x30636, x30635, x30634);
  nand n30638(x30638, x29434, x30637);
  nand n30639(x30639, x29433, x30636);
  nand n30640(x30640, x30639, x30638);
  nand n30642(x30642, x30634, x30638);
  nand n30643(x30643, x29436, x29438);
  nand n30644(x30644, x29435, x29437);
  nand n30645(x30645, x30644, x30643);
  nand n30647(x30647, x29440, x30646);
  nand n30648(x30648, x29439, x30645);
  nand n30649(x30649, x30648, x30647);
  nand n30651(x30651, x30643, x30647);
  nand n30652(x30652, x29442, x29444);
  nand n30653(x30653, x29441, x29443);
  nand n30654(x30654, x30653, x30652);
  nand n30656(x30656, x29446, x30655);
  nand n30657(x30657, x29445, x30654);
  nand n30658(x30658, x30657, x30656);
  nand n30660(x30660, x30652, x30656);
  nand n30661(x30661, x29448, x29450);
  nand n30662(x30662, x29447, x29449);
  nand n30663(x30663, x30662, x30661);
  nand n30665(x30665, x29452, x30664);
  nand n30666(x30666, x29451, x30663);
  nand n30667(x30667, x30666, x30665);
  nand n30669(x30669, x30661, x30665);
  nand n30670(x30670, x29454, x29456);
  nand n30671(x30671, x29453, x29455);
  nand n30672(x30672, x30671, x30670);
  nand n30674(x30674, x29458, x30673);
  nand n30675(x30675, x29457, x30672);
  nand n30676(x30676, x30675, x30674);
  nand n30678(x30678, x30670, x30674);
  nand n30679(x30679, x29460, x29462);
  nand n30680(x30680, x29459, x29461);
  nand n30681(x30681, x30680, x30679);
  nand n30683(x30683, x29464, x30682);
  nand n30684(x30684, x29463, x30681);
  nand n30685(x30685, x30684, x30683);
  nand n30686(x30686, x30679, x30683);
  nand n30687(x30687, x29466, x29468);
  nand n30688(x30688, x29465, x29467);
  nand n30689(x30689, x30688, x30687);
  nand n30691(x30691, x29470, x30690);
  nand n30692(x30692, x29469, x30689);
  nand n30693(x30693, x30692, x30691);
  nand n30695(x30695, x30687, x30691);
  nand n30696(x30696, x29472, x29474);
  nand n30697(x30697, x29471, x29473);
  nand n30698(x30698, x30697, x30696);
  nand n30700(x30700, x29476, x30699);
  nand n30701(x30701, x29475, x30698);
  nand n30702(x30702, x30701, x30700);
  nand n30704(x30704, x30696, x30700);
  nand n30705(x30705, x29478, x29480);
  nand n30706(x30706, x29477, x29479);
  nand n30707(x30707, x30706, x30705);
  nand n30709(x30709, x29482, x30708);
  nand n30710(x30710, x29481, x30707);
  nand n30711(x30711, x30710, x30709);
  nand n30713(x30713, x30705, x30709);
  nand n30714(x30714, x29484, x29486);
  nand n30715(x30715, x29483, x29485);
  nand n30716(x30716, x30715, x30714);
  nand n30718(x30718, x29488, x30717);
  nand n30719(x30719, x29487, x30716);
  nand n30720(x30720, x30719, x30718);
  nand n30722(x30722, x30714, x30718);
  nand n30723(x30723, x29490, x29492);
  nand n30724(x30724, x29489, x29491);
  nand n30725(x30725, x30724, x30723);
  nand n30727(x30727, x29494, x30726);
  nand n30728(x30728, x29493, x30725);
  nand n30729(x30729, x30728, x30727);
  nand n30731(x30731, x30723, x30727);
  nand n30732(x30732, x29496, x29498);
  nand n30733(x30733, x29495, x29497);
  nand n30734(x30734, x30733, x30732);
  nand n30736(x30736, x29500, x30735);
  nand n30737(x30737, x29499, x30734);
  nand n30738(x30738, x30737, x30736);
  nand n30740(x30740, x30732, x30736);
  nand n30741(x30741, x29503, x29505);
  nand n30742(x30742, x29502, x29504);
  nand n30743(x30743, x30742, x30741);
  nand n30745(x30745, x29507, x30744);
  nand n30746(x30746, x29506, x30743);
  nand n30747(x30747, x30746, x30745);
  nand n30748(x30748, x30741, x30745);
  nand n30749(x30749, x29509, x29511);
  nand n30750(x30750, x29508, x29510);
  nand n30751(x30751, x30750, x30749);
  nand n30753(x30753, x29513, x30752);
  nand n30754(x30754, x29512, x30751);
  nand n30755(x30755, x30754, x30753);
  nand n30757(x30757, x30749, x30753);
  nand n30758(x30758, x29515, x29517);
  nand n30759(x30759, x29514, x29516);
  nand n30760(x30760, x30759, x30758);
  nand n30762(x30762, x29519, x30761);
  nand n30763(x30763, x29518, x30760);
  nand n30764(x30764, x30763, x30762);
  nand n30766(x30766, x30758, x30762);
  nand n30767(x30767, x29521, x29523);
  nand n30768(x30768, x29520, x29522);
  nand n30769(x30769, x30768, x30767);
  nand n30771(x30771, x29525, x30770);
  nand n30772(x30772, x29524, x30769);
  nand n30773(x30773, x30772, x30771);
  nand n30775(x30775, x30767, x30771);
  nand n30776(x30776, x29527, x29529);
  nand n30777(x30777, x29526, x29528);
  nand n30778(x30778, x30777, x30776);
  nand n30780(x30780, x29531, x30779);
  nand n30781(x30781, x29530, x30778);
  nand n30782(x30782, x30781, x30780);
  nand n30784(x30784, x30776, x30780);
  nand n30785(x30785, x29533, x29535);
  nand n30786(x30786, x29532, x29534);
  nand n30787(x30787, x30786, x30785);
  nand n30789(x30789, x29537, x30788);
  nand n30790(x30790, x29536, x30787);
  nand n30791(x30791, x30790, x30789);
  nand n30793(x30793, x30785, x30789);
  nand n30794(x30794, x29539, x29541);
  nand n30795(x30795, x29538, x29540);
  nand n30796(x30796, x30795, x30794);
  nand n30798(x30798, x29543, x30797);
  nand n30799(x30799, x29542, x30796);
  nand n30800(x30800, x30799, x30798);
  nand n30802(x30802, x30794, x30798);
  nand n30803(x30803, x29545, x29547);
  nand n30804(x30804, x29544, x29546);
  nand n30805(x30805, x30804, x30803);
  nand n30806(x30806, x29549, x29551);
  nand n30807(x30807, x29548, x29550);
  nand n30808(x30808, x30807, x30806);
  nand n30810(x30810, x29553, x30809);
  nand n30811(x30811, x29552, x30808);
  nand n30812(x30812, x30811, x30810);
  nand n30813(x30813, x30806, x30810);
  nand n30814(x30814, x29555, x29557);
  nand n30815(x30815, x29554, x29556);
  nand n30816(x30816, x30815, x30814);
  nand n30818(x30818, x29559, x30817);
  nand n30819(x30819, x29558, x30816);
  nand n30820(x30820, x30819, x30818);
  nand n30822(x30822, x30814, x30818);
  nand n30823(x30823, x29561, x29563);
  nand n30824(x30824, x29560, x29562);
  nand n30825(x30825, x30824, x30823);
  nand n30827(x30827, x29565, x30826);
  nand n30828(x30828, x29564, x30825);
  nand n30829(x30829, x30828, x30827);
  nand n30831(x30831, x30823, x30827);
  nand n30832(x30832, x29567, x29569);
  nand n30833(x30833, x29566, x29568);
  nand n30834(x30834, x30833, x30832);
  nand n30836(x30836, x29571, x30835);
  nand n30837(x30837, x29570, x30834);
  nand n30838(x30838, x30837, x30836);
  nand n30840(x30840, x30832, x30836);
  nand n30841(x30841, x29573, x29575);
  nand n30842(x30842, x29572, x29574);
  nand n30843(x30843, x30842, x30841);
  nand n30845(x30845, x29577, x30844);
  nand n30846(x30846, x29576, x30843);
  nand n30847(x30847, x30846, x30845);
  nand n30849(x30849, x30841, x30845);
  nand n30850(x30850, x29579, x29581);
  nand n30851(x30851, x29578, x29580);
  nand n30852(x30852, x30851, x30850);
  nand n30854(x30854, x29583, x30853);
  nand n30855(x30855, x29582, x30852);
  nand n30856(x30856, x30855, x30854);
  nand n30858(x30858, x30850, x30854);
  nand n30859(x30859, x29585, x29587);
  nand n30860(x30860, x29584, x29586);
  nand n30861(x30861, x30860, x30859);
  nand n30863(x30863, x29589, x30862);
  nand n30864(x30864, x29588, x30861);
  nand n30865(x30865, x30864, x30863);
  nand n30867(x30867, x30859, x30863);
  nand n30868(x30868, x29591, x29593);
  nand n30869(x30869, x29590, x29592);
  nand n30870(x30870, x30869, x30868);
  nand n30872(x30872, x29595, x30871);
  nand n30873(x30873, x29594, x30870);
  nand n30874(x30874, x30873, x30872);
  nand n30875(x30875, x30868, x30872);
  nand n30876(x30876, x29597, x29599);
  nand n30877(x30877, x29596, x29598);
  nand n30878(x30878, x30877, x30876);
  nand n30880(x30880, x29601, x30879);
  nand n30881(x30881, x29600, x30878);
  nand n30882(x30882, x30881, x30880);
  nand n30883(x30883, x30876, x30880);
  nand n30884(x30884, x29603, x29605);
  nand n30885(x30885, x29602, x29604);
  nand n30886(x30886, x30885, x30884);
  nand n30888(x30888, x29607, x30887);
  nand n30889(x30889, x29606, x30886);
  nand n30890(x30890, x30889, x30888);
  nand n30892(x30892, x30884, x30888);
  nand n30893(x30893, x29609, x29611);
  nand n30894(x30894, x29608, x29610);
  nand n30895(x30895, x30894, x30893);
  nand n30897(x30897, x29613, x30896);
  nand n30898(x30898, x29612, x30895);
  nand n30899(x30899, x30898, x30897);
  nand n30901(x30901, x30893, x30897);
  nand n30902(x30902, x29615, x29617);
  nand n30903(x30903, x29614, x29616);
  nand n30904(x30904, x30903, x30902);
  nand n30906(x30906, x29619, x30905);
  nand n30907(x30907, x29618, x30904);
  nand n30908(x30908, x30907, x30906);
  nand n30910(x30910, x30902, x30906);
  nand n30911(x30911, x29621, x29623);
  nand n30912(x30912, x29620, x29622);
  nand n30913(x30913, x30912, x30911);
  nand n30915(x30915, x29625, x30914);
  nand n30916(x30916, x29624, x30913);
  nand n30917(x30917, x30916, x30915);
  nand n30919(x30919, x30911, x30915);
  nand n30920(x30920, x29627, x29629);
  nand n30921(x30921, x29626, x29628);
  nand n30922(x30922, x30921, x30920);
  nand n30924(x30924, x29631, x30923);
  nand n30925(x30925, x29630, x30922);
  nand n30926(x30926, x30925, x30924);
  nand n30928(x30928, x30920, x30924);
  nand n30929(x30929, x29633, x29635);
  nand n30930(x30930, x29632, x29634);
  nand n30931(x30931, x30930, x30929);
  nand n30933(x30933, x29637, x30932);
  nand n30934(x30934, x29636, x30931);
  nand n30935(x30935, x30934, x30933);
  nand n30937(x30937, x30929, x30933);
  nand n30938(x30938, x29639, x29641);
  nand n30939(x30939, x29638, x29640);
  nand n30940(x30940, x30939, x30938);
  nand n30942(x30942, x29643, x30941);
  nand n30943(x30943, x29642, x30940);
  nand n30944(x30944, x30943, x30942);
  nand n30946(x30946, x30938, x30942);
  nand n30947(x30947, x29646, x29648);
  nand n30948(x30948, x29645, x29647);
  nand n30949(x30949, x30948, x30947);
  nand n30951(x30951, x29650, x30950);
  nand n30952(x30952, x29649, x30949);
  nand n30953(x30953, x30952, x30951);
  nand n30954(x30954, x30947, x30951);
  nand n30955(x30955, x29652, x29654);
  nand n30956(x30956, x29651, x29653);
  nand n30957(x30957, x30956, x30955);
  nand n30959(x30959, x29656, x30958);
  nand n30960(x30960, x29655, x30957);
  nand n30961(x30961, x30960, x30959);
  nand n30963(x30963, x30955, x30959);
  nand n30964(x30964, x29658, x29660);
  nand n30965(x30965, x29657, x29659);
  nand n30966(x30966, x30965, x30964);
  nand n30968(x30968, x29662, x30967);
  nand n30969(x30969, x29661, x30966);
  nand n30970(x30970, x30969, x30968);
  nand n30972(x30972, x30964, x30968);
  nand n30973(x30973, x29664, x29666);
  nand n30974(x30974, x29663, x29665);
  nand n30975(x30975, x30974, x30973);
  nand n30977(x30977, x29668, x30976);
  nand n30978(x30978, x29667, x30975);
  nand n30979(x30979, x30978, x30977);
  nand n30981(x30981, x30973, x30977);
  nand n30982(x30982, x29670, x29672);
  nand n30983(x30983, x29669, x29671);
  nand n30984(x30984, x30983, x30982);
  nand n30986(x30986, x29674, x30985);
  nand n30987(x30987, x29673, x30984);
  nand n30988(x30988, x30987, x30986);
  nand n30990(x30990, x30982, x30986);
  nand n30991(x30991, x29676, x29678);
  nand n30992(x30992, x29675, x29677);
  nand n30993(x30993, x30992, x30991);
  nand n30995(x30995, x29680, x30994);
  nand n30996(x30996, x29679, x30993);
  nand n30997(x30997, x30996, x30995);
  nand n30999(x30999, x30991, x30995);
  nand n31000(x31000, x29682, x29684);
  nand n31001(x31001, x29681, x29683);
  nand n31002(x31002, x31001, x31000);
  nand n31004(x31004, x29686, x31003);
  nand n31005(x31005, x29685, x31002);
  nand n31006(x31006, x31005, x31004);
  nand n31008(x31008, x31000, x31004);
  nand n31009(x31009, x29688, x29690);
  nand n31010(x31010, x29687, x29689);
  nand n31011(x31011, x31010, x31009);
  nand n31013(x31013, x29692, x31012);
  nand n31014(x31014, x29691, x31011);
  nand n31015(x31015, x31014, x31013);
  nand n31017(x31017, x31009, x31013);
  nand n31018(x31018, x29694, x29696);
  nand n31019(x31019, x29693, x29695);
  nand n31020(x31020, x31019, x31018);
  nand n31021(x31021, x29698, x29700);
  nand n31022(x31022, x29697, x29699);
  nand n31023(x31023, x31022, x31021);
  nand n31025(x31025, x29702, x31024);
  nand n31026(x31026, x29701, x31023);
  nand n31027(x31027, x31026, x31025);
  nand n31028(x31028, x31021, x31025);
  nand n31029(x31029, x29704, x29706);
  nand n31030(x31030, x29703, x29705);
  nand n31031(x31031, x31030, x31029);
  nand n31033(x31033, x29708, x31032);
  nand n31034(x31034, x29707, x31031);
  nand n31035(x31035, x31034, x31033);
  nand n31037(x31037, x31029, x31033);
  nand n31038(x31038, x29710, x29712);
  nand n31039(x31039, x29709, x29711);
  nand n31040(x31040, x31039, x31038);
  nand n31042(x31042, x29714, x31041);
  nand n31043(x31043, x29713, x31040);
  nand n31044(x31044, x31043, x31042);
  nand n31046(x31046, x31038, x31042);
  nand n31047(x31047, x29716, x29718);
  nand n31048(x31048, x29715, x29717);
  nand n31049(x31049, x31048, x31047);
  nand n31051(x31051, x29720, x31050);
  nand n31052(x31052, x29719, x31049);
  nand n31053(x31053, x31052, x31051);
  nand n31055(x31055, x31047, x31051);
  nand n31056(x31056, x29722, x29724);
  nand n31057(x31057, x29721, x29723);
  nand n31058(x31058, x31057, x31056);
  nand n31060(x31060, x29726, x31059);
  nand n31061(x31061, x29725, x31058);
  nand n31062(x31062, x31061, x31060);
  nand n31064(x31064, x31056, x31060);
  nand n31065(x31065, x29728, x29730);
  nand n31066(x31066, x29727, x29729);
  nand n31067(x31067, x31066, x31065);
  nand n31069(x31069, x29732, x31068);
  nand n31070(x31070, x29731, x31067);
  nand n31071(x31071, x31070, x31069);
  nand n31073(x31073, x31065, x31069);
  nand n31074(x31074, x29734, x29736);
  nand n31075(x31075, x29733, x29735);
  nand n31076(x31076, x31075, x31074);
  nand n31078(x31078, x29738, x31077);
  nand n31079(x31079, x29737, x31076);
  nand n31080(x31080, x31079, x31078);
  nand n31082(x31082, x31074, x31078);
  nand n31083(x31083, x29740, x29742);
  nand n31084(x31084, x29739, x29741);
  nand n31085(x31085, x31084, x31083);
  nand n31087(x31087, x29744, x31086);
  nand n31088(x31088, x29743, x31085);
  nand n31089(x31089, x31088, x31087);
  nand n31091(x31091, x31083, x31087);
  nand n31092(x31092, x29746, x29748);
  nand n31093(x31093, x29745, x29747);
  nand n31094(x31094, x31093, x31092);
  nand n31096(x31096, x29750, x31095);
  nand n31097(x31097, x29749, x31094);
  nand n31098(x31098, x31097, x31096);
  nand n31100(x31100, x31092, x31096);
  nand n31101(x31101, x29752, x29754);
  nand n31102(x31102, x29751, x29753);
  nand n31103(x31103, x31102, x31101);
  nand n31105(x31105, x29756, x31104);
  nand n31106(x31106, x29755, x31103);
  nand n31107(x31107, x31106, x31105);
  nand n31108(x31108, x31101, x31105);
  nand n31109(x31109, x29758, x29760);
  nand n31110(x31110, x29757, x29759);
  nand n31111(x31111, x31110, x31109);
  nand n31113(x31113, x29762, x31112);
  nand n31114(x31114, x29761, x31111);
  nand n31115(x31115, x31114, x31113);
  nand n31117(x31117, x31109, x31113);
  nand n31118(x31118, x29764, x29766);
  nand n31119(x31119, x29763, x29765);
  nand n31120(x31120, x31119, x31118);
  nand n31122(x31122, x29768, x31121);
  nand n31123(x31123, x29767, x31120);
  nand n31124(x31124, x31123, x31122);
  nand n31126(x31126, x31118, x31122);
  nand n31127(x31127, x29770, x29772);
  nand n31128(x31128, x29769, x29771);
  nand n31129(x31129, x31128, x31127);
  nand n31131(x31131, x29774, x31130);
  nand n31132(x31132, x29773, x31129);
  nand n31133(x31133, x31132, x31131);
  nand n31135(x31135, x31127, x31131);
  nand n31136(x31136, x29776, x29778);
  nand n31137(x31137, x29775, x29777);
  nand n31138(x31138, x31137, x31136);
  nand n31140(x31140, x29780, x31139);
  nand n31141(x31141, x29779, x31138);
  nand n31142(x31142, x31141, x31140);
  nand n31144(x31144, x31136, x31140);
  nand n31145(x31145, x29782, x29784);
  nand n31146(x31146, x29781, x29783);
  nand n31147(x31147, x31146, x31145);
  nand n31149(x31149, x29786, x31148);
  nand n31150(x31150, x29785, x31147);
  nand n31151(x31151, x31150, x31149);
  nand n31153(x31153, x31145, x31149);
  nand n31154(x31154, x29788, x29790);
  nand n31155(x31155, x29787, x29789);
  nand n31156(x31156, x31155, x31154);
  nand n31158(x31158, x29792, x31157);
  nand n31159(x31159, x29791, x31156);
  nand n31160(x31160, x31159, x31158);
  nand n31162(x31162, x31154, x31158);
  nand n31163(x31163, x29794, x29796);
  nand n31164(x31164, x29793, x29795);
  nand n31165(x31165, x31164, x31163);
  nand n31167(x31167, x29798, x31166);
  nand n31168(x31168, x29797, x31165);
  nand n31169(x31169, x31168, x31167);
  nand n31171(x31171, x31163, x31167);
  nand n31172(x31172, x29800, x29802);
  nand n31173(x31173, x29799, x29801);
  nand n31174(x31174, x31173, x31172);
  nand n31176(x31176, x29804, x31175);
  nand n31177(x31177, x29803, x31174);
  nand n31178(x31178, x31177, x31176);
  nand n31180(x31180, x31172, x31176);
  nand n31181(x31181, x29807, x29809);
  nand n31182(x31182, x29806, x29808);
  nand n31183(x31183, x31182, x31181);
  nand n31185(x31185, x29811, x31184);
  nand n31186(x31186, x29810, x31183);
  nand n31187(x31187, x31186, x31185);
  nand n31188(x31188, x31181, x31185);
  nand n31189(x31189, x29813, x29815);
  nand n31190(x31190, x29812, x29814);
  nand n31191(x31191, x31190, x31189);
  nand n31193(x31193, x29817, x31192);
  nand n31194(x31194, x29816, x31191);
  nand n31195(x31195, x31194, x31193);
  nand n31197(x31197, x31189, x31193);
  nand n31198(x31198, x29819, x29821);
  nand n31199(x31199, x29818, x29820);
  nand n31200(x31200, x31199, x31198);
  nand n31202(x31202, x29823, x31201);
  nand n31203(x31203, x29822, x31200);
  nand n31204(x31204, x31203, x31202);
  nand n31206(x31206, x31198, x31202);
  nand n31207(x31207, x29825, x29827);
  nand n31208(x31208, x29824, x29826);
  nand n31209(x31209, x31208, x31207);
  nand n31211(x31211, x29829, x31210);
  nand n31212(x31212, x29828, x31209);
  nand n31213(x31213, x31212, x31211);
  nand n31215(x31215, x31207, x31211);
  nand n31216(x31216, x29831, x29833);
  nand n31217(x31217, x29830, x29832);
  nand n31218(x31218, x31217, x31216);
  nand n31220(x31220, x29835, x31219);
  nand n31221(x31221, x29834, x31218);
  nand n31222(x31222, x31221, x31220);
  nand n31224(x31224, x31216, x31220);
  nand n31225(x31225, x29837, x29839);
  nand n31226(x31226, x29836, x29838);
  nand n31227(x31227, x31226, x31225);
  nand n31229(x31229, x29841, x31228);
  nand n31230(x31230, x29840, x31227);
  nand n31231(x31231, x31230, x31229);
  nand n31233(x31233, x31225, x31229);
  nand n31234(x31234, x29843, x29845);
  nand n31235(x31235, x29842, x29844);
  nand n31236(x31236, x31235, x31234);
  nand n31238(x31238, x29847, x31237);
  nand n31239(x31239, x29846, x31236);
  nand n31240(x31240, x31239, x31238);
  nand n31242(x31242, x31234, x31238);
  nand n31243(x31243, x29849, x29851);
  nand n31244(x31244, x29848, x29850);
  nand n31245(x31245, x31244, x31243);
  nand n31247(x31247, x29853, x31246);
  nand n31248(x31248, x29852, x31245);
  nand n31249(x31249, x31248, x31247);
  nand n31251(x31251, x31243, x31247);
  nand n31252(x31252, x29855, x29857);
  nand n31253(x31253, x29854, x29856);
  nand n31254(x31254, x31253, x31252);
  nand n31256(x31256, x29859, x31255);
  nand n31257(x31257, x29858, x31254);
  nand n31258(x31258, x31257, x31256);
  nand n31260(x31260, x31252, x31256);
  nand n31261(x31261, x29861, x29863);
  nand n31262(x31262, x29860, x29862);
  nand n31263(x31263, x31262, x31261);
  nand n31264(x31264, x29865, x29867);
  nand n31265(x31265, x29864, x29866);
  nand n31266(x31266, x31265, x31264);
  nand n31268(x31268, x29869, x31267);
  nand n31269(x31269, x29868, x31266);
  nand n31270(x31270, x31269, x31268);
  nand n31272(x31272, x31264, x31268);
  nand n31273(x31273, x29871, x29873);
  nand n31274(x31274, x29870, x29872);
  nand n31275(x31275, x31274, x31273);
  nand n31277(x31277, x29875, x31276);
  nand n31278(x31278, x29874, x31275);
  nand n31279(x31279, x31278, x31277);
  nand n31281(x31281, x31273, x31277);
  nand n31282(x31282, x29877, x29879);
  nand n31283(x31283, x29876, x29878);
  nand n31284(x31284, x31283, x31282);
  nand n31286(x31286, x29881, x31285);
  nand n31287(x31287, x29880, x31284);
  nand n31288(x31288, x31287, x31286);
  nand n31290(x31290, x31282, x31286);
  nand n31291(x31291, x29883, x29885);
  nand n31292(x31292, x29882, x29884);
  nand n31293(x31293, x31292, x31291);
  nand n31295(x31295, x29887, x31294);
  nand n31296(x31296, x29886, x31293);
  nand n31297(x31297, x31296, x31295);
  nand n31299(x31299, x31291, x31295);
  nand n31300(x31300, x29889, x29891);
  nand n31301(x31301, x29888, x29890);
  nand n31302(x31302, x31301, x31300);
  nand n31304(x31304, x29893, x31303);
  nand n31305(x31305, x29892, x31302);
  nand n31306(x31306, x31305, x31304);
  nand n31308(x31308, x31300, x31304);
  nand n31309(x31309, x29895, x29897);
  nand n31310(x31310, x29894, x29896);
  nand n31311(x31311, x31310, x31309);
  nand n31313(x31313, x29899, x31312);
  nand n31314(x31314, x29898, x31311);
  nand n31315(x31315, x31314, x31313);
  nand n31317(x31317, x31309, x31313);
  nand n31318(x31318, x29901, x29903);
  nand n31319(x31319, x29900, x29902);
  nand n31320(x31320, x31319, x31318);
  nand n31322(x31322, x29905, x31321);
  nand n31323(x31323, x29904, x31320);
  nand n31324(x31324, x31323, x31322);
  nand n31326(x31326, x31318, x31322);
  nand n31327(x31327, x29907, x29909);
  nand n31328(x31328, x29906, x29908);
  nand n31329(x31329, x31328, x31327);
  nand n31331(x31331, x29911, x31330);
  nand n31332(x31332, x29910, x31329);
  nand n31333(x31333, x31332, x31331);
  nand n31335(x31335, x31327, x31331);
  nand n31336(x31336, x29913, x29915);
  nand n31337(x31337, x29912, x29914);
  nand n31338(x31338, x31337, x31336);
  nand n31340(x31340, x29917, x31339);
  nand n31341(x31341, x29916, x31338);
  nand n31342(x31342, x31341, x31340);
  nand n31344(x31344, x31336, x31340);
  nand n31345(x31345, x29919, x29921);
  nand n31346(x31346, x29918, x29920);
  nand n31347(x31347, x31346, x31345);
  nand n31349(x31349, x29923, x31348);
  nand n31350(x31350, x29922, x31347);
  nand n31351(x31351, x31350, x31349);
  nand n31353(x31353, x31345, x31349);
  nand n31354(x31354, x29925, x29927);
  nand n31355(x31355, x29924, x29926);
  nand n31356(x31356, x31355, x31354);
  nand n31358(x31358, x29929, x31357);
  nand n31359(x31359, x29928, x31356);
  nand n31360(x31360, x31359, x31358);
  nand n31362(x31362, x31354, x31358);
  nand n31363(x31363, x29931, x29933);
  nand n31364(x31364, x29930, x29932);
  nand n31365(x31365, x31364, x31363);
  nand n31367(x31367, x29935, x31366);
  nand n31368(x31368, x29934, x31365);
  nand n31369(x31369, x31368, x31367);
  nand n31371(x31371, x31363, x31367);
  nand n31372(x31372, x29937, x29939);
  nand n31373(x31373, x29936, x29938);
  nand n31374(x31374, x31373, x31372);
  nand n31376(x31376, x29941, x31375);
  nand n31377(x31377, x29940, x31374);
  nand n31378(x31378, x31377, x31376);
  nand n31380(x31380, x31372, x31376);
  nand n31381(x31381, x29943, x29945);
  nand n31382(x31382, x29942, x29944);
  nand n31383(x31383, x31382, x31381);
  nand n31385(x31385, x29947, x31384);
  nand n31386(x31386, x29946, x31383);
  nand n31387(x31387, x31386, x31385);
  nand n31389(x31389, x31381, x31385);
  nand n31390(x31390, x29949, x29951);
  nand n31391(x31391, x29948, x29950);
  nand n31392(x31392, x31391, x31390);
  nand n31394(x31394, x29953, x31393);
  nand n31395(x31395, x29952, x31392);
  nand n31396(x31396, x31395, x31394);
  nand n31398(x31398, x31390, x31394);
  nand n31399(x31399, x29955, x29957);
  nand n31400(x31400, x29954, x29956);
  nand n31401(x31401, x31400, x31399);
  nand n31403(x31403, x29959, x31402);
  nand n31404(x31404, x29958, x31401);
  nand n31405(x31405, x31404, x31403);
  nand n31407(x31407, x31399, x31403);
  nand n31408(x31408, x29961, x29963);
  nand n31409(x31409, x29960, x29962);
  nand n31410(x31410, x31409, x31408);
  nand n31412(x31412, x29965, x31411);
  nand n31413(x31413, x29964, x31410);
  nand n31414(x31414, x31413, x31412);
  nand n31416(x31416, x31408, x31412);
  nand n31417(x31417, x29967, x29969);
  nand n31418(x31418, x29966, x29968);
  nand n31419(x31419, x31418, x31417);
  nand n31421(x31421, x29971, x31420);
  nand n31422(x31422, x29970, x31419);
  nand n31423(x31423, x31422, x31421);
  nand n31425(x31425, x31417, x31421);
  nand n31426(x31426, x29973, x29975);
  nand n31427(x31427, x29972, x29974);
  nand n31428(x31428, x31427, x31426);
  nand n31430(x31430, x29977, x31429);
  nand n31431(x31431, x29976, x31428);
  nand n31432(x31432, x31431, x31430);
  nand n31434(x31434, x31426, x31430);
  nand n31435(x31435, x29979, x29981);
  nand n31436(x31436, x29978, x29980);
  nand n31437(x31437, x31436, x31435);
  nand n31439(x31439, x29983, x31438);
  nand n31440(x31440, x29982, x31437);
  nand n31441(x31441, x31440, x31439);
  nand n31443(x31443, x31435, x31439);
  nand n31444(x31444, x29986, x29988);
  nand n31445(x31445, x29985, x29987);
  nand n31446(x31446, x31445, x31444);
  nand n31448(x31448, x29990, x31447);
  nand n31449(x31449, x29989, x31446);
  nand n31450(x31450, x31449, x31448);
  nand n31452(x31452, x29992, x29994);
  nand n31453(x31453, x29991, x29993);
  nand n31454(x31454, x31453, x31452);
  nand n31456(x31456, x29996, x31455);
  nand n31457(x31457, x29995, x31454);
  nand n31458(x31458, x31457, x31456);
  nand n31460(x31460, x29998, x30000);
  nand n31461(x31461, x29997, x29999);
  nand n31462(x31462, x31461, x31460);
  nand n31464(x31464, x30002, x31463);
  nand n31465(x31465, x30001, x31462);
  nand n31466(x31466, x31465, x31464);
  nand n31468(x31468, x30004, x30006);
  nand n31469(x31469, x30003, x30005);
  nand n31470(x31470, x31469, x31468);
  nand n31472(x31472, x30008, x31471);
  nand n31473(x31473, x30007, x31470);
  nand n31474(x31474, x31473, x31472);
  nand n31476(x31476, x30010, x30012);
  nand n31477(x31477, x30009, x30011);
  nand n31478(x31478, x31477, x31476);
  nand n31480(x31480, x30014, x31479);
  nand n31481(x31481, x30013, x31478);
  nand n31482(x31482, x31481, x31480);
  nand n31484(x31484, x30016, x30018);
  nand n31485(x31485, x30015, x30017);
  nand n31486(x31486, x31485, x31484);
  nand n31488(x31488, x30020, x31487);
  nand n31489(x31489, x30019, x31486);
  nand n31490(x31490, x31489, x31488);
  nand n31492(x31492, x30022, x30024);
  nand n31493(x31493, x30021, x30023);
  nand n31494(x31494, x31493, x31492);
  nand n31496(x31496, x30026, x31495);
  nand n31497(x31497, x30025, x31494);
  nand n31498(x31498, x31497, x31496);
  nand n31500(x31500, x30028, x30030);
  nand n31501(x31501, x30027, x30029);
  nand n31502(x31502, x31501, x31500);
  nand n31504(x31504, x30032, x31503);
  nand n31505(x31505, x30031, x31502);
  nand n31506(x31506, x31505, x31504);
  nand n31508(x31508, x30034, x30036);
  nand n31509(x31509, x30033, x30035);
  nand n31510(x31510, x31509, x31508);
  nand n31512(x31512, x30038, x31511);
  nand n31513(x31513, x30037, x31510);
  nand n31514(x31514, x31513, x31512);
  nand n31516(x31516, x30040, x30042);
  nand n31517(x31517, x30039, x30041);
  nand n31518(x31518, x31517, x31516);
  nand n31520(x31520, x30044, x31519);
  nand n31521(x31521, x30043, x31518);
  nand n31522(x31522, x31521, x31520);
  nand n31524(x31524, x30046, x30048);
  nand n31525(x31525, x30045, x30047);
  nand n31526(x31526, x31525, x31524);
  nand n31530(x31530, x30075, x84289);
  nand n31532(x31532, x31531, x30076);
  nand n31533(x31533, x31532, x31530);
  nand n31534(x31534, x30086, x30094);
  nand n31537(x31537, x31536, x31535);
  nand n31538(x31538, x31537, x31534);
  nand n31539(x31539, x30110, x84290);
  nand n31540(x31540, x30109, x29056);
  nand n31541(x31541, x31540, x31539);
  nand n31542(x31542, x30102, x30111);
  nand n31545(x31545, x31544, x31543);
  nand n31546(x31546, x31545, x31542);
  nand n31547(x31547, x30127, x84291);
  nand n31548(x31548, x30126, x30131);
  nand n31549(x31549, x31548, x31547);
  nand n31550(x31550, x30119, x30128);
  nand n31553(x31553, x31552, x31551);
  nand n31554(x31554, x31553, x31550);
  nand n31556(x31556, x84292, x31555);
  nand n31557(x31557, x30129, x31554);
  nand n31558(x31558, x31557, x31556);
  nand n31559(x31559, x31550, x31556);
  nand n31560(x31560, x30147, x30156);
  nand n31561(x31561, x30146, x30155);
  nand n31562(x31562, x31561, x31560);
  nand n31563(x31563, x30139, x30148);
  nand n31566(x31566, x31565, x31564);
  nand n31567(x31567, x31566, x31563);
  nand n31569(x31569, x30157, x31568);
  nand n31571(x31571, x31570, x31567);
  nand n31572(x31572, x31571, x31569);
  nand n31573(x31573, x31563, x31569);
  nand n31574(x31574, x30173, x30182);
  nand n31575(x31575, x30172, x30181);
  nand n31576(x31576, x31575, x31574);
  nand n31578(x31578, x84293, x31577);
  nand n31579(x31579, x29109, x31576);
  nand n31580(x31580, x31579, x31578);
  nand n31582(x31582, x31574, x31578);
  nand n31583(x31583, x30165, x30174);
  nand n31586(x31586, x31585, x31584);
  nand n31587(x31587, x31586, x31583);
  nand n31589(x31589, x30183, x31588);
  nand n31591(x31591, x31590, x31587);
  nand n31592(x31592, x31591, x31589);
  nand n31593(x31593, x31583, x31589);
  nand n31594(x31594, x30199, x30208);
  nand n31595(x31595, x30198, x30207);
  nand n31596(x31596, x31595, x31594);
  nand n31598(x31598, x84294, x31597);
  nand n31599(x31599, x30212, x31596);
  nand n31600(x31600, x31599, x31598);
  nand n31602(x31602, x31594, x31598);
  nand n31603(x31603, x30191, x30200);
  nand n31606(x31606, x31605, x31604);
  nand n31607(x31607, x31606, x31603);
  nand n31609(x31609, x30209, x31608);
  nand n31611(x31611, x31610, x31607);
  nand n31612(x31612, x31611, x31609);
  nand n31613(x31613, x31603, x31609);
  nand n31614(x31614, x30228, x30237);
  nand n31615(x31615, x30227, x30236);
  nand n31616(x31616, x31615, x31614);
  nand n31618(x31618, x30246, x31617);
  nand n31619(x31619, x30245, x31616);
  nand n31620(x31620, x31619, x31618);
  nand n31622(x31622, x31614, x31618);
  nand n31623(x31623, x30220, x30229);
  nand n31626(x31626, x31625, x31624);
  nand n31627(x31627, x31626, x31623);
  nand n31629(x31629, x30238, x31628);
  nand n31631(x31631, x31630, x31627);
  nand n31632(x31632, x31631, x31629);
  nand n31633(x31633, x31623, x31629);
  nand n31635(x31635, x30263, x30272);
  nand n31636(x31636, x30262, x30271);
  nand n31637(x31637, x31636, x31635);
  nand n31639(x31639, x30281, x31638);
  nand n31640(x31640, x30280, x31637);
  nand n31641(x31641, x31640, x31639);
  nand n31643(x31643, x31635, x31639);
  nand n31644(x31644, x30255, x30264);
  nand n31647(x31647, x31646, x31645);
  nand n31648(x31648, x31647, x31644);
  nand n31650(x31650, x30273, x31649);
  nand n31652(x31652, x31651, x31648);
  nand n31653(x31653, x31652, x31650);
  nand n31654(x31654, x31644, x31650);
  nand n31656(x31656, x30298, x30307);
  nand n31657(x31657, x30297, x30306);
  nand n31658(x31658, x31657, x31656);
  nand n31660(x31660, x30316, x31659);
  nand n31661(x31661, x30315, x31658);
  nand n31662(x31662, x31661, x31660);
  nand n31664(x31664, x31656, x31660);
  nand n31665(x31665, x30290, x30299);
  nand n31668(x31668, x31667, x31666);
  nand n31669(x31669, x31668, x31665);
  nand n31671(x31671, x30308, x31670);
  nand n31673(x31673, x31672, x31669);
  nand n31674(x31674, x31673, x31671);
  nand n31675(x31675, x31665, x31671);
  nand n31676(x31676, x30317, x84295);
  nand n31678(x31678, x31677, x30318);
  nand n31679(x31679, x31678, x31676);
  nand n31680(x31680, x30336, x30345);
  nand n31681(x31681, x30335, x30344);
  nand n31682(x31682, x31681, x31680);
  nand n31684(x31684, x30354, x31683);
  nand n31685(x31685, x30353, x31682);
  nand n31686(x31686, x31685, x31684);
  nand n31688(x31688, x31680, x31684);
  nand n31689(x31689, x30328, x30337);
  nand n31692(x31692, x31691, x31690);
  nand n31693(x31693, x31692, x31689);
  nand n31695(x31695, x30346, x31694);
  nand n31697(x31697, x31696, x31693);
  nand n31698(x31698, x31697, x31695);
  nand n31699(x31699, x31689, x31695);
  nand n31700(x31700, x30355, x30363);
  nand n31703(x31703, x31702, x31701);
  nand n31704(x31704, x31703, x31700);
  nand n31705(x31705, x30379, x30388);
  nand n31706(x31706, x30378, x30387);
  nand n31707(x31707, x31706, x31705);
  nand n31709(x31709, x30397, x31708);
  nand n31710(x31710, x30396, x31707);
  nand n31711(x31711, x31710, x31709);
  nand n31713(x31713, x31705, x31709);
  nand n31714(x31714, x30406, x84296);
  nand n31715(x31715, x30405, x29269);
  nand n31716(x31716, x31715, x31714);
  nand n31717(x31717, x30371, x30380);
  nand n31720(x31720, x31719, x31718);
  nand n31721(x31721, x31720, x31717);
  nand n31723(x31723, x30389, x31722);
  nand n31725(x31725, x31724, x31721);
  nand n31726(x31726, x31725, x31723);
  nand n31727(x31727, x31717, x31723);
  nand n31728(x31728, x30398, x30407);
  nand n31731(x31731, x31730, x31729);
  nand n31732(x31732, x31731, x31728);
  nand n31733(x31733, x30423, x30432);
  nand n31734(x31734, x30422, x30431);
  nand n31735(x31735, x31734, x31733);
  nand n31737(x31737, x30441, x31736);
  nand n31738(x31738, x30440, x31735);
  nand n31739(x31739, x31738, x31737);
  nand n31741(x31741, x31733, x31737);
  nand n31742(x31742, x30450, x84297);
  nand n31743(x31743, x30449, x30454);
  nand n31744(x31744, x31743, x31742);
  nand n31745(x31745, x30415, x30424);
  nand n31748(x31748, x31747, x31746);
  nand n31749(x31749, x31748, x31745);
  nand n31751(x31751, x30433, x31750);
  nand n31753(x31753, x31752, x31749);
  nand n31754(x31754, x31753, x31751);
  nand n31755(x31755, x31745, x31751);
  nand n31756(x31756, x30442, x30451);
  nand n31759(x31759, x31758, x31757);
  nand n31760(x31760, x31759, x31756);
  nand n31762(x31762, x84298, x31761);
  nand n31763(x31763, x30452, x31760);
  nand n31764(x31764, x31763, x31762);
  nand n31766(x31766, x31756, x31762);
  nand n31767(x31767, x30470, x30479);
  nand n31768(x31768, x30469, x30478);
  nand n31769(x31769, x31768, x31767);
  nand n31771(x31771, x30488, x31770);
  nand n31772(x31772, x30487, x31769);
  nand n31773(x31773, x31772, x31771);
  nand n31775(x31775, x31767, x31771);
  nand n31776(x31776, x30497, x30506);
  nand n31777(x31777, x30496, x30505);
  nand n31778(x31778, x31777, x31776);
  nand n31779(x31779, x30462, x30471);
  nand n31782(x31782, x31781, x31780);
  nand n31783(x31783, x31782, x31779);
  nand n31785(x31785, x30480, x31784);
  nand n31787(x31787, x31786, x31783);
  nand n31788(x31788, x31787, x31785);
  nand n31789(x31789, x31779, x31785);
  nand n31790(x31790, x30489, x30498);
  nand n31793(x31793, x31792, x31791);
  nand n31794(x31794, x31793, x31790);
  nand n31796(x31796, x30507, x31795);
  nand n31798(x31798, x31797, x31794);
  nand n31799(x31799, x31798, x31796);
  nand n31801(x31801, x31790, x31796);
  nand n31802(x31802, x30523, x30532);
  nand n31803(x31803, x30522, x30531);
  nand n31804(x31804, x31803, x31802);
  nand n31806(x31806, x30541, x31805);
  nand n31807(x31807, x30540, x31804);
  nand n31808(x31808, x31807, x31806);
  nand n31810(x31810, x31802, x31806);
  nand n31811(x31811, x30550, x30559);
  nand n31812(x31812, x30549, x30558);
  nand n31813(x31813, x31812, x31811);
  nand n31815(x31815, x84299, x31814);
  nand n31816(x31816, x29376, x31813);
  nand n31817(x31817, x31816, x31815);
  nand n31818(x31818, x31811, x31815);
  nand n31819(x31819, x30515, x30524);
  nand n31822(x31822, x31821, x31820);
  nand n31823(x31823, x31822, x31819);
  nand n31825(x31825, x30533, x31824);
  nand n31827(x31827, x31826, x31823);
  nand n31828(x31828, x31827, x31825);
  nand n31829(x31829, x31819, x31825);
  nand n31830(x31830, x30542, x30551);
  nand n31833(x31833, x31832, x31831);
  nand n31834(x31834, x31833, x31830);
  nand n31836(x31836, x30560, x31835);
  nand n31838(x31838, x31837, x31834);
  nand n31839(x31839, x31838, x31836);
  nand n31841(x31841, x31830, x31836);
  nand n31842(x31842, x30576, x30585);
  nand n31843(x31843, x30575, x30584);
  nand n31844(x31844, x31843, x31842);
  nand n31846(x31846, x30594, x31845);
  nand n31847(x31847, x30593, x31844);
  nand n31848(x31848, x31847, x31846);
  nand n31850(x31850, x31842, x31846);
  nand n31851(x31851, x30603, x30612);
  nand n31852(x31852, x30602, x30611);
  nand n31853(x31853, x31852, x31851);
  nand n31855(x31855, x84300, x31854);
  nand n31856(x31856, x30616, x31853);
  nand n31857(x31857, x31856, x31855);
  nand n31858(x31858, x31851, x31855);
  nand n31859(x31859, x30568, x30577);
  nand n31862(x31862, x31861, x31860);
  nand n31863(x31863, x31862, x31859);
  nand n31865(x31865, x30586, x31864);
  nand n31867(x31867, x31866, x31863);
  nand n31868(x31868, x31867, x31865);
  nand n31869(x31869, x31859, x31865);
  nand n31870(x31870, x30595, x30604);
  nand n31873(x31873, x31872, x31871);
  nand n31874(x31874, x31873, x31870);
  nand n31876(x31876, x30613, x31875);
  nand n31878(x31878, x31877, x31874);
  nand n31879(x31879, x31878, x31876);
  nand n31881(x31881, x31870, x31876);
  nand n31882(x31882, x30632, x30641);
  nand n31883(x31883, x30631, x30640);
  nand n31884(x31884, x31883, x31882);
  nand n31886(x31886, x30650, x31885);
  nand n31887(x31887, x30649, x31884);
  nand n31888(x31888, x31887, x31886);
  nand n31890(x31890, x31882, x31886);
  nand n31891(x31891, x30659, x30668);
  nand n31892(x31892, x30658, x30667);
  nand n31893(x31893, x31892, x31891);
  nand n31895(x31895, x30677, x31894);
  nand n31896(x31896, x30676, x31893);
  nand n31897(x31897, x31896, x31895);
  nand n31898(x31898, x31891, x31895);
  nand n31899(x31899, x30624, x30633);
  nand n31902(x31902, x31901, x31900);
  nand n31903(x31903, x31902, x31899);
  nand n31905(x31905, x30642, x31904);
  nand n31907(x31907, x31906, x31903);
  nand n31908(x31908, x31907, x31905);
  nand n31909(x31909, x31899, x31905);
  nand n31910(x31910, x30651, x30660);
  nand n31913(x31913, x31912, x31911);
  nand n31914(x31914, x31913, x31910);
  nand n31916(x31916, x30669, x31915);
  nand n31918(x31918, x31917, x31914);
  nand n31919(x31919, x31918, x31916);
  nand n31921(x31921, x31910, x31916);
  nand n31923(x31923, x30694, x30703);
  nand n31924(x31924, x30693, x30702);
  nand n31925(x31925, x31924, x31923);
  nand n31927(x31927, x30712, x31926);
  nand n31928(x31928, x30711, x31925);
  nand n31929(x31929, x31928, x31927);
  nand n31931(x31931, x31923, x31927);
  nand n31932(x31932, x30721, x30730);
  nand n31933(x31933, x30720, x30729);
  nand n31934(x31934, x31933, x31932);
  nand n31936(x31936, x30739, x31935);
  nand n31937(x31937, x30738, x31934);
  nand n31938(x31938, x31937, x31936);
  nand n31940(x31940, x31932, x31936);
  nand n31941(x31941, x30686, x30695);
  nand n31944(x31944, x31943, x31942);
  nand n31945(x31945, x31944, x31941);
  nand n31947(x31947, x30704, x31946);
  nand n31949(x31949, x31948, x31945);
  nand n31950(x31950, x31949, x31947);
  nand n31951(x31951, x31941, x31947);
  nand n31952(x31952, x30713, x30722);
  nand n31955(x31955, x31954, x31953);
  nand n31956(x31956, x31955, x31952);
  nand n31958(x31958, x30731, x31957);
  nand n31960(x31960, x31959, x31956);
  nand n31961(x31961, x31960, x31958);
  nand n31963(x31963, x31952, x31958);
  nand n31965(x31965, x30756, x30765);
  nand n31966(x31966, x30755, x30764);
  nand n31967(x31967, x31966, x31965);
  nand n31969(x31969, x30774, x31968);
  nand n31970(x31970, x30773, x31967);
  nand n31971(x31971, x31970, x31969);
  nand n31973(x31973, x31965, x31969);
  nand n31974(x31974, x30783, x30792);
  nand n31975(x31975, x30782, x30791);
  nand n31976(x31976, x31975, x31974);
  nand n31978(x31978, x30801, x31977);
  nand n31979(x31979, x30800, x31976);
  nand n31980(x31980, x31979, x31978);
  nand n31982(x31982, x31974, x31978);
  nand n31983(x31983, x30748, x30757);
  nand n31986(x31986, x31985, x31984);
  nand n31987(x31987, x31986, x31983);
  nand n31989(x31989, x30766, x31988);
  nand n31991(x31991, x31990, x31987);
  nand n31992(x31992, x31991, x31989);
  nand n31993(x31993, x31983, x31989);
  nand n31994(x31994, x30775, x30784);
  nand n31997(x31997, x31996, x31995);
  nand n31998(x31998, x31997, x31994);
  nand n32000(x32000, x30793, x31999);
  nand n32002(x32002, x32001, x31998);
  nand n32003(x32003, x32002, x32000);
  nand n32005(x32005, x31994, x32000);
  nand n32006(x32006, x30802, x84301);
  nand n32008(x32008, x32007, x30803);
  nand n32009(x32009, x32008, x32006);
  nand n32010(x32010, x30821, x30830);
  nand n32011(x32011, x30820, x30829);
  nand n32012(x32012, x32011, x32010);
  nand n32014(x32014, x30839, x32013);
  nand n32015(x32015, x30838, x32012);
  nand n32016(x32016, x32015, x32014);
  nand n32018(x32018, x32010, x32014);
  nand n32019(x32019, x30848, x30857);
  nand n32020(x32020, x30847, x30856);
  nand n32021(x32021, x32020, x32019);
  nand n32023(x32023, x30866, x32022);
  nand n32024(x32024, x30865, x32021);
  nand n32025(x32025, x32024, x32023);
  nand n32027(x32027, x32019, x32023);
  nand n32028(x32028, x30813, x30822);
  nand n32031(x32031, x32030, x32029);
  nand n32032(x32032, x32031, x32028);
  nand n32034(x32034, x30831, x32033);
  nand n32036(x32036, x32035, x32032);
  nand n32037(x32037, x32036, x32034);
  nand n32038(x32038, x32028, x32034);
  nand n32039(x32039, x30840, x30849);
  nand n32042(x32042, x32041, x32040);
  nand n32043(x32043, x32042, x32039);
  nand n32045(x32045, x30858, x32044);
  nand n32047(x32047, x32046, x32043);
  nand n32048(x32048, x32047, x32045);
  nand n32050(x32050, x32039, x32045);
  nand n32051(x32051, x30867, x30875);
  nand n32054(x32054, x32053, x32052);
  nand n32055(x32055, x32054, x32051);
  nand n32056(x32056, x30891, x30900);
  nand n32057(x32057, x30890, x30899);
  nand n32058(x32058, x32057, x32056);
  nand n32060(x32060, x30909, x32059);
  nand n32061(x32061, x30908, x32058);
  nand n32062(x32062, x32061, x32060);
  nand n32064(x32064, x32056, x32060);
  nand n32065(x32065, x30918, x30927);
  nand n32066(x32066, x30917, x30926);
  nand n32067(x32067, x32066, x32065);
  nand n32069(x32069, x30936, x32068);
  nand n32070(x32070, x30935, x32067);
  nand n32071(x32071, x32070, x32069);
  nand n32073(x32073, x32065, x32069);
  nand n32074(x32074, x30945, x84302);
  nand n32075(x32075, x30944, x29644);
  nand n32076(x32076, x32075, x32074);
  nand n32077(x32077, x30883, x30892);
  nand n32080(x32080, x32079, x32078);
  nand n32081(x32081, x32080, x32077);
  nand n32083(x32083, x30901, x32082);
  nand n32085(x32085, x32084, x32081);
  nand n32086(x32086, x32085, x32083);
  nand n32088(x32088, x32077, x32083);
  nand n32089(x32089, x30910, x30919);
  nand n32092(x32092, x32091, x32090);
  nand n32093(x32093, x32092, x32089);
  nand n32095(x32095, x30928, x32094);
  nand n32097(x32097, x32096, x32093);
  nand n32098(x32098, x32097, x32095);
  nand n32100(x32100, x32089, x32095);
  nand n32101(x32101, x30937, x30946);
  nand n32104(x32104, x32103, x32102);
  nand n32105(x32105, x32104, x32101);
  nand n32106(x32106, x30962, x30971);
  nand n32107(x32107, x30961, x30970);
  nand n32108(x32108, x32107, x32106);
  nand n32110(x32110, x30980, x32109);
  nand n32111(x32111, x30979, x32108);
  nand n32112(x32112, x32111, x32110);
  nand n32114(x32114, x32106, x32110);
  nand n32115(x32115, x30989, x30998);
  nand n32116(x32116, x30988, x30997);
  nand n32117(x32117, x32116, x32115);
  nand n32119(x32119, x31007, x32118);
  nand n32120(x32120, x31006, x32117);
  nand n32121(x32121, x32120, x32119);
  nand n32123(x32123, x32115, x32119);
  nand n32124(x32124, x31016, x84303);
  nand n32125(x32125, x31015, x31020);
  nand n32126(x32126, x32125, x32124);
  nand n32127(x32127, x30954, x30963);
  nand n32130(x32130, x32129, x32128);
  nand n32131(x32131, x32130, x32127);
  nand n32133(x32133, x30972, x32132);
  nand n32135(x32135, x32134, x32131);
  nand n32136(x32136, x32135, x32133);
  nand n32138(x32138, x32127, x32133);
  nand n32139(x32139, x30981, x30990);
  nand n32142(x32142, x32141, x32140);
  nand n32143(x32143, x32142, x32139);
  nand n32145(x32145, x30999, x32144);
  nand n32147(x32147, x32146, x32143);
  nand n32148(x32148, x32147, x32145);
  nand n32150(x32150, x32139, x32145);
  nand n32151(x32151, x31008, x31017);
  nand n32154(x32154, x32153, x32152);
  nand n32155(x32155, x32154, x32151);
  nand n32157(x32157, x84304, x32156);
  nand n32158(x32158, x31018, x32155);
  nand n32159(x32159, x32158, x32157);
  nand n32161(x32161, x32151, x32157);
  nand n32162(x32162, x31036, x31045);
  nand n32163(x32163, x31035, x31044);
  nand n32164(x32164, x32163, x32162);
  nand n32166(x32166, x31054, x32165);
  nand n32167(x32167, x31053, x32164);
  nand n32168(x32168, x32167, x32166);
  nand n32170(x32170, x32162, x32166);
  nand n32171(x32171, x31063, x31072);
  nand n32172(x32172, x31062, x31071);
  nand n32173(x32173, x32172, x32171);
  nand n32175(x32175, x31081, x32174);
  nand n32176(x32176, x31080, x32173);
  nand n32177(x32177, x32176, x32175);
  nand n32179(x32179, x32171, x32175);
  nand n32180(x32180, x31090, x31099);
  nand n32181(x32181, x31089, x31098);
  nand n32182(x32182, x32181, x32180);
  nand n32183(x32183, x31028, x31037);
  nand n32186(x32186, x32185, x32184);
  nand n32187(x32187, x32186, x32183);
  nand n32189(x32189, x31046, x32188);
  nand n32191(x32191, x32190, x32187);
  nand n32192(x32192, x32191, x32189);
  nand n32194(x32194, x32183, x32189);
  nand n32195(x32195, x31055, x31064);
  nand n32198(x32198, x32197, x32196);
  nand n32199(x32199, x32198, x32195);
  nand n32201(x32201, x31073, x32200);
  nand n32203(x32203, x32202, x32199);
  nand n32204(x32204, x32203, x32201);
  nand n32206(x32206, x32195, x32201);
  nand n32207(x32207, x31082, x31091);
  nand n32210(x32210, x32209, x32208);
  nand n32211(x32211, x32210, x32207);
  nand n32213(x32213, x31100, x32212);
  nand n32215(x32215, x32214, x32211);
  nand n32216(x32216, x32215, x32213);
  nand n32218(x32218, x32207, x32213);
  nand n32219(x32219, x31116, x31125);
  nand n32220(x32220, x31115, x31124);
  nand n32221(x32221, x32220, x32219);
  nand n32223(x32223, x31134, x32222);
  nand n32224(x32224, x31133, x32221);
  nand n32225(x32225, x32224, x32223);
  nand n32227(x32227, x32219, x32223);
  nand n32228(x32228, x31143, x31152);
  nand n32229(x32229, x31142, x31151);
  nand n32230(x32230, x32229, x32228);
  nand n32232(x32232, x31161, x32231);
  nand n32233(x32233, x31160, x32230);
  nand n32234(x32234, x32233, x32232);
  nand n32236(x32236, x32228, x32232);
  nand n32237(x32237, x31170, x31179);
  nand n32238(x32238, x31169, x31178);
  nand n32239(x32239, x32238, x32237);
  nand n32241(x32241, x84305, x32240);
  nand n32242(x32242, x29805, x32239);
  nand n32243(x32243, x32242, x32241);
  nand n32245(x32245, x32237, x32241);
  nand n32246(x32246, x31108, x31117);
  nand n32249(x32249, x32248, x32247);
  nand n32250(x32250, x32249, x32246);
  nand n32252(x32252, x31126, x32251);
  nand n32254(x32254, x32253, x32250);
  nand n32255(x32255, x32254, x32252);
  nand n32257(x32257, x32246, x32252);
  nand n32258(x32258, x31135, x31144);
  nand n32261(x32261, x32260, x32259);
  nand n32262(x32262, x32261, x32258);
  nand n32264(x32264, x31153, x32263);
  nand n32266(x32266, x32265, x32262);
  nand n32267(x32267, x32266, x32264);
  nand n32269(x32269, x32258, x32264);
  nand n32270(x32270, x31162, x31171);
  nand n32273(x32273, x32272, x32271);
  nand n32274(x32274, x32273, x32270);
  nand n32276(x32276, x31180, x32275);
  nand n32278(x32278, x32277, x32274);
  nand n32279(x32279, x32278, x32276);
  nand n32281(x32281, x32270, x32276);
  nand n32282(x32282, x31196, x31205);
  nand n32283(x32283, x31195, x31204);
  nand n32284(x32284, x32283, x32282);
  nand n32286(x32286, x31214, x32285);
  nand n32287(x32287, x31213, x32284);
  nand n32288(x32288, x32287, x32286);
  nand n32290(x32290, x32282, x32286);
  nand n32291(x32291, x31223, x31232);
  nand n32292(x32292, x31222, x31231);
  nand n32293(x32293, x32292, x32291);
  nand n32295(x32295, x31241, x32294);
  nand n32296(x32296, x31240, x32293);
  nand n32297(x32297, x32296, x32295);
  nand n32299(x32299, x32291, x32295);
  nand n32300(x32300, x31250, x31259);
  nand n32301(x32301, x31249, x31258);
  nand n32302(x32302, x32301, x32300);
  nand n32304(x32304, x84306, x32303);
  nand n32305(x32305, x31263, x32302);
  nand n32306(x32306, x32305, x32304);
  nand n32308(x32308, x32300, x32304);
  nand n32309(x32309, x31188, x31197);
  nand n32312(x32312, x32311, x32310);
  nand n32313(x32313, x32312, x32309);
  nand n32315(x32315, x31206, x32314);
  nand n32317(x32317, x32316, x32313);
  nand n32318(x32318, x32317, x32315);
  nand n32320(x32320, x32309, x32315);
  nand n32321(x32321, x31215, x31224);
  nand n32324(x32324, x32323, x32322);
  nand n32325(x32325, x32324, x32321);
  nand n32327(x32327, x31233, x32326);
  nand n32329(x32329, x32328, x32325);
  nand n32330(x32330, x32329, x32327);
  nand n32332(x32332, x32321, x32327);
  nand n32333(x32333, x31242, x31251);
  nand n32336(x32336, x32335, x32334);
  nand n32337(x32337, x32336, x32333);
  nand n32339(x32339, x31260, x32338);
  nand n32341(x32341, x32340, x32337);
  nand n32342(x32342, x32341, x32339);
  nand n32344(x32344, x32333, x32339);
  nand n32345(x32345, x31271, x84349);
  nand n32346(x32346, x31270, x31261);
  nand n32347(x32347, x32346, x32345);
  nand n32349(x32349, x31280, x31289);
  nand n32350(x32350, x31279, x31288);
  nand n32351(x32351, x32350, x32349);
  nand n32353(x32353, x31298, x32352);
  nand n32354(x32354, x31297, x32351);
  nand n32355(x32355, x32354, x32353);
  nand n32357(x32357, x32349, x32353);
  nand n32358(x32358, x31307, x31316);
  nand n32359(x32359, x31306, x31315);
  nand n32360(x32360, x32359, x32358);
  nand n32362(x32362, x31325, x32361);
  nand n32363(x32363, x31324, x32360);
  nand n32364(x32364, x32363, x32362);
  nand n32366(x32366, x32358, x32362);
  nand n32367(x32367, x31334, x31343);
  nand n32368(x32368, x31333, x31342);
  nand n32369(x32369, x32368, x32367);
  nand n32371(x32371, x31352, x32370);
  nand n32372(x32372, x31351, x32369);
  nand n32373(x32373, x32372, x32371);
  nand n32375(x32375, x32367, x32371);
  nand n32376(x32376, x31272, x31281);
  nand n32379(x32379, x32378, x32377);
  nand n32380(x32380, x32379, x32376);
  nand n32382(x32382, x31290, x32381);
  nand n32384(x32384, x32383, x32380);
  nand n32385(x32385, x32384, x32382);
  nand n32387(x32387, x32376, x32382);
  nand n32388(x32388, x31299, x31308);
  nand n32391(x32391, x32390, x32389);
  nand n32392(x32392, x32391, x32388);
  nand n32394(x32394, x31317, x32393);
  nand n32396(x32396, x32395, x32392);
  nand n32397(x32397, x32396, x32394);
  nand n32399(x32399, x32388, x32394);
  nand n32400(x32400, x31326, x31335);
  nand n32403(x32403, x32402, x32401);
  nand n32404(x32404, x32403, x32400);
  nand n32406(x32406, x31344, x32405);
  nand n32408(x32408, x32407, x32404);
  nand n32409(x32409, x32408, x32406);
  nand n32411(x32411, x32400, x32406);
  nand n32413(x32413, x31361, x31353);
  nand n32414(x32414, x31360, x32412);
  nand n32415(x32415, x32414, x32413);
  nand n32417(x32417, x31370, x31379);
  nand n32418(x32418, x31369, x31378);
  nand n32419(x32419, x32418, x32417);
  nand n32421(x32421, x31388, x32420);
  nand n32422(x32422, x31387, x32419);
  nand n32423(x32423, x32422, x32421);
  nand n32425(x32425, x32417, x32421);
  nand n32426(x32426, x31397, x31406);
  nand n32427(x32427, x31396, x31405);
  nand n32428(x32428, x32427, x32426);
  nand n32430(x32430, x31415, x32429);
  nand n32431(x32431, x31414, x32428);
  nand n32432(x32432, x32431, x32430);
  nand n32434(x32434, x32426, x32430);
  nand n32435(x32435, x31424, x31433);
  nand n32436(x32436, x31423, x31432);
  nand n32437(x32437, x32436, x32435);
  nand n32439(x32439, x31442, x32438);
  nand n32440(x32440, x31441, x32437);
  nand n32441(x32441, x32440, x32439);
  nand n32443(x32443, x32435, x32439);
  nand n32444(x32444, x31362, x31371);
  nand n32447(x32447, x32446, x32445);
  nand n32448(x32448, x32447, x32444);
  nand n32450(x32450, x31380, x32449);
  nand n32452(x32452, x32451, x32448);
  nand n32453(x32453, x32452, x32450);
  nand n32455(x32455, x31389, x31398);
  nand n32458(x32458, x32457, x32456);
  nand n32459(x32459, x32458, x32455);
  nand n32461(x32461, x31407, x32460);
  nand n32463(x32463, x32462, x32459);
  nand n32464(x32464, x32463, x32461);
  nand n32466(x32466, x31416, x31425);
  nand n32469(x32469, x32468, x32467);
  nand n32470(x32470, x32469, x32466);
  nand n32472(x32472, x31434, x32471);
  nand n32474(x32474, x32473, x32470);
  nand n32475(x32475, x32474, x32472);
  nand n32478(x32478, x31451, x31443);
  nand n32479(x32479, x31450, x32477);
  nand n32480(x32480, x32479, x32478);
  nand n32482(x32482, x31459, x31467);
  nand n32483(x32483, x31458, x31466);
  nand n32484(x32484, x32483, x32482);
  nand n32486(x32486, x31475, x32485);
  nand n32487(x32487, x31474, x32484);
  nand n32488(x32488, x32487, x32486);
  nand n32490(x32490, x31483, x31491);
  nand n32491(x32491, x31482, x31490);
  nand n32492(x32492, x32491, x32490);
  nand n32494(x32494, x31499, x32493);
  nand n32495(x32495, x31498, x32492);
  nand n32496(x32496, x32495, x32494);
  nand n32498(x32498, x31507, x31515);
  nand n32499(x32499, x31506, x31514);
  nand n32500(x32500, x32499, x32498);
  nand n32502(x32502, x31523, x32501);
  nand n32503(x32503, x31522, x32500);
  nand n32504(x32504, x32503, x32502);
  nand n32506(x32506, x84308, x84354);
  nand n32507(x32507, x29021, x30066);
  nand n32508(x32508, x32507, x32506);
  nand n32510(x32510, x84309, x84355);
  nand n32511(x32511, x30078, x30074);
  nand n32512(x32512, x32511, x32510);
  nand n32514(x32514, x84310, x84356);
  nand n32515(x32515, x30093, x30085);
  nand n32516(x32516, x32515, x32514);
  nand n32518(x32518, x84311, x84358);
  nand n32519(x32519, x31541, x30101);
  nand n32520(x32520, x32519, x32518);
  nand n32522(x32522, x84312, x84362);
  nand n32523(x32523, x31549, x30118);
  nand n32524(x32524, x32523, x32522);
  nand n32526(x32526, x84313, x84366);
  nand n32527(x32527, x31562, x30138);
  nand n32528(x32528, x32527, x32526);
  nand n32531(x32531, x31581, x84369);
  nand n32532(x32532, x31580, x30164);
  nand n32533(x32533, x32532, x32531);
  nand n32537(x32537, x31601, x84371);
  nand n32538(x32538, x31600, x30190);
  nand n32539(x32539, x32538, x32537);
  nand n32543(x32543, x84314, x84372);
  nand n32544(x32544, x30210, x31612);
  nand n32545(x32545, x32544, x32543);
  nand n32547(x32547, x31621, x84373);
  nand n32548(x32548, x31620, x30219);
  nand n32549(x32549, x32548, x32547);
  nand n32553(x32553, x30247, x84374);
  nand n32554(x32554, x31634, x31632);
  nand n32555(x32555, x32554, x32553);
  nand n32557(x32557, x31642, x84375);
  nand n32558(x32558, x31641, x30254);
  nand n32559(x32559, x32558, x32557);
  nand n32563(x32563, x30282, x84377);
  nand n32564(x32564, x31655, x31653);
  nand n32565(x32565, x32564, x32563);
  nand n32567(x32567, x31663, x84378);
  nand n32568(x32568, x31662, x30289);
  nand n32569(x32569, x32568, x32567);
  nand n32573(x32573, x84315, x84380);
  nand n32574(x32574, x31679, x31674);
  nand n32575(x32575, x32574, x32573);
  nand n32577(x32577, x31687, x84381);
  nand n32578(x32578, x31686, x30327);
  nand n32579(x32579, x32578, x32577);
  nand n32581(x32581, x31675, x84316);
  nand n32583(x32583, x32582, x31676);
  nand n32584(x32584, x32583, x32581);
  nand n32586(x32586, x84317, x84384);
  nand n32587(x32587, x31704, x31698);
  nand n32588(x32588, x32587, x32586);
  nand n32590(x32590, x31712, x84386);
  nand n32591(x32591, x31711, x30370);
  nand n32592(x32592, x32591, x32590);
  nand n32594(x32594, x31699, x84318);
  nand n32596(x32596, x32595, x31700);
  nand n32597(x32597, x32596, x32594);
  nand n32599(x32599, x84319, x31713);
  nand n32600(x32600, x31714, x32598);
  nand n32601(x32601, x32600, x32599);
  nand n32603(x32603, x84320, x84391);
  nand n32604(x32604, x31732, x31726);
  nand n32605(x32605, x32604, x32603);
  nand n32607(x32607, x31740, x84393);
  nand n32608(x32608, x31739, x30414);
  nand n32609(x32609, x32608, x32607);
  nand n32611(x32611, x31727, x84321);
  nand n32613(x32613, x32612, x31728);
  nand n32614(x32614, x32613, x32611);
  nand n32616(x32616, x84322, x31741);
  nand n32617(x32617, x31742, x32615);
  nand n32618(x32618, x32617, x32616);
  nand n32620(x32620, x31765, x84398);
  nand n32621(x32621, x31764, x31754);
  nand n32622(x32622, x32621, x32620);
  nand n32624(x32624, x31774, x84400);
  nand n32625(x32625, x31773, x30461);
  nand n32626(x32626, x32625, x32624);
  nand n32628(x32628, x31755, x31766);
  nand n32631(x32631, x32630, x32629);
  nand n32632(x32632, x32631, x32628);
  nand n32634(x32634, x84323, x31775);
  nand n32635(x32635, x31776, x32633);
  nand n32636(x32636, x32635, x32634);
  nand n32638(x32638, x31800, x84405);
  nand n32639(x32639, x31799, x31788);
  nand n32640(x32640, x32639, x32638);
  nand n32642(x32642, x31809, x84407);
  nand n32643(x32643, x31808, x30514);
  nand n32644(x32644, x32643, x32642);
  nand n32646(x32646, x31789, x31801);
  nand n32649(x32649, x32648, x32647);
  nand n32650(x32650, x32649, x32646);
  nand n32652(x32652, x31818, x31810);
  nand n32654(x32654, x32653, x32651);
  nand n32655(x32655, x32654, x32652);
  nand n32657(x32657, x31840, x84412);
  nand n32658(x32658, x31839, x31828);
  nand n32659(x32659, x32658, x32657);
  nand n32661(x32661, x31849, x84414);
  nand n32662(x32662, x31848, x30567);
  nand n32663(x32663, x32662, x32661);
  nand n32665(x32665, x31829, x31841);
  nand n32668(x32668, x32667, x32666);
  nand n32669(x32669, x32668, x32665);
  nand n32671(x32671, x31858, x31850);
  nand n32673(x32673, x32672, x32670);
  nand n32674(x32674, x32673, x32671);
  nand n32676(x32676, x31880, x84419);
  nand n32677(x32677, x31879, x31868);
  nand n32678(x32678, x32677, x32676);
  nand n32680(x32680, x84324, x84325);
  nand n32681(x32681, x30614, x30623);
  nand n32682(x32682, x32681, x32680);
  nand n32684(x32684, x31889, x32683);
  nand n32685(x32685, x31888, x32682);
  nand n32686(x32686, x32685, x32684);
  nand n32688(x32688, x32680, x32684);
  nand n32689(x32689, x31869, x31881);
  nand n32692(x32692, x32691, x32690);
  nand n32693(x32693, x32692, x32689);
  nand n32695(x32695, x31898, x31890);
  nand n32697(x32697, x32696, x32694);
  nand n32698(x32698, x32697, x32695);
  nand n32700(x32700, x31920, x84425);
  nand n32701(x32701, x31919, x31908);
  nand n32702(x32702, x32701, x32700);
  nand n32704(x32704, x30678, x84326);
  nand n32705(x32705, x31922, x30685);
  nand n32706(x32706, x32705, x32704);
  nand n32708(x32708, x31930, x32707);
  nand n32709(x32709, x31929, x32706);
  nand n32710(x32710, x32709, x32708);
  nand n32712(x32712, x32704, x32708);
  nand n32713(x32713, x31939, x84327);
  nand n32714(x32714, x31938, x29501);
  nand n32715(x32715, x32714, x32713);
  nand n32716(x32716, x31909, x31921);
  nand n32719(x32719, x32718, x32717);
  nand n32720(x32720, x32719, x32716);
  nand n32722(x32722, x31940, x31931);
  nand n32724(x32724, x32723, x32721);
  nand n32725(x32725, x32724, x32722);
  nand n32727(x32727, x31962, x84432);
  nand n32728(x32728, x31961, x31950);
  nand n32729(x32729, x32728, x32727);
  nand n32731(x32731, x30740, x84328);
  nand n32732(x32732, x31964, x30747);
  nand n32733(x32733, x32732, x32731);
  nand n32735(x32735, x31972, x32734);
  nand n32736(x32736, x31971, x32733);
  nand n32737(x32737, x32736, x32735);
  nand n32739(x32739, x32731, x32735);
  nand n32740(x32740, x31981, x84329);
  nand n32741(x32741, x31980, x30805);
  nand n32742(x32742, x32741, x32740);
  nand n32743(x32743, x31951, x31963);
  nand n32746(x32746, x32745, x32744);
  nand n32747(x32747, x32746, x32743);
  nand n32749(x32749, x31982, x31973);
  nand n32751(x32751, x32750, x32748);
  nand n32752(x32752, x32751, x32749);
  nand n32754(x32754, x32004, x84439);
  nand n32755(x32755, x32003, x31992);
  nand n32756(x32756, x32755, x32754);
  nand n32758(x32758, x84330, x84332);
  nand n32759(x32759, x32009, x30812);
  nand n32760(x32760, x32759, x32758);
  nand n32762(x32762, x32017, x32761);
  nand n32763(x32763, x32016, x32760);
  nand n32764(x32764, x32763, x32762);
  nand n32766(x32766, x32758, x32762);
  nand n32767(x32767, x32026, x84333);
  nand n32768(x32768, x32025, x30874);
  nand n32769(x32769, x32768, x32767);
  nand n32770(x32770, x31993, x32005);
  nand n32773(x32773, x32772, x32771);
  nand n32774(x32774, x32773, x32770);
  nand n32776(x32776, x84331, x32775);
  nand n32777(x32777, x32006, x32774);
  nand n32778(x32778, x32777, x32776);
  nand n32780(x32780, x32770, x32776);
  nand n32782(x32782, x32027, x32018);
  nand n32784(x32784, x32783, x32781);
  nand n32785(x32785, x32784, x32782);
  nand n32787(x32787, x32049, x84444);
  nand n32788(x32788, x32048, x32037);
  nand n32789(x32789, x32788, x32787);
  nand n32791(x32791, x84334, x84336);
  nand n32792(x32792, x32055, x30882);
  nand n32793(x32793, x32792, x32791);
  nand n32795(x32795, x32063, x32794);
  nand n32796(x32796, x32062, x32793);
  nand n32797(x32797, x32796, x32795);
  nand n32799(x32799, x32791, x32795);
  nand n32800(x32800, x32072, x84337);
  nand n32801(x32801, x32071, x32076);
  nand n32802(x32802, x32801, x32800);
  nand n32803(x32803, x32038, x32050);
  nand n32806(x32806, x32805, x32804);
  nand n32807(x32807, x32806, x32803);
  nand n32809(x32809, x84335, x32808);
  nand n32810(x32810, x32051, x32807);
  nand n32811(x32811, x32810, x32809);
  nand n32813(x32813, x32803, x32809);
  nand n32815(x32815, x32073, x32064);
  nand n32817(x32817, x32816, x32814);
  nand n32818(x32818, x32817, x32815);
  nand n32820(x32820, x84338, x32087);
  nand n32821(x32821, x32074, x32086);
  nand n32822(x32822, x32821, x32820);
  nand n32824(x32824, x32099, x32823);
  nand n32825(x32825, x32098, x32822);
  nand n32826(x32826, x32825, x32824);
  nand n32828(x32828, x32820, x32824);
  nand n32829(x32829, x84339, x84341);
  nand n32830(x32830, x32105, x30953);
  nand n32831(x32831, x32830, x32829);
  nand n32833(x32833, x32113, x32832);
  nand n32834(x32834, x32112, x32831);
  nand n32835(x32835, x32834, x32833);
  nand n32837(x32837, x32829, x32833);
  nand n32838(x32838, x32122, x84342);
  nand n32839(x32839, x32121, x32126);
  nand n32840(x32840, x32839, x32838);
  nand n32841(x32841, x32088, x32100);
  nand n32844(x32844, x32843, x32842);
  nand n32845(x32845, x32844, x32841);
  nand n32847(x32847, x84340, x32846);
  nand n32848(x32848, x32101, x32845);
  nand n32849(x32849, x32848, x32847);
  nand n32851(x32851, x32841, x32847);
  nand n32853(x32853, x32123, x32114);
  nand n32855(x32855, x32854, x32852);
  nand n32856(x32856, x32855, x32853);
  nand n32858(x32858, x84343, x32137);
  nand n32859(x32859, x32124, x32136);
  nand n32860(x32860, x32859, x32858);
  nand n32862(x32862, x32149, x32861);
  nand n32863(x32863, x32148, x32860);
  nand n32864(x32864, x32863, x32862);
  nand n32866(x32866, x32858, x32862);
  nand n32867(x32867, x32160, x84344);
  nand n32868(x32868, x32159, x31027);
  nand n32869(x32869, x32868, x32867);
  nand n32871(x32871, x32169, x32870);
  nand n32872(x32872, x32168, x32869);
  nand n32873(x32873, x32872, x32871);
  nand n32875(x32875, x32867, x32871);
  nand n32876(x32876, x32178, x84345);
  nand n32877(x32877, x32177, x32182);
  nand n32878(x32878, x32877, x32876);
  nand n32879(x32879, x32138, x32150);
  nand n32882(x32882, x32881, x32880);
  nand n32883(x32883, x32882, x32879);
  nand n32885(x32885, x32161, x32884);
  nand n32887(x32887, x32886, x32883);
  nand n32888(x32888, x32887, x32885);
  nand n32890(x32890, x32879, x32885);
  nand n32892(x32892, x32179, x32170);
  nand n32894(x32894, x32893, x32891);
  nand n32895(x32895, x32894, x32892);
  nand n32897(x32897, x84346, x32193);
  nand n32898(x32898, x32180, x32192);
  nand n32899(x32899, x32898, x32897);
  nand n32901(x32901, x32205, x32900);
  nand n32902(x32902, x32204, x32899);
  nand n32903(x32903, x32902, x32901);
  nand n32905(x32905, x32897, x32901);
  nand n32906(x32906, x32217, x84347);
  nand n32907(x32907, x32216, x31107);
  nand n32908(x32908, x32907, x32906);
  nand n32910(x32910, x32226, x32909);
  nand n32911(x32911, x32225, x32908);
  nand n32912(x32912, x32911, x32910);
  nand n32914(x32914, x32906, x32910);
  nand n32915(x32915, x32235, x32244);
  nand n32916(x32916, x32234, x32243);
  nand n32917(x32917, x32916, x32915);
  nand n32918(x32918, x32194, x32206);
  nand n32921(x32921, x32920, x32919);
  nand n32922(x32922, x32921, x32918);
  nand n32924(x32924, x32218, x32923);
  nand n32926(x32926, x32925, x32922);
  nand n32927(x32927, x32926, x32924);
  nand n32929(x32929, x32918, x32924);
  nand n32931(x32931, x32236, x32227);
  nand n32933(x32933, x32932, x32930);
  nand n32934(x32934, x32933, x32931);
  nand n32936(x32936, x32245, x32256);
  nand n32938(x32938, x32937, x32255);
  nand n32939(x32939, x32938, x32936);
  nand n32941(x32941, x32268, x32940);
  nand n32942(x32942, x32267, x32939);
  nand n32943(x32943, x32942, x32941);
  nand n32945(x32945, x32936, x32941);
  nand n32946(x32946, x32280, x84348);
  nand n32947(x32947, x32279, x31187);
  nand n32948(x32948, x32947, x32946);
  nand n32950(x32950, x32289, x32949);
  nand n32951(x32951, x32288, x32948);
  nand n32952(x32952, x32951, x32950);
  nand n32954(x32954, x32946, x32950);
  nand n32955(x32955, x32298, x32307);
  nand n32956(x32956, x32297, x32306);
  nand n32957(x32957, x32956, x32955);
  nand n32958(x32958, x32257, x32269);
  nand n32961(x32961, x32960, x32959);
  nand n32962(x32962, x32961, x32958);
  nand n32964(x32964, x32281, x32963);
  nand n32966(x32966, x32965, x32962);
  nand n32967(x32967, x32966, x32964);
  nand n32969(x32969, x32958, x32964);
  nand n32971(x32971, x32299, x32290);
  nand n32973(x32973, x32972, x32970);
  nand n32974(x32974, x32973, x32971);
  nand n32976(x32976, x32308, x32319);
  nand n32978(x32978, x32977, x32318);
  nand n32979(x32979, x32978, x32976);
  nand n32981(x32981, x32331, x32980);
  nand n32982(x32982, x32330, x32979);
  nand n32983(x32983, x32982, x32981);
  nand n32985(x32985, x32976, x32981);
  nand n32986(x32986, x32343, x32348);
  nand n32987(x32987, x32342, x32347);
  nand n32988(x32988, x32987, x32986);
  nand n32990(x32990, x32356, x32989);
  nand n32991(x32991, x32355, x32988);
  nand n32992(x32992, x32991, x32990);
  nand n32994(x32994, x32986, x32990);
  nand n32995(x32995, x32365, x32374);
  nand n32996(x32996, x32364, x32373);
  nand n32997(x32997, x32996, x32995);
  nand n32998(x32998, x32320, x32332);
  nand n33001(x33001, x33000, x32999);
  nand n33002(x33002, x33001, x32998);
  nand n33004(x33004, x32344, x33003);
  nand n33006(x33006, x33005, x33002);
  nand n33007(x33007, x33006, x33004);
  nand n33009(x33009, x32998, x33004);
  nand n33010(x33010, x84350, x32357);
  nand n33012(x33012, x32345, x33011);
  nand n33013(x33013, x33012, x33010);
  nand n33015(x33015, x32366, x33014);
  nand n33017(x33017, x33016, x33013);
  nand n33018(x33018, x33017, x33015);
  nand n33020(x33020, x33010, x33015);
  nand n33021(x33021, x32375, x32386);
  nand n33023(x33023, x33022, x32385);
  nand n33024(x33024, x33023, x33021);
  nand n33026(x33026, x32398, x33025);
  nand n33027(x33027, x32397, x33024);
  nand n33028(x33028, x33027, x33026);
  nand n33030(x33030, x33021, x33026);
  nand n33031(x33031, x32410, x32416);
  nand n33032(x33032, x32409, x32415);
  nand n33033(x33033, x33032, x33031);
  nand n33035(x33035, x32424, x33034);
  nand n33036(x33036, x32423, x33033);
  nand n33037(x33037, x33036, x33035);
  nand n33039(x33039, x33031, x33035);
  nand n33040(x33040, x32433, x32442);
  nand n33041(x33041, x32432, x32441);
  nand n33042(x33042, x33041, x33040);
  nand n33044(x33044, x84307, x33043);
  nand n33045(x33045, x29984, x33042);
  nand n33046(x33046, x33045, x33044);
  nand n33048(x33048, x33040, x33044);
  nand n33049(x33049, x32387, x32399);
  nand n33052(x33052, x33051, x33050);
  nand n33053(x33053, x33052, x33049);
  nand n33055(x33055, x32411, x33054);
  nand n33057(x33057, x33056, x33053);
  nand n33058(x33058, x33057, x33055);
  nand n33060(x33060, x84351, x32425);
  nand n33062(x33062, x32413, x33061);
  nand n33063(x33063, x33062, x33060);
  nand n33065(x33065, x32434, x33064);
  nand n33067(x33067, x33066, x33063);
  nand n33068(x33068, x33067, x33065);
  nand n33070(x33070, x32443, x32454);
  nand n33072(x33072, x33071, x32453);
  nand n33073(x33073, x33072, x33070);
  nand n33075(x33075, x32465, x33074);
  nand n33076(x33076, x32464, x33073);
  nand n33077(x33077, x33076, x33075);
  nand n33079(x33079, x32476, x32481);
  nand n33080(x33080, x32475, x32480);
  nand n33081(x33081, x33080, x33079);
  nand n33083(x33083, x32489, x33082);
  nand n33084(x33084, x32488, x33081);
  nand n33085(x33085, x33084, x33083);
  nand n33087(x33087, x32497, x32505);
  nand n33088(x33088, x32496, x32504);
  nand n33089(x33089, x33088, x33087);
  nand n33091(x33091, x31527, x33090);
  nand n33092(x33092, x31526, x33089);
  nand n33093(x33093, x33092, x33091);
  nand n33095(x33095, x84352, x84353);
  nand n33096(x33096, x30049, x30058);
  nand n33097(x33097, x33096, x33095);
  nand n33098(x33098, x32509, x30059);
  nand n33099(x33099, x32508, x31528);
  nand n33100(x33100, x33099, x33098);
  nand n33101(x33101, x32513, x30067);
  nand n33102(x33102, x32512, x31529);
  nand n33103(x33103, x33102, x33101);
  nand n33105(x33105, x32517, x84463);
  nand n33106(x33106, x32516, x31533);
  nand n33107(x33107, x33106, x33105);
  nand n33109(x33109, x84357, x84464);
  nand n33110(x33110, x31530, x32514);
  nand n33111(x33111, x33110, x33109);
  nand n33112(x33112, x32521, x84465);
  nand n33113(x33113, x32520, x31538);
  nand n33114(x33114, x33113, x33112);
  nand n33116(x33116, x84359, x84467);
  nand n33117(x33117, x31534, x32518);
  nand n33118(x33118, x33117, x33116);
  nand n33119(x33119, x84360, x84361);
  nand n33120(x33120, x31539, x31546);
  nand n33121(x33121, x33120, x33119);
  nand n33123(x33123, x32525, x33122);
  nand n33124(x33124, x32524, x33121);
  nand n33125(x33125, x33124, x33123);
  nand n33127(x33127, x33119, x33123);
  nand n33128(x33128, x84363, x84468);
  nand n33129(x33129, x31542, x32522);
  nand n33130(x33130, x33129, x33128);
  nand n33131(x33131, x84364, x84365);
  nand n33132(x33132, x31547, x31558);
  nand n33133(x33133, x33132, x33131);
  nand n33135(x33135, x32529, x33134);
  nand n33136(x33136, x32528, x33133);
  nand n33137(x33137, x33136, x33135);
  nand n33139(x33139, x33131, x33135);
  nand n33140(x33140, x31559, x84469);
  nand n33141(x33141, x32530, x32526);
  nand n33142(x33142, x33141, x33140);
  nand n33143(x33143, x84367, x84368);
  nand n33144(x33144, x31560, x31572);
  nand n33145(x33145, x33144, x33143);
  nand n33147(x33147, x32534, x33146);
  nand n33148(x33148, x32533, x33145);
  nand n33149(x33149, x33148, x33147);
  nand n33151(x33151, x33143, x33147);
  nand n33152(x33152, x31573, x84470);
  nand n33153(x33153, x32535, x32531);
  nand n33154(x33154, x33153, x33152);
  nand n33155(x33155, x31582, x84370);
  nand n33156(x33156, x32536, x31592);
  nand n33157(x33157, x33156, x33155);
  nand n33159(x33159, x32540, x33158);
  nand n33160(x33160, x32539, x33157);
  nand n33161(x33161, x33160, x33159);
  nand n33163(x33163, x33155, x33159);
  nand n33164(x33164, x31593, x84471);
  nand n33165(x33165, x32541, x32537);
  nand n33166(x33166, x33165, x33164);
  nand n33167(x33167, x31602, x32546);
  nand n33168(x33168, x32542, x32545);
  nand n33169(x33169, x33168, x33167);
  nand n33171(x33171, x32550, x33170);
  nand n33172(x33172, x32549, x33169);
  nand n33173(x33173, x33172, x33171);
  nand n33175(x33175, x33167, x33171);
  nand n33176(x33176, x31613, x84473);
  nand n33177(x33177, x32551, x32547);
  nand n33178(x33178, x33177, x33176);
  nand n33180(x33180, x31622, x32556);
  nand n33181(x33181, x32552, x32555);
  nand n33182(x33182, x33181, x33180);
  nand n33184(x33184, x32560, x33183);
  nand n33185(x33185, x32559, x33182);
  nand n33186(x33186, x33185, x33184);
  nand n33188(x33188, x33180, x33184);
  nand n33189(x33189, x31633, x84475);
  nand n33190(x33190, x32561, x32557);
  nand n33191(x33191, x33190, x33189);
  nand n33193(x33193, x31643, x32566);
  nand n33194(x33194, x32562, x32565);
  nand n33195(x33195, x33194, x33193);
  nand n33197(x33197, x32570, x33196);
  nand n33198(x33198, x32569, x33195);
  nand n33199(x33199, x33198, x33197);
  nand n33201(x33201, x33193, x33197);
  nand n33202(x33202, x31654, x84477);
  nand n33203(x33203, x32571, x32567);
  nand n33204(x33204, x33203, x33202);
  nand n33206(x33206, x31664, x32576);
  nand n33207(x33207, x32572, x32575);
  nand n33208(x33208, x33207, x33206);
  nand n33210(x33210, x32580, x33209);
  nand n33211(x33211, x32579, x33208);
  nand n33212(x33212, x33211, x33210);
  nand n33214(x33214, x33206, x33210);
  nand n33215(x33215, x84383, x84479);
  nand n33216(x33216, x32584, x32577);
  nand n33217(x33217, x33216, x33215);
  nand n33219(x33219, x31688, x32589);
  nand n33220(x33220, x32585, x32588);
  nand n33221(x33221, x33220, x33219);
  nand n33223(x33223, x32593, x33222);
  nand n33224(x33224, x32592, x33221);
  nand n33225(x33225, x33224, x33223);
  nand n33227(x33227, x33219, x33223);
  nand n33228(x33228, x84385, x84480);
  nand n33229(x33229, x32586, x32581);
  nand n33230(x33230, x33229, x33228);
  nand n33232(x33232, x84388, x84482);
  nand n33233(x33233, x32597, x32590);
  nand n33234(x33234, x33233, x33232);
  nand n33236(x33236, x32602, x32606);
  nand n33237(x33237, x32601, x32605);
  nand n33238(x33238, x33237, x33236);
  nand n33240(x33240, x32610, x33239);
  nand n33241(x33241, x32609, x33238);
  nand n33242(x33242, x33241, x33240);
  nand n33244(x33244, x33236, x33240);
  nand n33245(x33245, x84389, x84390);
  nand n33246(x33246, x32594, x32599);
  nand n33247(x33247, x33246, x33245);
  nand n33249(x33249, x84392, x33248);
  nand n33250(x33250, x32603, x33247);
  nand n33251(x33251, x33250, x33249);
  nand n33253(x33253, x33245, x33249);
  nand n33254(x33254, x84395, x84484);
  nand n33255(x33255, x32614, x32607);
  nand n33256(x33256, x33255, x33254);
  nand n33258(x33258, x32619, x32623);
  nand n33259(x33259, x32618, x32622);
  nand n33260(x33260, x33259, x33258);
  nand n33262(x33262, x32627, x33261);
  nand n33263(x33263, x32626, x33260);
  nand n33264(x33264, x33263, x33262);
  nand n33266(x33266, x33258, x33262);
  nand n33267(x33267, x84396, x84397);
  nand n33268(x33268, x32611, x32616);
  nand n33269(x33269, x33268, x33267);
  nand n33271(x33271, x84399, x33270);
  nand n33272(x33272, x32620, x33269);
  nand n33273(x33273, x33272, x33271);
  nand n33275(x33275, x33267, x33271);
  nand n33276(x33276, x84402, x84486);
  nand n33277(x33277, x32632, x32624);
  nand n33278(x33278, x33277, x33276);
  nand n33280(x33280, x32637, x32641);
  nand n33281(x33281, x32636, x32640);
  nand n33282(x33282, x33281, x33280);
  nand n33284(x33284, x32645, x33283);
  nand n33285(x33285, x32644, x33282);
  nand n33286(x33286, x33285, x33284);
  nand n33288(x33288, x33280, x33284);
  nand n33289(x33289, x84403, x84404);
  nand n33290(x33290, x32628, x32634);
  nand n33291(x33291, x33290, x33289);
  nand n33293(x33293, x84406, x33292);
  nand n33294(x33294, x32638, x33291);
  nand n33295(x33295, x33294, x33293);
  nand n33297(x33297, x33289, x33293);
  nand n33298(x33298, x84409, x84488);
  nand n33299(x33299, x32650, x32642);
  nand n33300(x33300, x33299, x33298);
  nand n33302(x33302, x32656, x32660);
  nand n33303(x33303, x32655, x32659);
  nand n33304(x33304, x33303, x33302);
  nand n33306(x33306, x32664, x33305);
  nand n33307(x33307, x32663, x33304);
  nand n33308(x33308, x33307, x33306);
  nand n33310(x33310, x33302, x33306);
  nand n33311(x33311, x84410, x84411);
  nand n33312(x33312, x32646, x32652);
  nand n33313(x33313, x33312, x33311);
  nand n33315(x33315, x84413, x33314);
  nand n33316(x33316, x32657, x33313);
  nand n33317(x33317, x33316, x33315);
  nand n33319(x33319, x33311, x33315);
  nand n33320(x33320, x84416, x84490);
  nand n33321(x33321, x32669, x32661);
  nand n33322(x33322, x33321, x33320);
  nand n33324(x33324, x32675, x32679);
  nand n33325(x33325, x32674, x32678);
  nand n33326(x33326, x33325, x33324);
  nand n33328(x33328, x32687, x33327);
  nand n33329(x33329, x32686, x33326);
  nand n33330(x33330, x33329, x33328);
  nand n33332(x33332, x33324, x33328);
  nand n33333(x33333, x84417, x84418);
  nand n33334(x33334, x32665, x32671);
  nand n33335(x33335, x33334, x33333);
  nand n33337(x33337, x84420, x33336);
  nand n33338(x33338, x32676, x33335);
  nand n33339(x33339, x33338, x33337);
  nand n33341(x33341, x33333, x33337);
  nand n33343(x33343, x84422, x32688);
  nand n33344(x33344, x32693, x33342);
  nand n33345(x33345, x33344, x33343);
  nand n33347(x33347, x32699, x32703);
  nand n33348(x33348, x32698, x32702);
  nand n33349(x33349, x33348, x33347);
  nand n33351(x33351, x32711, x33350);
  nand n33352(x33352, x32710, x33349);
  nand n33353(x33353, x33352, x33351);
  nand n33355(x33355, x33347, x33351);
  nand n33356(x33356, x84423, x84424);
  nand n33357(x33357, x32689, x32695);
  nand n33358(x33358, x33357, x33356);
  nand n33360(x33360, x84426, x33359);
  nand n33361(x33361, x32700, x33358);
  nand n33362(x33362, x33361, x33360);
  nand n33364(x33364, x33356, x33360);
  nand n33365(x33365, x32712, x84428);
  nand n33367(x33367, x33366, x32713);
  nand n33368(x33368, x33367, x33365);
  nand n33370(x33370, x84429, x33369);
  nand n33371(x33371, x32720, x33368);
  nand n33372(x33372, x33371, x33370);
  nand n33374(x33374, x33365, x33370);
  nand n33375(x33375, x32726, x32730);
  nand n33376(x33376, x32725, x32729);
  nand n33377(x33377, x33376, x33375);
  nand n33379(x33379, x32738, x33378);
  nand n33380(x33380, x32737, x33377);
  nand n33381(x33381, x33380, x33379);
  nand n33383(x33383, x33375, x33379);
  nand n33384(x33384, x84430, x84431);
  nand n33385(x33385, x32716, x32722);
  nand n33386(x33386, x33385, x33384);
  nand n33388(x33388, x84433, x33387);
  nand n33389(x33389, x32727, x33386);
  nand n33390(x33390, x33389, x33388);
  nand n33392(x33392, x33384, x33388);
  nand n33393(x33393, x32739, x84435);
  nand n33395(x33395, x33394, x32740);
  nand n33396(x33396, x33395, x33393);
  nand n33398(x33398, x84436, x33397);
  nand n33399(x33399, x32747, x33396);
  nand n33400(x33400, x33399, x33398);
  nand n33402(x33402, x33393, x33398);
  nand n33403(x33403, x32753, x32757);
  nand n33404(x33404, x32752, x32756);
  nand n33405(x33405, x33404, x33403);
  nand n33407(x33407, x32765, x33406);
  nand n33408(x33408, x32764, x33405);
  nand n33409(x33409, x33408, x33407);
  nand n33411(x33411, x33403, x33407);
  nand n33412(x33412, x84437, x84438);
  nand n33413(x33413, x32743, x32749);
  nand n33414(x33414, x33413, x33412);
  nand n33416(x33416, x84440, x33415);
  nand n33417(x33417, x32754, x33414);
  nand n33418(x33418, x33417, x33416);
  nand n33420(x33420, x33412, x33416);
  nand n33421(x33421, x32766, x84442);
  nand n33423(x33423, x33422, x32767);
  nand n33424(x33424, x33423, x33421);
  nand n33426(x33426, x32779, x33425);
  nand n33427(x33427, x32778, x33424);
  nand n33428(x33428, x33427, x33426);
  nand n33430(x33430, x33421, x33426);
  nand n33431(x33431, x32786, x32790);
  nand n33432(x33432, x32785, x32789);
  nand n33433(x33433, x33432, x33431);
  nand n33435(x33435, x32798, x33434);
  nand n33436(x33436, x32797, x33433);
  nand n33437(x33437, x33436, x33435);
  nand n33439(x33439, x33431, x33435);
  nand n33440(x33440, x32780, x84443);
  nand n33442(x33442, x33441, x32782);
  nand n33443(x33443, x33442, x33440);
  nand n33445(x33445, x84445, x33444);
  nand n33446(x33446, x32787, x33443);
  nand n33447(x33447, x33446, x33445);
  nand n33449(x33449, x33440, x33445);
  nand n33450(x33450, x32799, x84447);
  nand n33452(x33452, x33451, x32800);
  nand n33453(x33453, x33452, x33450);
  nand n33455(x33455, x32812, x33454);
  nand n33456(x33456, x32811, x33453);
  nand n33457(x33457, x33456, x33455);
  nand n33459(x33459, x33450, x33455);
  nand n33460(x33460, x32819, x32827);
  nand n33461(x33461, x32818, x32826);
  nand n33462(x33462, x33461, x33460);
  nand n33464(x33464, x32836, x33463);
  nand n33465(x33465, x32835, x33462);
  nand n33466(x33466, x33465, x33464);
  nand n33468(x33468, x33460, x33464);
  nand n33469(x33469, x32813, x84448);
  nand n33471(x33471, x33470, x32815);
  nand n33472(x33472, x33471, x33469);
  nand n33474(x33474, x32828, x33473);
  nand n33476(x33476, x33475, x33472);
  nand n33477(x33477, x33476, x33474);
  nand n33479(x33479, x33469, x33474);
  nand n33480(x33480, x32837, x84450);
  nand n33482(x33482, x33481, x32838);
  nand n33483(x33483, x33482, x33480);
  nand n33485(x33485, x32850, x33484);
  nand n33486(x33486, x32849, x33483);
  nand n33487(x33487, x33486, x33485);
  nand n33489(x33489, x33480, x33485);
  nand n33490(x33490, x32857, x32865);
  nand n33491(x33491, x32856, x32864);
  nand n33492(x33492, x33491, x33490);
  nand n33494(x33494, x32874, x33493);
  nand n33495(x33495, x32873, x33492);
  nand n33496(x33496, x33495, x33494);
  nand n33498(x33498, x33490, x33494);
  nand n33499(x33499, x32851, x84451);
  nand n33501(x33501, x33500, x32853);
  nand n33502(x33502, x33501, x33499);
  nand n33504(x33504, x32866, x33503);
  nand n33506(x33506, x33505, x33502);
  nand n33507(x33507, x33506, x33504);
  nand n33509(x33509, x33499, x33504);
  nand n33510(x33510, x32875, x84453);
  nand n33512(x33512, x33511, x32876);
  nand n33513(x33513, x33512, x33510);
  nand n33515(x33515, x32889, x33514);
  nand n33516(x33516, x32888, x33513);
  nand n33517(x33517, x33516, x33515);
  nand n33519(x33519, x33510, x33515);
  nand n33520(x33520, x32896, x32904);
  nand n33521(x33521, x32895, x32903);
  nand n33522(x33522, x33521, x33520);
  nand n33524(x33524, x32913, x33523);
  nand n33525(x33525, x32912, x33522);
  nand n33526(x33526, x33525, x33524);
  nand n33528(x33528, x33520, x33524);
  nand n33529(x33529, x32890, x84454);
  nand n33531(x33531, x33530, x32892);
  nand n33532(x33532, x33531, x33529);
  nand n33534(x33534, x32905, x33533);
  nand n33536(x33536, x33535, x33532);
  nand n33537(x33537, x33536, x33534);
  nand n33539(x33539, x33529, x33534);
  nand n33540(x33540, x32914, x84456);
  nand n33542(x33542, x33541, x32915);
  nand n33543(x33543, x33542, x33540);
  nand n33545(x33545, x32928, x33544);
  nand n33546(x33546, x32927, x33543);
  nand n33547(x33547, x33546, x33545);
  nand n33549(x33549, x33540, x33545);
  nand n33550(x33550, x32935, x32944);
  nand n33551(x33551, x32934, x32943);
  nand n33552(x33552, x33551, x33550);
  nand n33554(x33554, x32953, x33553);
  nand n33555(x33555, x32952, x33552);
  nand n33556(x33556, x33555, x33554);
  nand n33558(x33558, x33550, x33554);
  nand n33559(x33559, x32929, x84457);
  nand n33561(x33561, x33560, x32931);
  nand n33562(x33562, x33561, x33559);
  nand n33564(x33564, x32945, x33563);
  nand n33566(x33566, x33565, x33562);
  nand n33567(x33567, x33566, x33564);
  nand n33569(x33569, x33559, x33564);
  nand n33570(x33570, x32954, x84459);
  nand n33572(x33572, x33571, x32955);
  nand n33573(x33573, x33572, x33570);
  nand n33575(x33575, x32968, x33574);
  nand n33576(x33576, x32967, x33573);
  nand n33577(x33577, x33576, x33575);
  nand n33579(x33579, x33570, x33575);
  nand n33580(x33580, x32975, x32984);
  nand n33581(x33581, x32974, x32983);
  nand n33582(x33582, x33581, x33580);
  nand n33584(x33584, x32993, x33583);
  nand n33585(x33585, x32992, x33582);
  nand n33586(x33586, x33585, x33584);
  nand n33588(x33588, x33580, x33584);
  nand n33589(x33589, x32969, x84460);
  nand n33591(x33591, x33590, x32971);
  nand n33592(x33592, x33591, x33589);
  nand n33594(x33594, x32985, x33593);
  nand n33596(x33596, x33595, x33592);
  nand n33597(x33597, x33596, x33594);
  nand n33599(x33599, x33589, x33594);
  nand n33600(x33600, x32994, x84462);
  nand n33602(x33602, x33601, x32995);
  nand n33603(x33603, x33602, x33600);
  nand n33605(x33605, x33008, x33604);
  nand n33606(x33606, x33007, x33603);
  nand n33607(x33607, x33606, x33605);
  nand n33609(x33609, x33600, x33605);
  nand n33610(x33610, x33019, x33029);
  nand n33611(x33611, x33018, x33028);
  nand n33612(x33612, x33611, x33610);
  nand n33614(x33614, x33038, x33613);
  nand n33615(x33615, x33037, x33612);
  nand n33616(x33616, x33615, x33614);
  nand n33618(x33618, x33610, x33614);
  nand n33619(x33619, x33009, x33020);
  nand n33622(x33622, x33621, x33620);
  nand n33623(x33623, x33622, x33619);
  nand n33625(x33625, x33030, x33624);
  nand n33627(x33627, x33626, x33623);
  nand n33628(x33628, x33627, x33625);
  nand n33630(x33630, x33039, x33048);
  nand n33633(x33633, x33632, x33631);
  nand n33634(x33634, x33633, x33630);
  nand n33636(x33636, x33059, x33635);
  nand n33637(x33637, x33058, x33634);
  nand n33638(x33638, x33637, x33636);
  nand n33640(x33640, x33069, x33078);
  nand n33641(x33641, x33068, x33077);
  nand n33642(x33642, x33641, x33640);
  nand n33644(x33644, x33086, x33643);
  nand n33645(x33645, x33085, x33642);
  nand n33646(x33646, x33645, x33644);
  nand n33648(x33648, x33104, x84493);
  nand n33649(x33649, x33103, x32506);
  nand n33650(x33650, x33649, x33648);
  nand n33651(x33651, x33108, x84495);
  nand n33652(x33652, x33107, x32510);
  nand n33653(x33653, x33652, x33651);
  nand n33654(x33654, x33115, x84497);
  nand n33655(x33655, x33114, x33111);
  nand n33656(x33656, x33655, x33654);
  nand n33657(x33657, x84466, x84498);
  nand n33658(x33658, x33112, x33109);
  nand n33659(x33659, x33658, x33657);
  nand n33661(x33661, x33126, x84500);
  nand n33662(x33662, x33125, x33118);
  nand n33663(x33663, x33662, x33661);
  nand n33664(x33664, x33127, x84502);
  nand n33666(x33666, x33665, x33116);
  nand n33667(x33667, x33666, x33664);
  nand n33669(x33669, x33138, x84504);
  nand n33670(x33670, x33137, x33130);
  nand n33671(x33671, x33670, x33669);
  nand n33672(x33672, x33139, x84506);
  nand n33674(x33674, x33673, x33128);
  nand n33675(x33675, x33674, x33672);
  nand n33677(x33677, x33150, x84508);
  nand n33678(x33678, x33149, x33142);
  nand n33679(x33679, x33678, x33677);
  nand n33680(x33680, x33151, x84510);
  nand n33682(x33682, x33681, x33140);
  nand n33683(x33683, x33682, x33680);
  nand n33685(x33685, x33162, x84512);
  nand n33686(x33686, x33161, x33154);
  nand n33687(x33687, x33686, x33685);
  nand n33688(x33688, x33163, x84514);
  nand n33690(x33690, x33689, x33152);
  nand n33691(x33691, x33690, x33688);
  nand n33693(x33693, x33174, x84516);
  nand n33694(x33694, x33173, x33166);
  nand n33695(x33695, x33694, x33693);
  nand n33696(x33696, x33175, x84518);
  nand n33698(x33698, x33697, x33164);
  nand n33699(x33699, x33698, x33696);
  nand n33701(x33701, x84472, x33179);
  nand n33702(x33702, x32543, x33178);
  nand n33703(x33703, x33702, x33701);
  nand n33705(x33705, x33187, x33704);
  nand n33706(x33706, x33186, x33703);
  nand n33707(x33707, x33706, x33705);
  nand n33709(x33709, x33701, x33705);
  nand n33710(x33710, x33188, x84520);
  nand n33712(x33712, x33711, x33176);
  nand n33713(x33713, x33712, x33710);
  nand n33715(x33715, x84474, x33192);
  nand n33716(x33716, x32553, x33191);
  nand n33717(x33717, x33716, x33715);
  nand n33719(x33719, x33200, x33718);
  nand n33720(x33720, x33199, x33717);
  nand n33721(x33721, x33720, x33719);
  nand n33723(x33723, x33715, x33719);
  nand n33724(x33724, x33201, x84522);
  nand n33726(x33726, x33725, x33189);
  nand n33727(x33727, x33726, x33724);
  nand n33729(x33729, x84476, x33205);
  nand n33730(x33730, x32563, x33204);
  nand n33731(x33731, x33730, x33729);
  nand n33733(x33733, x33213, x33732);
  nand n33734(x33734, x33212, x33731);
  nand n33735(x33735, x33734, x33733);
  nand n33737(x33737, x33729, x33733);
  nand n33738(x33738, x33214, x84524);
  nand n33740(x33740, x33739, x33202);
  nand n33741(x33741, x33740, x33738);
  nand n33743(x33743, x84478, x33218);
  nand n33744(x33744, x32573, x33217);
  nand n33745(x33745, x33744, x33743);
  nand n33747(x33747, x33226, x33746);
  nand n33748(x33748, x33225, x33745);
  nand n33749(x33749, x33748, x33747);
  nand n33751(x33751, x33743, x33747);
  nand n33752(x33752, x33227, x84526);
  nand n33754(x33754, x33753, x33215);
  nand n33755(x33755, x33754, x33752);
  nand n33757(x33757, x33231, x33235);
  nand n33758(x33758, x33230, x33234);
  nand n33759(x33759, x33758, x33757);
  nand n33761(x33761, x33243, x33760);
  nand n33762(x33762, x33242, x33759);
  nand n33763(x33763, x33762, x33761);
  nand n33765(x33765, x33757, x33761);
  nand n33766(x33766, x84481, x84483);
  nand n33767(x33767, x33228, x33232);
  nand n33768(x33768, x33767, x33766);
  nand n33770(x33770, x33244, x33769);
  nand n33772(x33772, x33771, x33768);
  nand n33773(x33773, x33772, x33770);
  nand n33775(x33775, x33766, x33770);
  nand n33776(x33776, x33252, x33257);
  nand n33777(x33777, x33251, x33256);
  nand n33778(x33778, x33777, x33776);
  nand n33780(x33780, x33265, x33779);
  nand n33781(x33781, x33264, x33778);
  nand n33782(x33782, x33781, x33780);
  nand n33784(x33784, x33776, x33780);
  nand n33785(x33785, x33253, x84485);
  nand n33787(x33787, x33786, x33254);
  nand n33788(x33788, x33787, x33785);
  nand n33790(x33790, x33266, x33789);
  nand n33792(x33792, x33791, x33788);
  nand n33793(x33793, x33792, x33790);
  nand n33795(x33795, x33785, x33790);
  nand n33796(x33796, x33274, x33279);
  nand n33797(x33797, x33273, x33278);
  nand n33798(x33798, x33797, x33796);
  nand n33800(x33800, x33287, x33799);
  nand n33801(x33801, x33286, x33798);
  nand n33802(x33802, x33801, x33800);
  nand n33804(x33804, x33796, x33800);
  nand n33805(x33805, x33275, x84487);
  nand n33807(x33807, x33806, x33276);
  nand n33808(x33808, x33807, x33805);
  nand n33810(x33810, x33288, x33809);
  nand n33812(x33812, x33811, x33808);
  nand n33813(x33813, x33812, x33810);
  nand n33815(x33815, x33805, x33810);
  nand n33816(x33816, x33296, x33301);
  nand n33817(x33817, x33295, x33300);
  nand n33818(x33818, x33817, x33816);
  nand n33820(x33820, x33309, x33819);
  nand n33821(x33821, x33308, x33818);
  nand n33822(x33822, x33821, x33820);
  nand n33824(x33824, x33816, x33820);
  nand n33825(x33825, x33297, x84489);
  nand n33827(x33827, x33826, x33298);
  nand n33828(x33828, x33827, x33825);
  nand n33830(x33830, x33310, x33829);
  nand n33832(x33832, x33831, x33828);
  nand n33833(x33833, x33832, x33830);
  nand n33835(x33835, x33825, x33830);
  nand n33836(x33836, x33318, x33323);
  nand n33837(x33837, x33317, x33322);
  nand n33838(x33838, x33837, x33836);
  nand n33840(x33840, x33331, x33839);
  nand n33841(x33841, x33330, x33838);
  nand n33842(x33842, x33841, x33840);
  nand n33844(x33844, x33836, x33840);
  nand n33845(x33845, x33319, x84491);
  nand n33847(x33847, x33846, x33320);
  nand n33848(x33848, x33847, x33845);
  nand n33850(x33850, x33332, x33849);
  nand n33852(x33852, x33851, x33848);
  nand n33853(x33853, x33852, x33850);
  nand n33855(x33855, x33845, x33850);
  nand n33856(x33856, x33340, x33346);
  nand n33857(x33857, x33339, x33345);
  nand n33858(x33858, x33857, x33856);
  nand n33860(x33860, x33354, x33859);
  nand n33861(x33861, x33353, x33858);
  nand n33862(x33862, x33861, x33860);
  nand n33864(x33864, x33856, x33860);
  nand n33865(x33865, x33341, x84492);
  nand n33867(x33867, x33866, x33343);
  nand n33868(x33868, x33867, x33865);
  nand n33870(x33870, x33355, x33869);
  nand n33872(x33872, x33871, x33868);
  nand n33873(x33873, x33872, x33870);
  nand n33875(x33875, x33865, x33870);
  nand n33876(x33876, x33363, x33373);
  nand n33877(x33877, x33362, x33372);
  nand n33878(x33878, x33877, x33876);
  nand n33880(x33880, x33382, x33879);
  nand n33881(x33881, x33381, x33878);
  nand n33882(x33882, x33881, x33880);
  nand n33884(x33884, x33876, x33880);
  nand n33885(x33885, x33364, x33374);
  nand n33888(x33888, x33887, x33886);
  nand n33889(x33889, x33888, x33885);
  nand n33891(x33891, x33383, x33890);
  nand n33893(x33893, x33892, x33889);
  nand n33894(x33894, x33893, x33891);
  nand n33896(x33896, x33885, x33891);
  nand n33897(x33897, x33391, x33401);
  nand n33898(x33898, x33390, x33400);
  nand n33899(x33899, x33898, x33897);
  nand n33901(x33901, x33410, x33900);
  nand n33902(x33902, x33409, x33899);
  nand n33903(x33903, x33902, x33901);
  nand n33905(x33905, x33897, x33901);
  nand n33906(x33906, x33392, x33402);
  nand n33909(x33909, x33908, x33907);
  nand n33910(x33910, x33909, x33906);
  nand n33912(x33912, x33411, x33911);
  nand n33914(x33914, x33913, x33910);
  nand n33915(x33915, x33914, x33912);
  nand n33917(x33917, x33906, x33912);
  nand n33918(x33918, x33419, x33429);
  nand n33919(x33919, x33418, x33428);
  nand n33920(x33920, x33919, x33918);
  nand n33922(x33922, x33438, x33921);
  nand n33923(x33923, x33437, x33920);
  nand n33924(x33924, x33923, x33922);
  nand n33926(x33926, x33918, x33922);
  nand n33927(x33927, x33420, x33430);
  nand n33930(x33930, x33929, x33928);
  nand n33931(x33931, x33930, x33927);
  nand n33933(x33933, x33439, x33932);
  nand n33935(x33935, x33934, x33931);
  nand n33936(x33936, x33935, x33933);
  nand n33938(x33938, x33927, x33933);
  nand n33939(x33939, x33448, x33458);
  nand n33940(x33940, x33447, x33457);
  nand n33941(x33941, x33940, x33939);
  nand n33943(x33943, x33467, x33942);
  nand n33944(x33944, x33466, x33941);
  nand n33945(x33945, x33944, x33943);
  nand n33947(x33947, x33939, x33943);
  nand n33948(x33948, x33449, x33459);
  nand n33951(x33951, x33950, x33949);
  nand n33952(x33952, x33951, x33948);
  nand n33954(x33954, x33468, x33953);
  nand n33956(x33956, x33955, x33952);
  nand n33957(x33957, x33956, x33954);
  nand n33959(x33959, x33948, x33954);
  nand n33960(x33960, x33478, x33488);
  nand n33961(x33961, x33477, x33487);
  nand n33962(x33962, x33961, x33960);
  nand n33964(x33964, x33497, x33963);
  nand n33965(x33965, x33496, x33962);
  nand n33966(x33966, x33965, x33964);
  nand n33968(x33968, x33960, x33964);
  nand n33969(x33969, x33479, x33489);
  nand n33972(x33972, x33971, x33970);
  nand n33973(x33973, x33972, x33969);
  nand n33975(x33975, x33498, x33974);
  nand n33977(x33977, x33976, x33973);
  nand n33978(x33978, x33977, x33975);
  nand n33980(x33980, x33969, x33975);
  nand n33981(x33981, x33508, x33518);
  nand n33982(x33982, x33507, x33517);
  nand n33983(x33983, x33982, x33981);
  nand n33985(x33985, x33527, x33984);
  nand n33986(x33986, x33526, x33983);
  nand n33987(x33987, x33986, x33985);
  nand n33989(x33989, x33981, x33985);
  nand n33990(x33990, x33509, x33519);
  nand n33993(x33993, x33992, x33991);
  nand n33994(x33994, x33993, x33990);
  nand n33996(x33996, x33528, x33995);
  nand n33998(x33998, x33997, x33994);
  nand n33999(x33999, x33998, x33996);
  nand n34001(x34001, x33990, x33996);
  nand n34002(x34002, x33538, x33548);
  nand n34003(x34003, x33537, x33547);
  nand n34004(x34004, x34003, x34002);
  nand n34006(x34006, x33557, x34005);
  nand n34007(x34007, x33556, x34004);
  nand n34008(x34008, x34007, x34006);
  nand n34010(x34010, x34002, x34006);
  nand n34011(x34011, x33539, x33549);
  nand n34014(x34014, x34013, x34012);
  nand n34015(x34015, x34014, x34011);
  nand n34017(x34017, x33558, x34016);
  nand n34019(x34019, x34018, x34015);
  nand n34020(x34020, x34019, x34017);
  nand n34022(x34022, x34011, x34017);
  nand n34023(x34023, x33568, x33578);
  nand n34024(x34024, x33567, x33577);
  nand n34025(x34025, x34024, x34023);
  nand n34027(x34027, x33587, x34026);
  nand n34028(x34028, x33586, x34025);
  nand n34029(x34029, x34028, x34027);
  nand n34031(x34031, x34023, x34027);
  nand n34032(x34032, x33569, x33579);
  nand n34035(x34035, x34034, x34033);
  nand n34036(x34036, x34035, x34032);
  nand n34038(x34038, x33588, x34037);
  nand n34040(x34040, x34039, x34036);
  nand n34041(x34041, x34040, x34038);
  nand n34043(x34043, x34032, x34038);
  nand n34044(x34044, x33598, x33608);
  nand n34045(x34045, x33597, x33607);
  nand n34046(x34046, x34045, x34044);
  nand n34048(x34048, x33617, x34047);
  nand n34049(x34049, x33616, x34046);
  nand n34050(x34050, x34049, x34048);
  nand n34052(x34052, x34044, x34048);
  nand n34053(x34053, x33599, x33609);
  nand n34056(x34056, x34055, x34054);
  nand n34057(x34057, x34056, x34053);
  nand n34059(x34059, x33618, x34058);
  nand n34061(x34061, x34060, x34057);
  nand n34062(x34062, x34061, x34059);
  nand n34064(x34064, x33629, x33639);
  nand n34065(x34065, x33628, x33638);
  nand n34066(x34066, x34065, x34064);
  nand n34068(x34068, x33647, x34067);
  nand n34069(x34069, x33646, x34066);
  nand n34070(x34070, x34069, x34068);
  nand n34072(x34072, x84494, x84530);
  nand n34073(x34073, x33101, x33648);
  nand n34074(x34074, x34073, x34072);
  nand n34075(x34075, x84496, x84532);
  nand n34076(x34076, x33105, x33651);
  nand n34077(x34077, x34076, x34075);
  nand n34079(x34079, x33660, x84534);
  nand n34080(x34080, x33659, x33654);
  nand n34081(x34081, x34080, x34079);
  nand n34083(x34083, x84499, x84501);
  nand n34084(x34084, x33657, x33661);
  nand n34085(x34085, x34084, x34083);
  nand n34087(x34087, x33668, x34086);
  nand n34088(x34088, x33667, x34085);
  nand n34089(x34089, x34088, x34087);
  nand n34091(x34091, x34083, x34087);
  nand n34092(x34092, x84503, x84505);
  nand n34093(x34093, x33664, x33669);
  nand n34094(x34094, x34093, x34092);
  nand n34096(x34096, x33676, x34095);
  nand n34097(x34097, x33675, x34094);
  nand n34098(x34098, x34097, x34096);
  nand n34100(x34100, x34092, x34096);
  nand n34101(x34101, x84507, x84509);
  nand n34102(x34102, x33672, x33677);
  nand n34103(x34103, x34102, x34101);
  nand n34105(x34105, x33684, x34104);
  nand n34106(x34106, x33683, x34103);
  nand n34107(x34107, x34106, x34105);
  nand n34109(x34109, x34101, x34105);
  nand n34110(x34110, x84511, x84513);
  nand n34111(x34111, x33680, x33685);
  nand n34112(x34112, x34111, x34110);
  nand n34114(x34114, x33692, x34113);
  nand n34115(x34115, x33691, x34112);
  nand n34116(x34116, x34115, x34114);
  nand n34118(x34118, x34110, x34114);
  nand n34119(x34119, x84515, x84517);
  nand n34120(x34120, x33688, x33693);
  nand n34121(x34121, x34120, x34119);
  nand n34123(x34123, x33700, x34122);
  nand n34124(x34124, x33699, x34121);
  nand n34125(x34125, x34124, x34123);
  nand n34127(x34127, x34119, x34123);
  nand n34128(x34128, x33708, x84376);
  nand n34129(x34129, x33707, x29180);
  nand n34130(x34130, x34129, x34128);
  nand n34133(x34133, x84519, x33709);
  nand n34135(x34135, x33696, x34134);
  nand n34136(x34136, x34135, x34133);
  nand n34138(x34138, x33714, x34137);
  nand n34139(x34139, x33713, x34136);
  nand n34140(x34140, x34139, x34138);
  nand n34142(x34142, x34133, x34138);
  nand n34143(x34143, x33722, x84379);
  nand n34144(x34144, x33721, x30320);
  nand n34145(x34145, x34144, x34143);
  nand n34148(x34148, x84521, x33723);
  nand n34150(x34150, x33710, x34149);
  nand n34151(x34151, x34150, x34148);
  nand n34153(x34153, x33728, x34152);
  nand n34154(x34154, x33727, x34151);
  nand n34155(x34155, x34154, x34153);
  nand n34157(x34157, x34148, x34153);
  nand n34158(x34158, x33736, x84382);
  nand n34159(x34159, x33735, x30362);
  nand n34160(x34160, x34159, x34158);
  nand n34163(x34163, x84523, x33737);
  nand n34165(x34165, x33724, x34164);
  nand n34166(x34166, x34165, x34163);
  nand n34168(x34168, x33742, x34167);
  nand n34169(x34169, x33741, x34166);
  nand n34170(x34170, x34169, x34168);
  nand n34172(x34172, x34163, x34168);
  nand n34173(x34173, x33750, x84387);
  nand n34174(x34174, x33749, x31716);
  nand n34175(x34175, x34174, x34173);
  nand n34178(x34178, x84525, x33751);
  nand n34180(x34180, x33738, x34179);
  nand n34181(x34181, x34180, x34178);
  nand n34183(x34183, x33756, x34182);
  nand n34184(x34184, x33755, x34181);
  nand n34185(x34185, x34184, x34183);
  nand n34187(x34187, x34178, x34183);
  nand n34188(x34188, x33764, x84394);
  nand n34189(x34189, x33763, x31744);
  nand n34190(x34190, x34189, x34188);
  nand n34193(x34193, x84527, x33765);
  nand n34195(x34195, x33752, x34194);
  nand n34196(x34196, x34195, x34193);
  nand n34198(x34198, x33774, x34197);
  nand n34199(x34199, x33773, x34196);
  nand n34200(x34200, x34199, x34198);
  nand n34202(x34202, x34193, x34198);
  nand n34203(x34203, x33783, x84401);
  nand n34204(x34204, x33782, x31778);
  nand n34205(x34205, x34204, x34203);
  nand n34208(x34208, x33775, x33784);
  nand n34211(x34211, x34210, x34209);
  nand n34212(x34212, x34211, x34208);
  nand n34214(x34214, x33794, x34213);
  nand n34215(x34215, x33793, x34212);
  nand n34216(x34216, x34215, x34214);
  nand n34218(x34218, x34208, x34214);
  nand n34219(x34219, x33803, x84408);
  nand n34220(x34220, x33802, x31817);
  nand n34221(x34221, x34220, x34219);
  nand n34224(x34224, x33795, x33804);
  nand n34227(x34227, x34226, x34225);
  nand n34228(x34228, x34227, x34224);
  nand n34230(x34230, x33814, x34229);
  nand n34231(x34231, x33813, x34228);
  nand n34232(x34232, x34231, x34230);
  nand n34234(x34234, x34224, x34230);
  nand n34235(x34235, x33823, x84415);
  nand n34236(x34236, x33822, x31857);
  nand n34237(x34237, x34236, x34235);
  nand n34240(x34240, x33815, x33824);
  nand n34243(x34243, x34242, x34241);
  nand n34244(x34244, x34243, x34240);
  nand n34246(x34246, x33834, x34245);
  nand n34247(x34247, x33833, x34244);
  nand n34248(x34248, x34247, x34246);
  nand n34250(x34250, x34240, x34246);
  nand n34251(x34251, x33843, x84421);
  nand n34252(x34252, x33842, x31897);
  nand n34253(x34253, x34252, x34251);
  nand n34256(x34256, x33835, x33844);
  nand n34259(x34259, x34258, x34257);
  nand n34260(x34260, x34259, x34256);
  nand n34262(x34262, x33854, x34261);
  nand n34263(x34263, x33853, x34260);
  nand n34264(x34264, x34263, x34262);
  nand n34266(x34266, x34256, x34262);
  nand n34267(x34267, x33863, x84427);
  nand n34268(x34268, x33862, x32715);
  nand n34269(x34269, x34268, x34267);
  nand n34272(x34272, x33855, x33864);
  nand n34275(x34275, x34274, x34273);
  nand n34276(x34276, x34275, x34272);
  nand n34278(x34278, x33874, x34277);
  nand n34279(x34279, x33873, x34276);
  nand n34280(x34280, x34279, x34278);
  nand n34282(x34282, x34272, x34278);
  nand n34283(x34283, x33883, x84434);
  nand n34284(x34284, x33882, x32742);
  nand n34285(x34285, x34284, x34283);
  nand n34288(x34288, x33875, x33884);
  nand n34291(x34291, x34290, x34289);
  nand n34292(x34292, x34291, x34288);
  nand n34294(x34294, x33895, x34293);
  nand n34295(x34295, x33894, x34292);
  nand n34296(x34296, x34295, x34294);
  nand n34298(x34298, x34288, x34294);
  nand n34299(x34299, x33904, x84441);
  nand n34300(x34300, x33903, x32769);
  nand n34301(x34301, x34300, x34299);
  nand n34304(x34304, x33896, x33905);
  nand n34307(x34307, x34306, x34305);
  nand n34308(x34308, x34307, x34304);
  nand n34310(x34310, x33916, x34309);
  nand n34311(x34311, x33915, x34308);
  nand n34312(x34312, x34311, x34310);
  nand n34314(x34314, x34304, x34310);
  nand n34315(x34315, x33925, x84446);
  nand n34316(x34316, x33924, x32802);
  nand n34317(x34317, x34316, x34315);
  nand n34320(x34320, x33917, x33926);
  nand n34323(x34323, x34322, x34321);
  nand n34324(x34324, x34323, x34320);
  nand n34326(x34326, x33937, x34325);
  nand n34327(x34327, x33936, x34324);
  nand n34328(x34328, x34327, x34326);
  nand n34330(x34330, x34320, x34326);
  nand n34331(x34331, x33946, x84449);
  nand n34332(x34332, x33945, x32840);
  nand n34333(x34333, x34332, x34331);
  nand n34336(x34336, x33938, x33947);
  nand n34339(x34339, x34338, x34337);
  nand n34340(x34340, x34339, x34336);
  nand n34342(x34342, x33958, x34341);
  nand n34343(x34343, x33957, x34340);
  nand n34344(x34344, x34343, x34342);
  nand n34346(x34346, x34336, x34342);
  nand n34347(x34347, x33967, x84452);
  nand n34348(x34348, x33966, x32878);
  nand n34349(x34349, x34348, x34347);
  nand n34352(x34352, x33959, x33968);
  nand n34355(x34355, x34354, x34353);
  nand n34356(x34356, x34355, x34352);
  nand n34358(x34358, x33979, x34357);
  nand n34359(x34359, x33978, x34356);
  nand n34360(x34360, x34359, x34358);
  nand n34362(x34362, x34352, x34358);
  nand n34363(x34363, x33988, x84455);
  nand n34364(x34364, x33987, x32917);
  nand n34365(x34365, x34364, x34363);
  nand n34368(x34368, x33980, x33989);
  nand n34371(x34371, x34370, x34369);
  nand n34372(x34372, x34371, x34368);
  nand n34374(x34374, x34000, x34373);
  nand n34375(x34375, x33999, x34372);
  nand n34376(x34376, x34375, x34374);
  nand n34378(x34378, x34368, x34374);
  nand n34379(x34379, x34009, x84458);
  nand n34380(x34380, x34008, x32957);
  nand n34381(x34381, x34380, x34379);
  nand n34384(x34384, x34001, x34010);
  nand n34387(x34387, x34386, x34385);
  nand n34388(x34388, x34387, x34384);
  nand n34390(x34390, x34021, x34389);
  nand n34391(x34391, x34020, x34388);
  nand n34392(x34392, x34391, x34390);
  nand n34394(x34394, x34384, x34390);
  nand n34395(x34395, x34030, x84461);
  nand n34396(x34396, x34029, x32997);
  nand n34397(x34397, x34396, x34395);
  nand n34400(x34400, x34022, x34031);
  nand n34403(x34403, x34402, x34401);
  nand n34404(x34404, x34403, x34400);
  nand n34406(x34406, x34042, x34405);
  nand n34407(x34407, x34041, x34404);
  nand n34408(x34408, x34407, x34406);
  nand n34410(x34410, x34400, x34406);
  nand n34411(x34411, x34051, x33047);
  nand n34412(x34412, x34050, x33046);
  nand n34413(x34413, x34412, x34411);
  nand n34416(x34416, x34043, x34052);
  nand n34419(x34419, x34418, x34417);
  nand n34420(x34420, x34419, x34416);
  nand n34422(x34422, x34063, x34421);
  nand n34423(x34423, x34062, x34420);
  nand n34424(x34424, x34423, x34422);
  nand n34426(x34426, x34071, x33094);
  nand n34427(x34427, x34070, x33093);
  nand n34428(x34428, x34427, x34426);
  nand n34430(x34430, x84528, x84540);
  nand n34431(x34431, x33100, x33095);
  nand n34432(x34432, x34431, x34430);
  nand n34433(x34433, x34078, x84543);
  nand n34434(x34434, x34077, x34072);
  nand n34435(x34435, x34434, x34433);
  nand n34436(x34436, x34082, x84545);
  nand n34437(x34437, x34081, x34075);
  nand n34438(x34438, x34437, x34436);
  nand n34440(x34440, x34090, x84547);
  nand n34441(x34441, x34089, x34079);
  nand n34442(x34442, x34441, x34440);
  nand n34445(x34445, x34099, x34091);
  nand n34446(x34446, x34098, x34444);
  nand n34447(x34447, x34446, x34445);
  nand n34450(x34450, x34108, x34100);
  nand n34451(x34451, x34107, x34449);
  nand n34452(x34452, x34451, x34450);
  nand n34455(x34455, x34117, x34109);
  nand n34456(x34456, x34116, x34454);
  nand n34457(x34457, x34456, x34455);
  nand n34460(x34460, x34126, x34118);
  nand n34461(x34461, x34125, x34459);
  nand n34462(x34462, x34461, x34460);
  nand n34464(x34464, x34127, x34132);
  nand n34466(x34466, x34465, x34128);
  nand n34467(x34467, x34466, x34464);
  nand n34469(x34469, x34141, x34468);
  nand n34470(x34470, x34140, x34467);
  nand n34471(x34471, x34470, x34469);
  nand n34473(x34473, x34464, x34469);
  nand n34474(x34474, x34142, x34147);
  nand n34476(x34476, x34475, x34143);
  nand n34477(x34477, x34476, x34474);
  nand n34479(x34479, x34156, x34478);
  nand n34480(x34480, x34155, x34477);
  nand n34481(x34481, x34480, x34479);
  nand n34483(x34483, x34474, x34479);
  nand n34484(x34484, x34157, x34162);
  nand n34486(x34486, x34485, x34158);
  nand n34487(x34487, x34486, x34484);
  nand n34489(x34489, x34171, x34488);
  nand n34490(x34490, x34170, x34487);
  nand n34491(x34491, x34490, x34489);
  nand n34493(x34493, x34484, x34489);
  nand n34494(x34494, x34172, x34177);
  nand n34496(x34496, x34495, x34173);
  nand n34497(x34497, x34496, x34494);
  nand n34499(x34499, x34186, x34498);
  nand n34500(x34500, x34185, x34497);
  nand n34501(x34501, x34500, x34499);
  nand n34503(x34503, x34494, x34499);
  nand n34504(x34504, x34187, x34192);
  nand n34506(x34506, x34505, x34188);
  nand n34507(x34507, x34506, x34504);
  nand n34509(x34509, x34201, x34508);
  nand n34510(x34510, x34200, x34507);
  nand n34511(x34511, x34510, x34509);
  nand n34513(x34513, x34504, x34509);
  nand n34514(x34514, x34202, x34207);
  nand n34516(x34516, x34515, x34203);
  nand n34517(x34517, x34516, x34514);
  nand n34519(x34519, x34217, x34518);
  nand n34520(x34520, x34216, x34517);
  nand n34521(x34521, x34520, x34519);
  nand n34523(x34523, x34514, x34519);
  nand n34524(x34524, x34218, x34223);
  nand n34526(x34526, x34525, x34219);
  nand n34527(x34527, x34526, x34524);
  nand n34529(x34529, x34233, x34528);
  nand n34530(x34530, x34232, x34527);
  nand n34531(x34531, x34530, x34529);
  nand n34533(x34533, x34524, x34529);
  nand n34534(x34534, x34234, x34239);
  nand n34536(x34536, x34535, x34235);
  nand n34537(x34537, x34536, x34534);
  nand n34539(x34539, x34249, x34538);
  nand n34540(x34540, x34248, x34537);
  nand n34541(x34541, x34540, x34539);
  nand n34543(x34543, x34534, x34539);
  nand n34544(x34544, x34250, x34255);
  nand n34546(x34546, x34545, x34251);
  nand n34547(x34547, x34546, x34544);
  nand n34549(x34549, x34265, x34548);
  nand n34550(x34550, x34264, x34547);
  nand n34551(x34551, x34550, x34549);
  nand n34553(x34553, x34544, x34549);
  nand n34554(x34554, x34266, x34271);
  nand n34556(x34556, x34555, x34267);
  nand n34557(x34557, x34556, x34554);
  nand n34559(x34559, x34281, x34558);
  nand n34560(x34560, x34280, x34557);
  nand n34561(x34561, x34560, x34559);
  nand n34563(x34563, x34554, x34559);
  nand n34564(x34564, x34282, x34287);
  nand n34566(x34566, x34565, x34283);
  nand n34567(x34567, x34566, x34564);
  nand n34569(x34569, x34297, x34568);
  nand n34570(x34570, x34296, x34567);
  nand n34571(x34571, x34570, x34569);
  nand n34573(x34573, x34564, x34569);
  nand n34574(x34574, x34298, x34303);
  nand n34576(x34576, x34575, x34299);
  nand n34577(x34577, x34576, x34574);
  nand n34579(x34579, x34313, x34578);
  nand n34580(x34580, x34312, x34577);
  nand n34581(x34581, x34580, x34579);
  nand n34583(x34583, x34574, x34579);
  nand n34584(x34584, x34314, x34319);
  nand n34586(x34586, x34585, x34315);
  nand n34587(x34587, x34586, x34584);
  nand n34589(x34589, x34329, x34588);
  nand n34590(x34590, x34328, x34587);
  nand n34591(x34591, x34590, x34589);
  nand n34593(x34593, x34584, x34589);
  nand n34594(x34594, x34330, x34335);
  nand n34596(x34596, x34595, x34331);
  nand n34597(x34597, x34596, x34594);
  nand n34599(x34599, x34345, x34598);
  nand n34600(x34600, x34344, x34597);
  nand n34601(x34601, x34600, x34599);
  nand n34603(x34603, x34594, x34599);
  nand n34604(x34604, x34346, x34351);
  nand n34606(x34606, x34605, x34347);
  nand n34607(x34607, x34606, x34604);
  nand n34609(x34609, x34361, x34608);
  nand n34610(x34610, x34360, x34607);
  nand n34611(x34611, x34610, x34609);
  nand n34613(x34613, x34604, x34609);
  nand n34614(x34614, x34362, x34367);
  nand n34616(x34616, x34615, x34363);
  nand n34617(x34617, x34616, x34614);
  nand n34619(x34619, x34377, x34618);
  nand n34620(x34620, x34376, x34617);
  nand n34621(x34621, x34620, x34619);
  nand n34623(x34623, x34614, x34619);
  nand n34624(x34624, x34378, x34383);
  nand n34626(x34626, x34625, x34379);
  nand n34627(x34627, x34626, x34624);
  nand n34629(x34629, x34393, x34628);
  nand n34630(x34630, x34392, x34627);
  nand n34631(x34631, x34630, x34629);
  nand n34633(x34633, x34624, x34629);
  nand n34634(x34634, x34394, x34399);
  nand n34636(x34636, x34635, x34395);
  nand n34637(x34637, x34636, x34634);
  nand n34639(x34639, x34409, x34638);
  nand n34640(x34640, x34408, x34637);
  nand n34641(x34641, x34640, x34639);
  nand n34643(x34643, x34634, x34639);
  nand n34644(x34644, x34410, x34415);
  nand n34646(x34646, x34645, x34411);
  nand n34647(x34647, x34646, x34644);
  nand n34649(x34649, x34425, x34648);
  nand n34650(x34650, x34424, x34647);
  nand n34651(x34651, x34650, x34649);
  nand n34653(x34653, x84541, x84542);
  nand n34654(x34654, x34430, x33098);
  nand n34655(x34655, x34654, x34653);
  nand n34657(x34657, x84529, x34656);
  nand n34658(x34658, x33650, x34655);
  nand n34659(x34659, x34658, x34657);
  nand n34660(x34660, x34653, x34657);
  nand n34661(x34661, x84531, x84553);
  nand n34662(x34662, x33653, x34074);
  nand n34663(x34663, x34662, x34661);
  nand n34665(x34665, x84533, x84555);
  nand n34666(x34666, x33656, x34435);
  nand n34667(x34667, x34666, x34665);
  nand n34669(x34669, x84544, x34439);
  nand n34670(x34670, x34433, x34438);
  nand n34671(x34671, x34670, x34669);
  nand n34673(x34673, x84535, x34672);
  nand n34674(x34674, x33663, x34671);
  nand n34675(x34675, x34674, x34673);
  nand n34677(x34677, x34669, x34673);
  nand n34678(x34678, x84546, x34443);
  nand n34679(x34679, x34436, x34442);
  nand n34680(x34680, x34679, x34678);
  nand n34682(x34682, x84536, x34681);
  nand n34683(x34683, x33671, x34680);
  nand n34684(x34684, x34683, x34682);
  nand n34686(x34686, x34678, x34682);
  nand n34687(x34687, x84548, x34448);
  nand n34688(x34688, x34440, x34447);
  nand n34689(x34689, x34688, x34687);
  nand n34691(x34691, x84537, x34690);
  nand n34692(x34692, x33679, x34689);
  nand n34693(x34693, x34692, x34691);
  nand n34695(x34695, x34687, x34691);
  nand n34696(x34696, x84549, x34453);
  nand n34697(x34697, x34445, x34452);
  nand n34698(x34698, x34697, x34696);
  nand n34700(x34700, x84538, x34699);
  nand n34701(x34701, x33687, x34698);
  nand n34702(x34702, x34701, x34700);
  nand n34704(x34704, x34696, x34700);
  nand n34705(x34705, x84550, x34458);
  nand n34706(x34706, x34450, x34457);
  nand n34707(x34707, x34706, x34705);
  nand n34709(x34709, x84539, x34708);
  nand n34710(x34710, x33695, x34707);
  nand n34711(x34711, x34710, x34709);
  nand n34713(x34713, x34705, x34709);
  nand n34714(x34714, x84551, x34463);
  nand n34715(x34715, x34455, x34462);
  nand n34716(x34716, x34715, x34714);
  nand n34718(x34718, x34131, x34717);
  nand n34719(x34719, x34130, x34716);
  nand n34720(x34720, x34719, x34718);
  nand n34722(x34722, x34714, x34718);
  nand n34723(x34723, x84552, x34472);
  nand n34724(x34724, x34460, x34471);
  nand n34725(x34725, x34724, x34723);
  nand n34727(x34727, x34146, x34726);
  nand n34728(x34728, x34145, x34725);
  nand n34729(x34729, x34728, x34727);
  nand n34731(x34731, x34723, x34727);
  nand n34732(x34732, x34473, x34482);
  nand n34734(x34734, x34733, x34481);
  nand n34735(x34735, x34734, x34732);
  nand n34737(x34737, x34161, x34736);
  nand n34738(x34738, x34160, x34735);
  nand n34739(x34739, x34738, x34737);
  nand n34741(x34741, x34732, x34737);
  nand n34742(x34742, x34483, x34492);
  nand n34744(x34744, x34743, x34491);
  nand n34745(x34745, x34744, x34742);
  nand n34747(x34747, x34176, x34746);
  nand n34748(x34748, x34175, x34745);
  nand n34749(x34749, x34748, x34747);
  nand n34751(x34751, x34742, x34747);
  nand n34752(x34752, x34493, x34502);
  nand n34754(x34754, x34753, x34501);
  nand n34755(x34755, x34754, x34752);
  nand n34757(x34757, x34191, x34756);
  nand n34758(x34758, x34190, x34755);
  nand n34759(x34759, x34758, x34757);
  nand n34761(x34761, x34752, x34757);
  nand n34762(x34762, x34503, x34512);
  nand n34764(x34764, x34763, x34511);
  nand n34765(x34765, x34764, x34762);
  nand n34767(x34767, x34206, x34766);
  nand n34768(x34768, x34205, x34765);
  nand n34769(x34769, x34768, x34767);
  nand n34771(x34771, x34762, x34767);
  nand n34772(x34772, x34513, x34522);
  nand n34774(x34774, x34773, x34521);
  nand n34775(x34775, x34774, x34772);
  nand n34777(x34777, x34222, x34776);
  nand n34778(x34778, x34221, x34775);
  nand n34779(x34779, x34778, x34777);
  nand n34781(x34781, x34772, x34777);
  nand n34782(x34782, x34523, x34532);
  nand n34784(x34784, x34783, x34531);
  nand n34785(x34785, x34784, x34782);
  nand n34787(x34787, x34238, x34786);
  nand n34788(x34788, x34237, x34785);
  nand n34789(x34789, x34788, x34787);
  nand n34791(x34791, x34782, x34787);
  nand n34792(x34792, x34533, x34542);
  nand n34794(x34794, x34793, x34541);
  nand n34795(x34795, x34794, x34792);
  nand n34797(x34797, x34254, x34796);
  nand n34798(x34798, x34253, x34795);
  nand n34799(x34799, x34798, x34797);
  nand n34801(x34801, x34792, x34797);
  nand n34802(x34802, x34543, x34552);
  nand n34804(x34804, x34803, x34551);
  nand n34805(x34805, x34804, x34802);
  nand n34807(x34807, x34270, x34806);
  nand n34808(x34808, x34269, x34805);
  nand n34809(x34809, x34808, x34807);
  nand n34811(x34811, x34802, x34807);
  nand n34812(x34812, x34553, x34562);
  nand n34814(x34814, x34813, x34561);
  nand n34815(x34815, x34814, x34812);
  nand n34817(x34817, x34286, x34816);
  nand n34818(x34818, x34285, x34815);
  nand n34819(x34819, x34818, x34817);
  nand n34821(x34821, x34812, x34817);
  nand n34822(x34822, x34563, x34572);
  nand n34824(x34824, x34823, x34571);
  nand n34825(x34825, x34824, x34822);
  nand n34827(x34827, x34302, x34826);
  nand n34828(x34828, x34301, x34825);
  nand n34829(x34829, x34828, x34827);
  nand n34831(x34831, x34822, x34827);
  nand n34832(x34832, x34573, x34582);
  nand n34834(x34834, x34833, x34581);
  nand n34835(x34835, x34834, x34832);
  nand n34837(x34837, x34318, x34836);
  nand n34838(x34838, x34317, x34835);
  nand n34839(x34839, x34838, x34837);
  nand n34841(x34841, x34832, x34837);
  nand n34842(x34842, x34583, x34592);
  nand n34844(x34844, x34843, x34591);
  nand n34845(x34845, x34844, x34842);
  nand n34847(x34847, x34334, x34846);
  nand n34848(x34848, x34333, x34845);
  nand n34849(x34849, x34848, x34847);
  nand n34851(x34851, x34842, x34847);
  nand n34852(x34852, x34593, x34602);
  nand n34854(x34854, x34853, x34601);
  nand n34855(x34855, x34854, x34852);
  nand n34857(x34857, x34350, x34856);
  nand n34858(x34858, x34349, x34855);
  nand n34859(x34859, x34858, x34857);
  nand n34861(x34861, x34852, x34857);
  nand n34862(x34862, x34603, x34612);
  nand n34864(x34864, x34863, x34611);
  nand n34865(x34865, x34864, x34862);
  nand n34867(x34867, x34366, x34866);
  nand n34868(x34868, x34365, x34865);
  nand n34869(x34869, x34868, x34867);
  nand n34871(x34871, x34862, x34867);
  nand n34872(x34872, x34613, x34622);
  nand n34874(x34874, x34873, x34621);
  nand n34875(x34875, x34874, x34872);
  nand n34877(x34877, x34382, x34876);
  nand n34878(x34878, x34381, x34875);
  nand n34879(x34879, x34878, x34877);
  nand n34881(x34881, x34872, x34877);
  nand n34882(x34882, x34623, x34632);
  nand n34884(x34884, x34883, x34631);
  nand n34885(x34885, x34884, x34882);
  nand n34887(x34887, x34398, x34886);
  nand n34888(x34888, x34397, x34885);
  nand n34889(x34889, x34888, x34887);
  nand n34891(x34891, x34882, x34887);
  nand n34892(x34892, x34633, x34642);
  nand n34894(x34894, x34893, x34641);
  nand n34895(x34895, x34894, x34892);
  nand n34897(x34897, x34414, x34896);
  nand n34898(x34898, x34413, x34895);
  nand n34899(x34899, x34898, x34897);
  nand n34901(x34901, x34892, x34897);
  nand n34902(x34902, x34643, x34652);
  nand n34904(x34904, x34903, x34651);
  nand n34905(x34905, x34904, x34902);
  nand n34907(x34907, x34429, x34906);
  nand n34908(x34908, x34428, x34905);
  nand n34909(x34909, x34908, x34907);
  nand n34911(x34911, x34660, x34664);
  nand n34913(x34913, x34912, x34663);
  nand n34914(x34914, x34913, x34911);
  nand n34915(x34915, x84554, x34668);
  nand n34916(x34916, x34661, x34667);
  nand n34917(x34917, x34916, x34915);
  nand n34919(x34919, x84556, x34676);
  nand n34920(x34920, x34665, x34675);
  nand n34921(x34921, x34920, x34919);
  nand n34923(x34923, x34677, x34685);
  nand n34925(x34925, x34924, x34684);
  nand n34926(x34926, x34925, x34923);
  nand n34928(x34928, x34686, x34694);
  nand n34930(x34930, x34929, x34693);
  nand n34931(x34931, x34930, x34928);
  nand n34933(x34933, x34695, x34703);
  nand n34935(x34935, x34934, x34702);
  nand n34936(x34936, x34935, x34933);
  nand n34938(x34938, x34704, x34712);
  nand n34940(x34940, x34939, x34711);
  nand n34941(x34941, x34940, x34938);
  nand n34943(x34943, x34713, x34721);
  nand n34945(x34945, x34944, x34720);
  nand n34946(x34946, x34945, x34943);
  nand n34948(x34948, x34722, x34730);
  nand n34950(x34950, x34949, x34729);
  nand n34951(x34951, x34950, x34948);
  nand n34953(x34953, x34731, x34740);
  nand n34955(x34955, x34954, x34739);
  nand n34956(x34956, x34955, x34953);
  nand n34958(x34958, x34741, x34750);
  nand n34960(x34960, x34959, x34749);
  nand n34961(x34961, x34960, x34958);
  nand n34963(x34963, x34751, x34760);
  nand n34965(x34965, x34964, x34759);
  nand n34966(x34966, x34965, x34963);
  nand n34968(x34968, x34761, x34770);
  nand n34970(x34970, x34969, x34769);
  nand n34971(x34971, x34970, x34968);
  nand n34973(x34973, x34771, x34780);
  nand n34975(x34975, x34974, x34779);
  nand n34976(x34976, x34975, x34973);
  nand n34978(x34978, x34781, x34790);
  nand n34980(x34980, x34979, x34789);
  nand n34981(x34981, x34980, x34978);
  nand n34983(x34983, x34791, x34800);
  nand n34985(x34985, x34984, x34799);
  nand n34986(x34986, x34985, x34983);
  nand n34988(x34988, x34801, x34810);
  nand n34990(x34990, x34989, x34809);
  nand n34991(x34991, x34990, x34988);
  nand n34993(x34993, x34811, x34820);
  nand n34995(x34995, x34994, x34819);
  nand n34996(x34996, x34995, x34993);
  nand n34998(x34998, x34821, x34830);
  nand n35000(x35000, x34999, x34829);
  nand n35001(x35001, x35000, x34998);
  nand n35003(x35003, x34831, x34840);
  nand n35005(x35005, x35004, x34839);
  nand n35006(x35006, x35005, x35003);
  nand n35008(x35008, x34841, x34850);
  nand n35010(x35010, x35009, x34849);
  nand n35011(x35011, x35010, x35008);
  nand n35013(x35013, x34851, x34860);
  nand n35015(x35015, x35014, x34859);
  nand n35016(x35016, x35015, x35013);
  nand n35018(x35018, x34861, x34870);
  nand n35020(x35020, x35019, x34869);
  nand n35021(x35021, x35020, x35018);
  nand n35023(x35023, x34871, x34880);
  nand n35025(x35025, x35024, x34879);
  nand n35026(x35026, x35025, x35023);
  nand n35028(x35028, x34881, x34890);
  nand n35030(x35030, x35029, x34889);
  nand n35031(x35031, x35030, x35028);
  nand n35033(x35033, x34891, x34900);
  nand n35035(x35035, x35034, x34899);
  nand n35036(x35036, x35035, x35033);
  nand n35038(x35038, x34901, x34910);
  nand n35040(x35040, x35039, x34909);
  nand n35041(x35041, x35040, x35038);
  nand n35068(x35068, x34918, x35043);
  nand n35069(x35069, x35068, x34915);
  nand n35070(x35070, x34922, x35044);
  nand n35071(x35071, x35070, x34919);
  nand n35072(x35072, x34922, x34918);
  nand n35074(x35074, x34927, x35045);
  nand n35075(x35075, x35074, x34923);
  nand n35076(x35076, x34927, x34922);
  nand n35078(x35078, x34932, x35046);
  nand n35079(x35079, x35078, x34928);
  nand n35080(x35080, x34932, x34927);
  nand n35082(x35082, x34937, x35047);
  nand n35083(x35083, x35082, x34933);
  nand n35084(x35084, x34937, x34932);
  nand n35086(x35086, x34942, x35048);
  nand n35087(x35087, x35086, x34938);
  nand n35088(x35088, x34942, x34937);
  nand n35090(x35090, x34947, x35049);
  nand n35091(x35091, x35090, x34943);
  nand n35092(x35092, x34947, x34942);
  nand n35094(x35094, x34952, x35050);
  nand n35095(x35095, x35094, x34948);
  nand n35096(x35096, x34952, x34947);
  nand n35098(x35098, x34957, x35051);
  nand n35099(x35099, x35098, x34953);
  nand n35100(x35100, x34957, x34952);
  nand n35102(x35102, x34962, x35052);
  nand n35103(x35103, x35102, x34958);
  nand n35104(x35104, x34962, x34957);
  nand n35106(x35106, x34967, x35053);
  nand n35107(x35107, x35106, x34963);
  nand n35108(x35108, x34967, x34962);
  nand n35110(x35110, x34972, x35054);
  nand n35111(x35111, x35110, x34968);
  nand n35112(x35112, x34972, x34967);
  nand n35114(x35114, x34977, x35055);
  nand n35115(x35115, x35114, x34973);
  nand n35116(x35116, x34977, x34972);
  nand n35118(x35118, x34982, x35056);
  nand n35119(x35119, x35118, x34978);
  nand n35120(x35120, x34982, x34977);
  nand n35122(x35122, x34987, x35057);
  nand n35123(x35123, x35122, x34983);
  nand n35124(x35124, x34987, x34982);
  nand n35126(x35126, x34992, x35058);
  nand n35127(x35127, x35126, x34988);
  nand n35128(x35128, x34992, x34987);
  nand n35130(x35130, x34997, x35059);
  nand n35131(x35131, x35130, x34993);
  nand n35132(x35132, x34997, x34992);
  nand n35134(x35134, x35002, x35060);
  nand n35135(x35135, x35134, x34998);
  nand n35136(x35136, x35002, x34997);
  nand n35138(x35138, x35007, x35061);
  nand n35139(x35139, x35138, x35003);
  nand n35140(x35140, x35007, x35002);
  nand n35142(x35142, x35012, x35062);
  nand n35143(x35143, x35142, x35008);
  nand n35144(x35144, x35012, x35007);
  nand n35146(x35146, x35017, x35063);
  nand n35147(x35147, x35146, x35013);
  nand n35148(x35148, x35017, x35012);
  nand n35150(x35150, x35022, x35064);
  nand n35151(x35151, x35150, x35018);
  nand n35152(x35152, x35022, x35017);
  nand n35154(x35154, x35027, x35065);
  nand n35155(x35155, x35154, x35023);
  nand n35156(x35156, x35027, x35022);
  nand n35158(x35158, x35032, x35066);
  nand n35159(x35159, x35158, x35028);
  nand n35160(x35160, x35032, x35027);
  nand n35162(x35162, x35037, x35067);
  nand n35163(x35163, x35162, x35033);
  nand n35164(x35164, x35037, x35032);
  nand n35167(x35167, x35073, x35043);
  nand n35169(x35169, x35167, x35168);
  nand n35170(x35170, x35077, x35069);
  nand n35172(x35172, x35170, x35171);
  nand n35173(x35173, x35081, x35071);
  nand n35175(x35175, x35173, x35174);
  nand n35176(x35176, x35081, x35073);
  nand n35178(x35178, x35085, x35075);
  nand n35180(x35180, x35178, x35179);
  nand n35181(x35181, x35085, x35077);
  nand n35183(x35183, x35089, x35079);
  nand n35185(x35185, x35183, x35184);
  nand n35186(x35186, x35089, x35081);
  nand n35188(x35188, x35093, x35083);
  nand n35190(x35190, x35188, x35189);
  nand n35191(x35191, x35093, x35085);
  nand n35193(x35193, x35097, x35087);
  nand n35195(x35195, x35193, x35194);
  nand n35196(x35196, x35097, x35089);
  nand n35198(x35198, x35101, x35091);
  nand n35200(x35200, x35198, x35199);
  nand n35201(x35201, x35101, x35093);
  nand n35203(x35203, x35105, x35095);
  nand n35205(x35205, x35203, x35204);
  nand n35206(x35206, x35105, x35097);
  nand n35208(x35208, x35109, x35099);
  nand n35210(x35210, x35208, x35209);
  nand n35211(x35211, x35109, x35101);
  nand n35213(x35213, x35113, x35103);
  nand n35215(x35215, x35213, x35214);
  nand n35216(x35216, x35113, x35105);
  nand n35218(x35218, x35117, x35107);
  nand n35220(x35220, x35218, x35219);
  nand n35221(x35221, x35117, x35109);
  nand n35223(x35223, x35121, x35111);
  nand n35225(x35225, x35223, x35224);
  nand n35226(x35226, x35121, x35113);
  nand n35228(x35228, x35125, x35115);
  nand n35230(x35230, x35228, x35229);
  nand n35231(x35231, x35125, x35117);
  nand n35233(x35233, x35129, x35119);
  nand n35235(x35235, x35233, x35234);
  nand n35236(x35236, x35129, x35121);
  nand n35238(x35238, x35133, x35123);
  nand n35240(x35240, x35238, x35239);
  nand n35241(x35241, x35133, x35125);
  nand n35243(x35243, x35137, x35127);
  nand n35245(x35245, x35243, x35244);
  nand n35246(x35246, x35137, x35129);
  nand n35248(x35248, x35141, x35131);
  nand n35250(x35250, x35248, x35249);
  nand n35251(x35251, x35141, x35133);
  nand n35253(x35253, x35145, x35135);
  nand n35255(x35255, x35253, x35254);
  nand n35256(x35256, x35145, x35137);
  nand n35258(x35258, x35149, x35139);
  nand n35260(x35260, x35258, x35259);
  nand n35261(x35261, x35149, x35141);
  nand n35263(x35263, x35153, x35143);
  nand n35265(x35265, x35263, x35264);
  nand n35266(x35266, x35153, x35145);
  nand n35268(x35268, x35157, x35147);
  nand n35270(x35270, x35268, x35269);
  nand n35271(x35271, x35157, x35149);
  nand n35273(x35273, x35161, x35151);
  nand n35275(x35275, x35273, x35274);
  nand n35276(x35276, x35161, x35153);
  nand n35278(x35278, x35165, x35155);
  nand n35280(x35280, x35278, x35279);
  nand n35281(x35281, x35165, x35157);
  nand n35285(x35285, x35177, x35043);
  nand n35287(x35287, x35285, x35286);
  nand n35288(x35288, x35182, x35069);
  nand n35290(x35290, x35288, x35289);
  nand n35291(x35291, x35187, x35169);
  nand n35293(x35293, x35291, x35292);
  nand n35294(x35294, x35192, x35172);
  nand n35296(x35296, x35294, x35295);
  nand n35297(x35297, x35197, x35175);
  nand n35299(x35299, x35297, x35298);
  nand n35300(x35300, x35197, x35177);
  nand n35302(x35302, x35202, x35180);
  nand n35304(x35304, x35302, x35303);
  nand n35305(x35305, x35202, x35182);
  nand n35307(x35307, x35207, x35185);
  nand n35309(x35309, x35307, x35308);
  nand n35310(x35310, x35207, x35187);
  nand n35312(x35312, x35212, x35190);
  nand n35314(x35314, x35312, x35313);
  nand n35315(x35315, x35212, x35192);
  nand n35317(x35317, x35217, x35195);
  nand n35319(x35319, x35317, x35318);
  nand n35320(x35320, x35217, x35197);
  nand n35322(x35322, x35222, x35200);
  nand n35324(x35324, x35322, x35323);
  nand n35325(x35325, x35222, x35202);
  nand n35327(x35327, x35227, x35205);
  nand n35329(x35329, x35327, x35328);
  nand n35330(x35330, x35227, x35207);
  nand n35332(x35332, x35232, x35210);
  nand n35334(x35334, x35332, x35333);
  nand n35335(x35335, x35232, x35212);
  nand n35337(x35337, x35237, x35215);
  nand n35339(x35339, x35337, x35338);
  nand n35340(x35340, x35237, x35217);
  nand n35342(x35342, x35242, x35220);
  nand n35344(x35344, x35342, x35343);
  nand n35345(x35345, x35242, x35222);
  nand n35347(x35347, x35247, x35225);
  nand n35349(x35349, x35347, x35348);
  nand n35350(x35350, x35247, x35227);
  nand n35352(x35352, x35252, x35230);
  nand n35354(x35354, x35352, x35353);
  nand n35355(x35355, x35252, x35232);
  nand n35357(x35357, x35257, x35235);
  nand n35359(x35359, x35357, x35358);
  nand n35360(x35360, x35257, x35237);
  nand n35362(x35362, x35262, x35240);
  nand n35364(x35364, x35362, x35363);
  nand n35365(x35365, x35262, x35242);
  nand n35367(x35367, x35267, x35245);
  nand n35369(x35369, x35367, x35368);
  nand n35370(x35370, x35267, x35247);
  nand n35372(x35372, x35272, x35250);
  nand n35374(x35374, x35372, x35373);
  nand n35375(x35375, x35272, x35252);
  nand n35377(x35377, x35277, x35255);
  nand n35379(x35379, x35377, x35378);
  nand n35380(x35380, x35277, x35257);
  nand n35382(x35382, x35282, x35260);
  nand n35384(x35384, x35382, x35383);
  nand n35385(x35385, x35282, x35262);
  nand n35391(x35391, x35301, x35043);
  nand n35393(x35393, x35391, x35392);
  nand n35394(x35394, x35306, x35069);
  nand n35396(x35396, x35394, x35395);
  nand n35397(x35397, x35311, x35169);
  nand n35399(x35399, x35397, x35398);
  nand n35400(x35400, x35316, x35172);
  nand n35402(x35402, x35400, x35401);
  nand n35403(x35403, x35321, x35287);
  nand n35405(x35405, x35403, x35404);
  nand n35406(x35406, x35326, x35290);
  nand n35408(x35408, x35406, x35407);
  nand n35409(x35409, x35331, x35293);
  nand n35411(x35411, x35409, x35410);
  nand n35412(x35412, x35336, x35296);
  nand n35414(x35414, x35412, x35413);
  nand n35415(x35415, x35341, x35299);
  nand n35417(x35417, x35415, x35416);
  nand n35418(x35418, x35341, x35301);
  nand n35420(x35420, x35346, x35304);
  nand n35422(x35422, x35420, x35421);
  nand n35423(x35423, x35346, x35306);
  nand n35425(x35425, x35351, x35309);
  nand n35427(x35427, x35425, x35426);
  nand n35428(x35428, x35351, x35311);
  nand n35430(x35430, x35356, x35314);
  nand n35432(x35432, x35430, x35431);
  nand n35433(x35433, x35356, x35316);
  nand n35435(x35435, x35361, x35319);
  nand n35437(x35437, x35435, x35436);
  nand n35438(x35438, x35361, x35321);
  nand n35440(x35440, x35366, x35324);
  nand n35442(x35442, x35440, x35441);
  nand n35443(x35443, x35366, x35326);
  nand n35445(x35445, x35371, x35329);
  nand n35447(x35447, x35445, x35446);
  nand n35448(x35448, x35371, x35331);
  nand n35450(x35450, x35376, x35334);
  nand n35452(x35452, x35450, x35451);
  nand n35453(x35453, x35376, x35336);
  nand n35455(x35455, x35381, x35339);
  nand n35457(x35457, x35455, x35456);
  nand n35458(x35458, x35381, x35341);
  nand n35460(x35460, x35386, x35344);
  nand n35462(x35462, x35460, x35461);
  nand n35463(x35463, x35386, x35346);
  nand n35471(x35471, x35419, x35043);
  nand n35473(x35473, x35471, x35472);
  nand n35474(x35474, x35424, x35069);
  nand n35476(x35476, x35474, x35475);
  nand n35477(x35477, x35429, x35169);
  nand n35479(x35479, x35477, x35478);
  nand n35480(x35480, x35434, x35172);
  nand n35482(x35482, x35480, x35481);
  nand n35483(x35483, x35439, x35287);
  nand n35485(x35485, x35483, x35484);
  nand n35486(x35486, x35444, x35290);
  nand n35488(x35488, x35486, x35487);
  nand n35489(x35489, x35449, x35293);
  nand n35491(x35491, x35489, x35490);
  nand n35492(x35492, x35454, x35296);
  nand n35494(x35494, x35492, x35493);
  nand n35495(x35495, x35459, x35393);
  nand n35497(x35497, x35495, x35496);
  nand n35498(x35498, x35464, x35396);
  nand n35500(x35500, x35498, x35499);
  nand n35501(x35501, x34917, x34911);
  nand n35502(x35502, x35501, x35068);
  nand n35504(x35504, x34922, x35069);
  nand n35505(x35505, x34921, x35166);
  nand n35506(x35506, x35505, x35504);
  nand n35508(x35508, x34927, x35169);
  nand n35509(x35509, x34926, x35283);
  nand n35510(x35510, x35509, x35508);
  nand n35512(x35512, x34932, x35172);
  nand n35513(x35513, x34931, x35284);
  nand n35514(x35514, x35513, x35512);
  nand n35516(x35516, x34937, x35287);
  nand n35517(x35517, x34936, x35387);
  nand n35518(x35518, x35517, x35516);
  nand n35520(x35520, x34942, x35290);
  nand n35521(x35521, x34941, x35388);
  nand n35522(x35522, x35521, x35520);
  nand n35524(x35524, x34947, x35293);
  nand n35525(x35525, x34946, x35389);
  nand n35526(x35526, x35525, x35524);
  nand n35528(x35528, x34952, x35296);
  nand n35529(x35529, x34951, x35390);
  nand n35530(x35530, x35529, x35528);
  nand n35532(x35532, x34957, x35393);
  nand n35534(x35534, x34956, x35533);
  nand n35535(x35535, x35534, x35532);
  nand n35537(x35537, x34962, x35396);
  nand n35539(x35539, x34961, x35538);
  nand n35540(x35540, x35539, x35537);
  nand n35542(x35542, x34967, x35399);
  nand n35543(x35543, x34966, x35465);
  nand n35544(x35544, x35543, x35542);
  nand n35546(x35546, x34972, x35402);
  nand n35547(x35547, x34971, x35466);
  nand n35548(x35548, x35547, x35546);
  nand n35550(x35550, x34977, x35405);
  nand n35551(x35551, x34976, x35467);
  nand n35552(x35552, x35551, x35550);
  nand n35554(x35554, x34982, x35408);
  nand n35555(x35555, x34981, x35468);
  nand n35556(x35556, x35555, x35554);
  nand n35558(x35558, x34987, x35411);
  nand n35559(x35559, x34986, x35469);
  nand n35560(x35560, x35559, x35558);
  nand n35562(x35562, x34992, x35414);
  nand n35563(x35563, x34991, x35470);
  nand n35564(x35564, x35563, x35562);
  nand n35566(x35566, x34997, x35473);
  nand n35568(x35568, x34996, x35567);
  nand n35569(x35569, x35568, x35566);
  nand n35571(x35571, x35002, x35476);
  nand n35573(x35573, x35001, x35572);
  nand n35574(x35574, x35573, x35571);
  nand n35576(x35576, x35007, x35479);
  nand n35578(x35578, x35006, x35577);
  nand n35579(x35579, x35578, x35576);
  nand n35581(x35581, x35012, x35482);
  nand n35583(x35583, x35011, x35582);
  nand n35584(x35584, x35583, x35581);
  nand n35586(x35586, x35017, x35485);
  nand n35588(x35588, x35016, x35587);
  nand n35589(x35589, x35588, x35586);
  nand n35591(x35591, x35022, x35488);
  nand n35593(x35593, x35021, x35592);
  nand n35594(x35594, x35593, x35591);
  nand n35596(x35596, x35027, x35491);
  nand n35598(x35598, x35026, x35597);
  nand n35599(x35599, x35598, x35596);
  nand n35601(x35601, x35032, x35494);
  nand n35603(x35603, x35031, x35602);
  nand n35604(x35604, x35603, x35601);
  nand n35606(x35606, x35037, x35497);
  nand n35608(x35608, x35036, x35607);
  nand n35609(x35609, x35608, x35606);
  nand n35611(x35611, x35042, x35500);
  nand n35613(x35613, x35041, x35612);
  nand n35614(x35614, x35613, x35611);
  nand n35616(x35616, x28080, x28074);
  nand n35618(x35618, x28086, x28080);
  nand n35620(x35620, x28092, x28086);
  nand n35622(x35622, x28098, x28092);
  nand n35624(x35624, x28104, x28098);
  nand n35626(x35626, x28110, x28104);
  nand n35628(x35628, x28116, x28110);
  nand n35630(x35630, x28122, x28116);
  nand n35632(x35632, x28128, x28122);
  nand n35634(x35634, x28134, x28128);
  nand n35636(x35636, x28140, x28134);
  nand n35638(x35638, x28146, x28140);
  nand n35640(x35640, x28152, x28146);
  nand n35642(x35642, x28158, x28152);
  nand n35644(x35644, x28164, x28158);
  nand n35646(x35646, x28170, x28164);
  nand n35648(x35648, x28176, x28170);
  nand n35650(x35650, x28182, x28176);
  nand n35652(x35652, x28188, x28182);
  nand n35654(x35654, x28194, x28188);
  nand n35656(x35656, x28200, x28194);
  nand n35658(x35658, x28206, x28200);
  nand n35660(x35660, x28212, x28206);
  nand n35662(x35662, x28218, x28212);
  nand n35664(x35664, x28224, x28218);
  nand n35666(x35666, x28230, x28224);
  nand n35668(x35668, x28236, x28230);
  nand n35670(x35670, x28242, x28236);
  nand n35672(x35672, x28248, x28242);
  nand n35674(x35674, x28254, x28248);
  nand n35676(x35676, x35619, x28074);
  nand n35677(x35677, x35621, x35617);
  nand n35679(x35679, x35623, x35619);
  nand n35681(x35681, x35625, x35621);
  nand n35683(x35683, x35627, x35623);
  nand n35685(x35685, x35629, x35625);
  nand n35687(x35687, x35631, x35627);
  nand n35689(x35689, x35633, x35629);
  nand n35691(x35691, x35635, x35631);
  nand n35693(x35693, x35637, x35633);
  nand n35695(x35695, x35639, x35635);
  nand n35697(x35697, x35641, x35637);
  nand n35699(x35699, x35643, x35639);
  nand n35701(x35701, x35645, x35641);
  nand n35703(x35703, x35647, x35643);
  nand n35705(x35705, x35649, x35645);
  nand n35707(x35707, x35651, x35647);
  nand n35709(x35709, x35653, x35649);
  nand n35711(x35711, x35655, x35651);
  nand n35713(x35713, x35657, x35653);
  nand n35715(x35715, x35659, x35655);
  nand n35717(x35717, x35661, x35657);
  nand n35719(x35719, x35663, x35659);
  nand n35721(x35721, x35665, x35661);
  nand n35723(x35723, x35667, x35663);
  nand n35725(x35725, x35669, x35665);
  nand n35727(x35727, x35671, x35667);
  nand n35729(x35729, x35673, x35669);
  nand n35731(x35731, x35675, x35671);
  nand n35733(x35733, x35680, x28074);
  nand n35734(x35734, x35682, x35617);
  nand n35735(x35735, x35684, x84562);
  nand n35736(x35736, x35686, x35678);
  nand n35738(x35738, x35688, x35680);
  nand n35740(x35740, x35690, x35682);
  nand n35742(x35742, x35692, x35684);
  nand n35744(x35744, x35694, x35686);
  nand n35746(x35746, x35696, x35688);
  nand n35748(x35748, x35698, x35690);
  nand n35750(x35750, x35700, x35692);
  nand n35752(x35752, x35702, x35694);
  nand n35754(x35754, x35704, x35696);
  nand n35756(x35756, x35706, x35698);
  nand n35758(x35758, x35708, x35700);
  nand n35760(x35760, x35710, x35702);
  nand n35762(x35762, x35712, x35704);
  nand n35764(x35764, x35714, x35706);
  nand n35766(x35766, x35716, x35708);
  nand n35768(x35768, x35718, x35710);
  nand n35770(x35770, x35720, x35712);
  nand n35772(x35772, x35722, x35714);
  nand n35774(x35774, x35724, x35716);
  nand n35776(x35776, x35726, x35718);
  nand n35778(x35778, x35728, x35720);
  nand n35780(x35780, x35730, x35722);
  nand n35782(x35782, x35732, x35724);
  nand n35784(x35784, x35739, x28074);
  nand n35785(x35785, x35741, x35617);
  nand n35786(x35786, x35743, x84562);
  nand n35787(x35787, x35745, x35678);
  nand n35788(x35788, x35747, x84563);
  nand n35789(x35789, x35749, x84564);
  nand n35790(x35790, x35751, x84565);
  nand n35791(x35791, x35753, x35737);
  nand n35792(x35792, x35755, x35739);
  nand n35794(x35794, x35757, x35741);
  nand n35796(x35796, x35759, x35743);
  nand n35798(x35798, x35761, x35745);
  nand n35800(x35800, x35763, x35747);
  nand n35802(x35802, x35765, x35749);
  nand n35804(x35804, x35767, x35751);
  nand n35806(x35806, x35769, x35753);
  nand n35808(x35808, x35771, x35755);
  nand n35810(x35810, x35773, x35757);
  nand n35812(x35812, x35775, x35759);
  nand n35814(x35814, x35777, x35761);
  nand n35816(x35816, x35779, x35763);
  nand n35818(x35818, x35781, x35765);
  nand n35820(x35820, x35783, x35767);
  nand n35822(x35822, x35793, x28074);
  nand n35823(x35823, x35795, x35617);
  nand n35824(x35824, x35797, x84562);
  nand n35825(x35825, x35799, x35678);
  nand n35826(x35826, x35801, x84563);
  nand n35827(x35827, x35803, x84564);
  nand n35828(x35828, x35805, x84565);
  nand n35829(x35829, x35807, x35737);
  nand n35830(x35830, x35809, x84566);
  nand n35831(x35831, x35811, x84567);
  nand n35832(x35832, x35813, x84568);
  nand n35833(x35833, x35815, x84569);
  nand n35834(x35834, x35817, x84570);
  nand n35835(x35835, x35819, x84571);
  nand n35836(x35836, x35821, x84572);
  nand n35837(x35837, x72542, x72537);
  nand n35838(x35838, x35837, x35616);
  nand n35840(x35840, x28086, x35617);
  nand n35841(x35841, x72547, x35616);
  nand n35842(x35842, x35841, x35840);
  nand n35844(x35844, x28092, x84562);
  nand n35845(x35845, x72552, x35676);
  nand n35846(x35846, x35845, x35844);
  nand n35848(x35848, x28098, x35678);
  nand n35849(x35849, x72557, x35677);
  nand n35850(x35850, x35849, x35848);
  nand n35852(x35852, x28104, x84563);
  nand n35853(x35853, x72562, x35733);
  nand n35854(x35854, x35853, x35852);
  nand n35856(x35856, x28110, x84564);
  nand n35857(x35857, x72567, x35734);
  nand n35858(x35858, x35857, x35856);
  nand n35860(x35860, x28116, x84565);
  nand n35861(x35861, x72572, x35735);
  nand n35862(x35862, x35861, x35860);
  nand n35864(x35864, x28122, x35737);
  nand n35865(x35865, x72577, x35736);
  nand n35866(x35866, x35865, x35864);
  nand n35868(x35868, x28128, x84566);
  nand n35869(x35869, x72582, x35784);
  nand n35870(x35870, x35869, x35868);
  nand n35872(x35872, x28134, x84567);
  nand n35873(x35873, x72587, x35785);
  nand n35874(x35874, x35873, x35872);
  nand n35876(x35876, x28140, x84568);
  nand n35877(x35877, x72592, x35786);
  nand n35878(x35878, x35877, x35876);
  nand n35880(x35880, x28146, x84569);
  nand n35881(x35881, x72597, x35787);
  nand n35882(x35882, x35881, x35880);
  nand n35884(x35884, x28152, x84570);
  nand n35885(x35885, x72602, x35788);
  nand n35886(x35886, x35885, x35884);
  nand n35888(x35888, x28158, x84571);
  nand n35889(x35889, x72607, x35789);
  nand n35890(x35890, x35889, x35888);
  nand n35892(x35892, x28164, x84572);
  nand n35893(x35893, x72612, x35790);
  nand n35894(x35894, x35893, x35892);
  nand n35896(x35896, x28170, x84573);
  nand n35897(x35897, x72617, x35791);
  nand n35898(x35898, x35897, x35896);
  nand n35900(x35900, x28176, x84574);
  nand n35901(x35901, x72622, x35822);
  nand n35902(x35902, x35901, x35900);
  nand n35904(x35904, x28182, x84575);
  nand n35905(x35905, x72627, x35823);
  nand n35906(x35906, x35905, x35904);
  nand n35908(x35908, x28188, x84576);
  nand n35909(x35909, x72632, x35824);
  nand n35910(x35910, x35909, x35908);
  nand n35912(x35912, x28194, x84577);
  nand n35913(x35913, x72637, x35825);
  nand n35914(x35914, x35913, x35912);
  nand n35916(x35916, x28200, x84578);
  nand n35917(x35917, x72642, x35826);
  nand n35918(x35918, x35917, x35916);
  nand n35920(x35920, x28206, x84579);
  nand n35921(x35921, x72647, x35827);
  nand n35922(x35922, x35921, x35920);
  nand n35924(x35924, x28212, x84580);
  nand n35925(x35925, x72652, x35828);
  nand n35926(x35926, x35925, x35924);
  nand n35928(x35928, x28218, x84581);
  nand n35929(x35929, x72657, x35829);
  nand n35930(x35930, x35929, x35928);
  nand n35932(x35932, x28224, x84582);
  nand n35933(x35933, x72662, x35830);
  nand n35934(x35934, x35933, x35932);
  nand n35936(x35936, x28230, x84583);
  nand n35937(x35937, x72667, x35831);
  nand n35938(x35938, x35937, x35936);
  nand n35940(x35940, x28236, x84584);
  nand n35941(x35941, x72672, x35832);
  nand n35942(x35942, x35941, x35940);
  nand n35944(x35944, x28242, x84585);
  nand n35945(x35945, x72677, x35833);
  nand n35946(x35946, x35945, x35944);
  nand n35948(x35948, x28248, x84586);
  nand n35949(x35949, x72682, x35834);
  nand n35950(x35950, x35949, x35948);
  nand n35952(x35952, x28254, x84587);
  nand n35953(x35953, x72687, x35835);
  nand n35954(x35954, x35953, x35952);
  nand n35956(x35956, x28260, x84588);
  nand n35957(x35957, x72692, x35836);
  nand n35958(x35958, x35957, x35956);
  nand n35961(x35961, x72617, x27913);
  nand n35963(x35963, x72622, x27915);
  nand n35965(x35965, x72627, x27917);
  nand n35967(x35967, x72632, x27919);
  nand n35969(x35969, x72637, x27921);
  nand n35971(x35971, x72642, x27923);
  nand n35973(x35973, x72647, x27925);
  nand n35975(x35975, x72652, x27927);
  nand n35977(x35977, x72657, x27929);
  nand n35979(x35979, x72662, x27931);
  nand n35981(x35981, x72667, x27933);
  nand n35983(x35983, x72672, x27935);
  nand n35985(x35985, x72677, x27937);
  nand n35987(x35987, x72682, x27939);
  nand n35989(x35989, x72687, x27941);
  nand n35991(x35991, x72692, x27943);
  nand n35993(x35993, x28074, x27944);
  nand n35994(x35994, x28080, x27945);
  nand n35995(x35995, x28086, x27946);
  nand n35996(x35996, x28092, x27947);
  nand n35997(x35997, x28098, x27948);
  nand n35998(x35998, x28104, x27949);
  nand n35999(x35999, x28110, x27950);
  nand n36000(x36000, x28116, x27951);
  nand n36001(x36001, x28122, x27952);
  nand n36002(x36002, x28128, x27953);
  nand n36003(x36003, x28134, x27954);
  nand n36004(x36004, x28140, x27955);
  nand n36005(x36005, x28146, x27956);
  nand n36006(x36006, x28152, x27957);
  nand n36007(x36007, x28158, x27958);
  nand n36008(x36008, x28164, x27959);
  nand n36009(x36009, x28170, x27960);
  nand n36010(x36010, x28176, x27961);
  nand n36011(x36011, x28182, x27962);
  nand n36012(x36012, x28188, x27963);
  nand n36013(x36013, x28194, x27964);
  nand n36014(x36014, x28200, x27965);
  nand n36015(x36015, x28206, x27966);
  nand n36016(x36016, x28212, x27967);
  nand n36017(x36017, x28218, x27968);
  nand n36018(x36018, x28224, x27969);
  nand n36019(x36019, x28230, x27970);
  nand n36020(x36020, x28236, x27971);
  nand n36021(x36021, x28242, x27972);
  nand n36022(x36022, x28248, x27973);
  nand n36023(x36023, x28254, x27974);
  nand n36024(x36024, x28260, x27975);
  nand n36025(x36025, x35993, x29004);
  nand n36027(x36027, x35994, x29011);
  nand n36029(x36029, x35995, x29026);
  nand n36031(x36031, x35996, x29050);
  nand n36033(x36033, x35997, x29081);
  nand n36035(x36035, x35998, x29120);
  nand n36037(x36037, x35999, x29168);
  nand n36039(x36039, x36000, x29223);
  nand n36041(x36041, x36001, x29286);
  nand n36043(x36043, x36002, x29358);
  nand n36045(x36045, x36003, x29437);
  nand n36047(x36047, x36004, x29524);
  nand n36049(x36049, x36005, x29620);
  nand n36051(x36051, x36006, x29723);
  nand n36053(x36053, x36007, x29834);
  nand n36055(x36055, x36008, x29954);
  nand n36057(x36057, x36009, x35961);
  nand n36059(x36059, x36010, x35963);
  nand n36061(x36061, x36011, x35965);
  nand n36063(x36063, x36012, x35967);
  nand n36065(x36065, x36013, x35969);
  nand n36067(x36067, x36014, x35971);
  nand n36069(x36069, x36015, x35973);
  nand n36071(x36071, x36016, x35975);
  nand n36073(x36073, x36017, x35977);
  nand n36075(x36075, x36018, x35979);
  nand n36077(x36077, x36019, x35981);
  nand n36079(x36079, x36020, x35983);
  nand n36081(x36081, x36021, x35985);
  nand n36083(x36083, x36022, x35987);
  nand n36085(x36085, x36023, x35989);
  nand n36087(x36087, x36024, x35991);
  nand n36089(x36089, x27944, x72537);
  nand n36090(x36090, x27944, x72542);
  nand n36091(x36091, x36090, x29004);
  nand n36092(x36092, x27944, x72547);
  nand n36093(x36093, x36092, x29005);
  nand n36094(x36094, x27944, x72552);
  nand n36095(x36095, x36094, x29009);
  nand n36096(x36096, x27944, x72557);
  nand n36097(x36097, x36096, x29015);
  nand n36098(x36098, x27944, x72562);
  nand n36099(x36099, x36098, x29022);
  nand n36100(x36100, x27944, x72567);
  nand n36101(x36101, x36100, x29032);
  nand n36102(x36102, x27944, x72572);
  nand n36103(x36103, x36102, x29044);
  nand n36104(x36104, x27944, x72577);
  nand n36105(x36105, x36104, x29057);
  nand n36106(x36106, x27944, x72582);
  nand n36107(x36107, x36106, x29073);
  nand n36108(x36108, x27944, x72587);
  nand n36109(x36109, x36108, x29091);
  nand n36110(x36110, x27944, x72592);
  nand n36111(x36111, x36110, x29110);
  nand n36112(x36112, x27944, x72597);
  nand n36113(x36113, x36112, x29132);
  nand n36114(x36114, x27944, x72602);
  nand n36115(x36115, x36114, x29156);
  nand n36116(x36116, x27944, x72607);
  nand n36117(x36117, x36116, x29181);
  nand n36118(x36118, x27944, x72612);
  nand n36119(x36119, x36118, x29209);
  nand n36120(x36120, x27944, x72617);
  nand n36121(x36121, x36120, x29239);
  nand n36122(x36122, x27944, x72622);
  nand n36123(x36123, x36122, x29270);
  nand n36124(x36124, x27944, x72627);
  nand n36125(x36125, x36124, x29304);
  nand n36126(x36126, x27944, x72632);
  nand n36127(x36127, x36126, x29340);
  nand n36128(x36128, x27944, x72637);
  nand n36129(x36129, x36128, x29377);
  nand n36130(x36130, x27944, x72642);
  nand n36131(x36131, x36130, x29417);
  nand n36132(x36132, x27944, x72647);
  nand n36133(x36133, x36132, x29459);
  nand n36134(x36134, x27944, x72652);
  nand n36135(x36135, x36134, x29502);
  nand n36136(x36136, x27944, x72657);
  nand n36137(x36137, x36136, x29548);
  nand n36138(x36138, x27944, x72662);
  nand n36139(x36139, x36138, x29596);
  nand n36140(x36140, x27944, x72667);
  nand n36141(x36141, x36140, x29645);
  nand n36142(x36142, x27944, x72672);
  nand n36143(x36143, x36142, x29697);
  nand n36144(x36144, x27944, x72677);
  nand n36145(x36145, x36144, x29751);
  nand n36146(x36146, x27944, x72682);
  nand n36147(x36147, x36146, x29806);
  nand n36148(x36148, x27944, x72687);
  nand n36149(x36149, x36148, x29864);
  nand n36150(x36150, x27944, x72692);
  nand n36151(x36151, x36150, x29924);
  nand n36152(x36152, x27945, x84589);
  nand n36153(x36153, x27945, x36091);
  nand n36154(x36154, x27883, x84589);
  nand n36155(x36155, x27945, x36093);
  nand n36156(x36156, x36155, x36154);
  nand n36157(x36157, x27883, x36091);
  nand n36158(x36158, x27945, x36095);
  nand n36159(x36159, x36158, x36157);
  nand n36160(x36160, x27883, x36093);
  nand n36161(x36161, x27945, x36097);
  nand n36162(x36162, x36161, x36160);
  nand n36163(x36163, x27883, x36095);
  nand n36164(x36164, x27945, x36099);
  nand n36165(x36165, x36164, x36163);
  nand n36166(x36166, x27883, x36097);
  nand n36167(x36167, x27945, x36101);
  nand n36168(x36168, x36167, x36166);
  nand n36169(x36169, x27883, x36099);
  nand n36170(x36170, x27945, x36103);
  nand n36171(x36171, x36170, x36169);
  nand n36172(x36172, x27883, x36101);
  nand n36173(x36173, x27945, x36105);
  nand n36174(x36174, x36173, x36172);
  nand n36175(x36175, x27883, x36103);
  nand n36176(x36176, x27945, x36107);
  nand n36177(x36177, x36176, x36175);
  nand n36178(x36178, x27883, x36105);
  nand n36179(x36179, x27945, x36109);
  nand n36180(x36180, x36179, x36178);
  nand n36181(x36181, x27883, x36107);
  nand n36182(x36182, x27945, x36111);
  nand n36183(x36183, x36182, x36181);
  nand n36184(x36184, x27883, x36109);
  nand n36185(x36185, x27945, x36113);
  nand n36186(x36186, x36185, x36184);
  nand n36187(x36187, x27883, x36111);
  nand n36188(x36188, x27945, x36115);
  nand n36189(x36189, x36188, x36187);
  nand n36190(x36190, x27883, x36113);
  nand n36191(x36191, x27945, x36117);
  nand n36192(x36192, x36191, x36190);
  nand n36193(x36193, x27883, x36115);
  nand n36194(x36194, x27945, x36119);
  nand n36195(x36195, x36194, x36193);
  nand n36196(x36196, x27883, x36117);
  nand n36197(x36197, x27945, x36121);
  nand n36198(x36198, x36197, x36196);
  nand n36199(x36199, x27883, x36119);
  nand n36200(x36200, x27945, x36123);
  nand n36201(x36201, x36200, x36199);
  nand n36202(x36202, x27883, x36121);
  nand n36203(x36203, x27945, x36125);
  nand n36204(x36204, x36203, x36202);
  nand n36205(x36205, x27883, x36123);
  nand n36206(x36206, x27945, x36127);
  nand n36207(x36207, x36206, x36205);
  nand n36208(x36208, x27883, x36125);
  nand n36209(x36209, x27945, x36129);
  nand n36210(x36210, x36209, x36208);
  nand n36211(x36211, x27883, x36127);
  nand n36212(x36212, x27945, x36131);
  nand n36213(x36213, x36212, x36211);
  nand n36214(x36214, x27883, x36129);
  nand n36215(x36215, x27945, x36133);
  nand n36216(x36216, x36215, x36214);
  nand n36217(x36217, x27883, x36131);
  nand n36218(x36218, x27945, x36135);
  nand n36219(x36219, x36218, x36217);
  nand n36220(x36220, x27883, x36133);
  nand n36221(x36221, x27945, x36137);
  nand n36222(x36222, x36221, x36220);
  nand n36223(x36223, x27883, x36135);
  nand n36224(x36224, x27945, x36139);
  nand n36225(x36225, x36224, x36223);
  nand n36226(x36226, x27883, x36137);
  nand n36227(x36227, x27945, x36141);
  nand n36228(x36228, x36227, x36226);
  nand n36229(x36229, x27883, x36139);
  nand n36230(x36230, x27945, x36143);
  nand n36231(x36231, x36230, x36229);
  nand n36232(x36232, x27883, x36141);
  nand n36233(x36233, x27945, x36145);
  nand n36234(x36234, x36233, x36232);
  nand n36235(x36235, x27883, x36143);
  nand n36236(x36236, x27945, x36147);
  nand n36237(x36237, x36236, x36235);
  nand n36238(x36238, x27883, x36145);
  nand n36239(x36239, x27945, x36149);
  nand n36240(x36240, x36239, x36238);
  nand n36241(x36241, x27883, x36147);
  nand n36242(x36242, x27945, x36151);
  nand n36243(x36243, x36242, x36241);
  nand n36244(x36244, x27946, x84590);
  nand n36245(x36245, x27946, x84591);
  nand n36246(x36246, x27946, x36156);
  nand n36247(x36247, x27946, x36159);
  nand n36248(x36248, x27885, x84590);
  nand n36249(x36249, x27946, x36162);
  nand n36250(x36250, x36249, x36248);
  nand n36251(x36251, x27885, x84591);
  nand n36252(x36252, x27946, x36165);
  nand n36253(x36253, x36252, x36251);
  nand n36254(x36254, x27885, x36156);
  nand n36255(x36255, x27946, x36168);
  nand n36256(x36256, x36255, x36254);
  nand n36257(x36257, x27885, x36159);
  nand n36258(x36258, x27946, x36171);
  nand n36259(x36259, x36258, x36257);
  nand n36260(x36260, x27885, x36162);
  nand n36261(x36261, x27946, x36174);
  nand n36262(x36262, x36261, x36260);
  nand n36263(x36263, x27885, x36165);
  nand n36264(x36264, x27946, x36177);
  nand n36265(x36265, x36264, x36263);
  nand n36266(x36266, x27885, x36168);
  nand n36267(x36267, x27946, x36180);
  nand n36268(x36268, x36267, x36266);
  nand n36269(x36269, x27885, x36171);
  nand n36270(x36270, x27946, x36183);
  nand n36271(x36271, x36270, x36269);
  nand n36272(x36272, x27885, x36174);
  nand n36273(x36273, x27946, x36186);
  nand n36274(x36274, x36273, x36272);
  nand n36275(x36275, x27885, x36177);
  nand n36276(x36276, x27946, x36189);
  nand n36277(x36277, x36276, x36275);
  nand n36278(x36278, x27885, x36180);
  nand n36279(x36279, x27946, x36192);
  nand n36280(x36280, x36279, x36278);
  nand n36281(x36281, x27885, x36183);
  nand n36282(x36282, x27946, x36195);
  nand n36283(x36283, x36282, x36281);
  nand n36284(x36284, x27885, x36186);
  nand n36285(x36285, x27946, x36198);
  nand n36286(x36286, x36285, x36284);
  nand n36287(x36287, x27885, x36189);
  nand n36288(x36288, x27946, x36201);
  nand n36289(x36289, x36288, x36287);
  nand n36290(x36290, x27885, x36192);
  nand n36291(x36291, x27946, x36204);
  nand n36292(x36292, x36291, x36290);
  nand n36293(x36293, x27885, x36195);
  nand n36294(x36294, x27946, x36207);
  nand n36295(x36295, x36294, x36293);
  nand n36296(x36296, x27885, x36198);
  nand n36297(x36297, x27946, x36210);
  nand n36298(x36298, x36297, x36296);
  nand n36299(x36299, x27885, x36201);
  nand n36300(x36300, x27946, x36213);
  nand n36301(x36301, x36300, x36299);
  nand n36302(x36302, x27885, x36204);
  nand n36303(x36303, x27946, x36216);
  nand n36304(x36304, x36303, x36302);
  nand n36305(x36305, x27885, x36207);
  nand n36306(x36306, x27946, x36219);
  nand n36307(x36307, x36306, x36305);
  nand n36308(x36308, x27885, x36210);
  nand n36309(x36309, x27946, x36222);
  nand n36310(x36310, x36309, x36308);
  nand n36311(x36311, x27885, x36213);
  nand n36312(x36312, x27946, x36225);
  nand n36313(x36313, x36312, x36311);
  nand n36314(x36314, x27885, x36216);
  nand n36315(x36315, x27946, x36228);
  nand n36316(x36316, x36315, x36314);
  nand n36317(x36317, x27885, x36219);
  nand n36318(x36318, x27946, x36231);
  nand n36319(x36319, x36318, x36317);
  nand n36320(x36320, x27885, x36222);
  nand n36321(x36321, x27946, x36234);
  nand n36322(x36322, x36321, x36320);
  nand n36323(x36323, x27885, x36225);
  nand n36324(x36324, x27946, x36237);
  nand n36325(x36325, x36324, x36323);
  nand n36326(x36326, x27885, x36228);
  nand n36327(x36327, x27946, x36240);
  nand n36328(x36328, x36327, x36326);
  nand n36329(x36329, x27885, x36231);
  nand n36330(x36330, x27946, x36243);
  nand n36331(x36331, x36330, x36329);
  nand n36332(x36332, x27947, x84592);
  nand n36333(x36333, x27947, x84593);
  nand n36334(x36334, x27947, x84594);
  nand n36335(x36335, x27947, x84595);
  nand n36336(x36336, x27947, x36250);
  nand n36337(x36337, x27947, x36253);
  nand n36338(x36338, x27947, x36256);
  nand n36339(x36339, x27947, x36259);
  nand n36340(x36340, x27887, x84592);
  nand n36341(x36341, x27947, x36262);
  nand n36342(x36342, x36341, x36340);
  nand n36343(x36343, x27887, x84593);
  nand n36344(x36344, x27947, x36265);
  nand n36345(x36345, x36344, x36343);
  nand n36346(x36346, x27887, x84594);
  nand n36347(x36347, x27947, x36268);
  nand n36348(x36348, x36347, x36346);
  nand n36349(x36349, x27887, x84595);
  nand n36350(x36350, x27947, x36271);
  nand n36351(x36351, x36350, x36349);
  nand n36352(x36352, x27887, x36250);
  nand n36353(x36353, x27947, x36274);
  nand n36354(x36354, x36353, x36352);
  nand n36355(x36355, x27887, x36253);
  nand n36356(x36356, x27947, x36277);
  nand n36357(x36357, x36356, x36355);
  nand n36358(x36358, x27887, x36256);
  nand n36359(x36359, x27947, x36280);
  nand n36360(x36360, x36359, x36358);
  nand n36361(x36361, x27887, x36259);
  nand n36362(x36362, x27947, x36283);
  nand n36363(x36363, x36362, x36361);
  nand n36364(x36364, x27887, x36262);
  nand n36365(x36365, x27947, x36286);
  nand n36366(x36366, x36365, x36364);
  nand n36367(x36367, x27887, x36265);
  nand n36368(x36368, x27947, x36289);
  nand n36369(x36369, x36368, x36367);
  nand n36370(x36370, x27887, x36268);
  nand n36371(x36371, x27947, x36292);
  nand n36372(x36372, x36371, x36370);
  nand n36373(x36373, x27887, x36271);
  nand n36374(x36374, x27947, x36295);
  nand n36375(x36375, x36374, x36373);
  nand n36376(x36376, x27887, x36274);
  nand n36377(x36377, x27947, x36298);
  nand n36378(x36378, x36377, x36376);
  nand n36379(x36379, x27887, x36277);
  nand n36380(x36380, x27947, x36301);
  nand n36381(x36381, x36380, x36379);
  nand n36382(x36382, x27887, x36280);
  nand n36383(x36383, x27947, x36304);
  nand n36384(x36384, x36383, x36382);
  nand n36385(x36385, x27887, x36283);
  nand n36386(x36386, x27947, x36307);
  nand n36387(x36387, x36386, x36385);
  nand n36388(x36388, x27887, x36286);
  nand n36389(x36389, x27947, x36310);
  nand n36390(x36390, x36389, x36388);
  nand n36391(x36391, x27887, x36289);
  nand n36392(x36392, x27947, x36313);
  nand n36393(x36393, x36392, x36391);
  nand n36394(x36394, x27887, x36292);
  nand n36395(x36395, x27947, x36316);
  nand n36396(x36396, x36395, x36394);
  nand n36397(x36397, x27887, x36295);
  nand n36398(x36398, x27947, x36319);
  nand n36399(x36399, x36398, x36397);
  nand n36400(x36400, x27887, x36298);
  nand n36401(x36401, x27947, x36322);
  nand n36402(x36402, x36401, x36400);
  nand n36403(x36403, x27887, x36301);
  nand n36404(x36404, x27947, x36325);
  nand n36405(x36405, x36404, x36403);
  nand n36406(x36406, x27887, x36304);
  nand n36407(x36407, x27947, x36328);
  nand n36408(x36408, x36407, x36406);
  nand n36409(x36409, x27887, x36307);
  nand n36410(x36410, x27947, x36331);
  nand n36411(x36411, x36410, x36409);
  nand n36412(x36412, x27948, x84596);
  nand n36413(x36413, x27948, x84597);
  nand n36414(x36414, x27948, x84598);
  nand n36415(x36415, x27948, x84599);
  nand n36416(x36416, x27948, x84600);
  nand n36417(x36417, x27948, x84601);
  nand n36418(x36418, x27948, x84602);
  nand n36419(x36419, x27948, x84603);
  nand n36420(x36420, x27948, x36342);
  nand n36421(x36421, x27948, x36345);
  nand n36422(x36422, x27948, x36348);
  nand n36423(x36423, x27948, x36351);
  nand n36424(x36424, x27948, x36354);
  nand n36425(x36425, x27948, x36357);
  nand n36426(x36426, x27948, x36360);
  nand n36427(x36427, x27948, x36363);
  nand n36428(x36428, x27889, x84596);
  nand n36429(x36429, x27948, x36366);
  nand n36430(x36430, x36429, x36428);
  nand n36431(x36431, x27889, x84597);
  nand n36432(x36432, x27948, x36369);
  nand n36433(x36433, x36432, x36431);
  nand n36434(x36434, x27889, x84598);
  nand n36435(x36435, x27948, x36372);
  nand n36436(x36436, x36435, x36434);
  nand n36437(x36437, x27889, x84599);
  nand n36438(x36438, x27948, x36375);
  nand n36439(x36439, x36438, x36437);
  nand n36440(x36440, x27889, x84600);
  nand n36441(x36441, x27948, x36378);
  nand n36442(x36442, x36441, x36440);
  nand n36443(x36443, x27889, x84601);
  nand n36444(x36444, x27948, x36381);
  nand n36445(x36445, x36444, x36443);
  nand n36446(x36446, x27889, x84602);
  nand n36447(x36447, x27948, x36384);
  nand n36448(x36448, x36447, x36446);
  nand n36449(x36449, x27889, x84603);
  nand n36450(x36450, x27948, x36387);
  nand n36451(x36451, x36450, x36449);
  nand n36452(x36452, x27889, x36342);
  nand n36453(x36453, x27948, x36390);
  nand n36454(x36454, x36453, x36452);
  nand n36455(x36455, x27889, x36345);
  nand n36456(x36456, x27948, x36393);
  nand n36457(x36457, x36456, x36455);
  nand n36458(x36458, x27889, x36348);
  nand n36459(x36459, x27948, x36396);
  nand n36460(x36460, x36459, x36458);
  nand n36461(x36461, x27889, x36351);
  nand n36462(x36462, x27948, x36399);
  nand n36463(x36463, x36462, x36461);
  nand n36464(x36464, x27889, x36354);
  nand n36465(x36465, x27948, x36402);
  nand n36466(x36466, x36465, x36464);
  nand n36467(x36467, x27889, x36357);
  nand n36468(x36468, x27948, x36405);
  nand n36469(x36469, x36468, x36467);
  nand n36470(x36470, x27889, x36360);
  nand n36471(x36471, x27948, x36408);
  nand n36472(x36472, x36471, x36470);
  nand n36473(x36473, x27889, x36363);
  nand n36474(x36474, x27948, x36411);
  nand n36475(x36475, x36474, x36473);
  nand n36476(x36476, x36089, x29005);
  nand n36477(x36477, x36090, x29009);
  nand n36478(x36478, x36092, x29015);
  nand n36479(x36479, x36094, x29022);
  nand n36480(x36480, x36096, x29032);
  nand n36481(x36481, x36098, x29044);
  nand n36482(x36482, x36100, x29057);
  nand n36483(x36483, x36102, x29073);
  nand n36484(x36484, x36104, x29091);
  nand n36485(x36485, x36106, x29110);
  nand n36486(x36486, x36108, x29132);
  nand n36487(x36487, x36110, x29156);
  nand n36488(x36488, x36112, x29181);
  nand n36489(x36489, x36114, x29209);
  nand n36490(x36490, x36116, x29239);
  nand n36491(x36491, x36118, x29270);
  nand n36492(x36492, x36120, x29304);
  nand n36493(x36493, x36122, x29340);
  nand n36494(x36494, x36124, x29377);
  nand n36495(x36495, x36126, x29417);
  nand n36496(x36496, x36128, x29459);
  nand n36497(x36497, x36130, x29502);
  nand n36498(x36498, x36132, x29548);
  nand n36499(x36499, x36134, x29596);
  nand n36500(x36500, x36136, x29645);
  nand n36501(x36501, x36138, x29697);
  nand n36502(x36502, x36140, x29751);
  nand n36503(x36503, x36142, x29806);
  nand n36504(x36504, x36144, x29864);
  nand n36505(x36505, x36146, x29924);
  nand n36506(x36506, x36148, x29985);
  nand n36507(x36507, x27883, x36478);
  nand n36508(x36508, x27945, x36476);
  nand n36509(x36509, x36508, x36507);
  nand n36510(x36510, x27883, x36479);
  nand n36511(x36511, x27945, x36477);
  nand n36512(x36512, x36511, x36510);
  nand n36513(x36513, x27883, x36480);
  nand n36514(x36514, x27945, x36478);
  nand n36515(x36515, x36514, x36513);
  nand n36516(x36516, x27883, x36481);
  nand n36517(x36517, x27945, x36479);
  nand n36518(x36518, x36517, x36516);
  nand n36519(x36519, x27883, x36482);
  nand n36520(x36520, x27945, x36480);
  nand n36521(x36521, x36520, x36519);
  nand n36522(x36522, x27883, x36483);
  nand n36523(x36523, x27945, x36481);
  nand n36524(x36524, x36523, x36522);
  nand n36525(x36525, x27883, x36484);
  nand n36526(x36526, x27945, x36482);
  nand n36527(x36527, x36526, x36525);
  nand n36528(x36528, x27883, x36485);
  nand n36529(x36529, x27945, x36483);
  nand n36530(x36530, x36529, x36528);
  nand n36531(x36531, x27883, x36486);
  nand n36532(x36532, x27945, x36484);
  nand n36533(x36533, x36532, x36531);
  nand n36534(x36534, x27883, x36487);
  nand n36535(x36535, x27945, x36485);
  nand n36536(x36536, x36535, x36534);
  nand n36537(x36537, x27883, x36488);
  nand n36538(x36538, x27945, x36486);
  nand n36539(x36539, x36538, x36537);
  nand n36540(x36540, x27883, x36489);
  nand n36541(x36541, x27945, x36487);
  nand n36542(x36542, x36541, x36540);
  nand n36543(x36543, x27883, x36490);
  nand n36544(x36544, x27945, x36488);
  nand n36545(x36545, x36544, x36543);
  nand n36546(x36546, x27883, x36491);
  nand n36547(x36547, x27945, x36489);
  nand n36548(x36548, x36547, x36546);
  nand n36549(x36549, x27883, x36492);
  nand n36550(x36550, x27945, x36490);
  nand n36551(x36551, x36550, x36549);
  nand n36552(x36552, x27883, x36493);
  nand n36553(x36553, x27945, x36491);
  nand n36554(x36554, x36553, x36552);
  nand n36555(x36555, x27883, x36494);
  nand n36556(x36556, x27945, x36492);
  nand n36557(x36557, x36556, x36555);
  nand n36558(x36558, x27883, x36495);
  nand n36559(x36559, x27945, x36493);
  nand n36560(x36560, x36559, x36558);
  nand n36561(x36561, x27883, x36496);
  nand n36562(x36562, x27945, x36494);
  nand n36563(x36563, x36562, x36561);
  nand n36564(x36564, x27883, x36497);
  nand n36565(x36565, x27945, x36495);
  nand n36566(x36566, x36565, x36564);
  nand n36567(x36567, x27883, x36498);
  nand n36568(x36568, x27945, x36496);
  nand n36569(x36569, x36568, x36567);
  nand n36570(x36570, x27883, x36499);
  nand n36571(x36571, x27945, x36497);
  nand n36572(x36572, x36571, x36570);
  nand n36573(x36573, x27883, x36500);
  nand n36574(x36574, x27945, x36498);
  nand n36575(x36575, x36574, x36573);
  nand n36576(x36576, x27883, x36501);
  nand n36577(x36577, x27945, x36499);
  nand n36578(x36578, x36577, x36576);
  nand n36579(x36579, x27883, x36502);
  nand n36580(x36580, x27945, x36500);
  nand n36581(x36581, x36580, x36579);
  nand n36582(x36582, x27883, x36503);
  nand n36583(x36583, x27945, x36501);
  nand n36584(x36584, x36583, x36582);
  nand n36585(x36585, x27883, x36504);
  nand n36586(x36586, x27945, x36502);
  nand n36587(x36587, x36586, x36585);
  nand n36588(x36588, x27883, x36505);
  nand n36589(x36589, x27945, x36503);
  nand n36590(x36590, x36589, x36588);
  nand n36591(x36591, x27883, x36506);
  nand n36592(x36592, x27945, x36504);
  nand n36593(x36593, x36592, x36591);
  nand n36594(x36594, x27883, x84620);
  nand n36595(x36595, x27945, x36505);
  nand n36596(x36596, x36595, x36594);
  nand n36597(x36597, x27945, x36506);
  nand n36598(x36598, x27945, x84620);
  nand n36599(x36599, x27885, x36521);
  nand n36600(x36600, x27946, x36509);
  nand n36601(x36601, x36600, x36599);
  nand n36602(x36602, x27885, x36524);
  nand n36603(x36603, x27946, x36512);
  nand n36604(x36604, x36603, x36602);
  nand n36605(x36605, x27885, x36527);
  nand n36606(x36606, x27946, x36515);
  nand n36607(x36607, x36606, x36605);
  nand n36608(x36608, x27885, x36530);
  nand n36609(x36609, x27946, x36518);
  nand n36610(x36610, x36609, x36608);
  nand n36611(x36611, x27885, x36533);
  nand n36612(x36612, x27946, x36521);
  nand n36613(x36613, x36612, x36611);
  nand n36614(x36614, x27885, x36536);
  nand n36615(x36615, x27946, x36524);
  nand n36616(x36616, x36615, x36614);
  nand n36617(x36617, x27885, x36539);
  nand n36618(x36618, x27946, x36527);
  nand n36619(x36619, x36618, x36617);
  nand n36620(x36620, x27885, x36542);
  nand n36621(x36621, x27946, x36530);
  nand n36622(x36622, x36621, x36620);
  nand n36623(x36623, x27885, x36545);
  nand n36624(x36624, x27946, x36533);
  nand n36625(x36625, x36624, x36623);
  nand n36626(x36626, x27885, x36548);
  nand n36627(x36627, x27946, x36536);
  nand n36628(x36628, x36627, x36626);
  nand n36629(x36629, x27885, x36551);
  nand n36630(x36630, x27946, x36539);
  nand n36631(x36631, x36630, x36629);
  nand n36632(x36632, x27885, x36554);
  nand n36633(x36633, x27946, x36542);
  nand n36634(x36634, x36633, x36632);
  nand n36635(x36635, x27885, x36557);
  nand n36636(x36636, x27946, x36545);
  nand n36637(x36637, x36636, x36635);
  nand n36638(x36638, x27885, x36560);
  nand n36639(x36639, x27946, x36548);
  nand n36640(x36640, x36639, x36638);
  nand n36641(x36641, x27885, x36563);
  nand n36642(x36642, x27946, x36551);
  nand n36643(x36643, x36642, x36641);
  nand n36644(x36644, x27885, x36566);
  nand n36645(x36645, x27946, x36554);
  nand n36646(x36646, x36645, x36644);
  nand n36647(x36647, x27885, x36569);
  nand n36648(x36648, x27946, x36557);
  nand n36649(x36649, x36648, x36647);
  nand n36650(x36650, x27885, x36572);
  nand n36651(x36651, x27946, x36560);
  nand n36652(x36652, x36651, x36650);
  nand n36653(x36653, x27885, x36575);
  nand n36654(x36654, x27946, x36563);
  nand n36655(x36655, x36654, x36653);
  nand n36656(x36656, x27885, x36578);
  nand n36657(x36657, x27946, x36566);
  nand n36658(x36658, x36657, x36656);
  nand n36659(x36659, x27885, x36581);
  nand n36660(x36660, x27946, x36569);
  nand n36661(x36661, x36660, x36659);
  nand n36662(x36662, x27885, x36584);
  nand n36663(x36663, x27946, x36572);
  nand n36664(x36664, x36663, x36662);
  nand n36665(x36665, x27885, x36587);
  nand n36666(x36666, x27946, x36575);
  nand n36667(x36667, x36666, x36665);
  nand n36668(x36668, x27885, x36590);
  nand n36669(x36669, x27946, x36578);
  nand n36670(x36670, x36669, x36668);
  nand n36671(x36671, x27885, x36593);
  nand n36672(x36672, x27946, x36581);
  nand n36673(x36673, x36672, x36671);
  nand n36674(x36674, x27885, x36596);
  nand n36675(x36675, x27946, x36584);
  nand n36676(x36676, x36675, x36674);
  nand n36677(x36677, x27885, x84621);
  nand n36678(x36678, x27946, x36587);
  nand n36679(x36679, x36678, x36677);
  nand n36680(x36680, x27885, x84622);
  nand n36681(x36681, x27946, x36590);
  nand n36682(x36682, x36681, x36680);
  nand n36683(x36683, x27946, x36593);
  nand n36684(x36684, x27946, x36596);
  nand n36685(x36685, x27946, x84621);
  nand n36686(x36686, x27946, x84622);
  nand n36687(x36687, x27887, x36625);
  nand n36688(x36688, x27947, x36601);
  nand n36689(x36689, x36688, x36687);
  nand n36690(x36690, x27887, x36628);
  nand n36691(x36691, x27947, x36604);
  nand n36692(x36692, x36691, x36690);
  nand n36693(x36693, x27887, x36631);
  nand n36694(x36694, x27947, x36607);
  nand n36695(x36695, x36694, x36693);
  nand n36696(x36696, x27887, x36634);
  nand n36697(x36697, x27947, x36610);
  nand n36698(x36698, x36697, x36696);
  nand n36699(x36699, x27887, x36637);
  nand n36700(x36700, x27947, x36613);
  nand n36701(x36701, x36700, x36699);
  nand n36702(x36702, x27887, x36640);
  nand n36703(x36703, x27947, x36616);
  nand n36704(x36704, x36703, x36702);
  nand n36705(x36705, x27887, x36643);
  nand n36706(x36706, x27947, x36619);
  nand n36707(x36707, x36706, x36705);
  nand n36708(x36708, x27887, x36646);
  nand n36709(x36709, x27947, x36622);
  nand n36710(x36710, x36709, x36708);
  nand n36711(x36711, x27887, x36649);
  nand n36712(x36712, x27947, x36625);
  nand n36713(x36713, x36712, x36711);
  nand n36714(x36714, x27887, x36652);
  nand n36715(x36715, x27947, x36628);
  nand n36716(x36716, x36715, x36714);
  nand n36717(x36717, x27887, x36655);
  nand n36718(x36718, x27947, x36631);
  nand n36719(x36719, x36718, x36717);
  nand n36720(x36720, x27887, x36658);
  nand n36721(x36721, x27947, x36634);
  nand n36722(x36722, x36721, x36720);
  nand n36723(x36723, x27887, x36661);
  nand n36724(x36724, x27947, x36637);
  nand n36725(x36725, x36724, x36723);
  nand n36726(x36726, x27887, x36664);
  nand n36727(x36727, x27947, x36640);
  nand n36728(x36728, x36727, x36726);
  nand n36729(x36729, x27887, x36667);
  nand n36730(x36730, x27947, x36643);
  nand n36731(x36731, x36730, x36729);
  nand n36732(x36732, x27887, x36670);
  nand n36733(x36733, x27947, x36646);
  nand n36734(x36734, x36733, x36732);
  nand n36735(x36735, x27887, x36673);
  nand n36736(x36736, x27947, x36649);
  nand n36737(x36737, x36736, x36735);
  nand n36738(x36738, x27887, x36676);
  nand n36739(x36739, x27947, x36652);
  nand n36740(x36740, x36739, x36738);
  nand n36741(x36741, x27887, x36679);
  nand n36742(x36742, x27947, x36655);
  nand n36743(x36743, x36742, x36741);
  nand n36744(x36744, x27887, x36682);
  nand n36745(x36745, x27947, x36658);
  nand n36746(x36746, x36745, x36744);
  nand n36747(x36747, x27887, x84623);
  nand n36748(x36748, x27947, x36661);
  nand n36749(x36749, x36748, x36747);
  nand n36750(x36750, x27887, x84624);
  nand n36751(x36751, x27947, x36664);
  nand n36752(x36752, x36751, x36750);
  nand n36753(x36753, x27887, x84625);
  nand n36754(x36754, x27947, x36667);
  nand n36755(x36755, x36754, x36753);
  nand n36756(x36756, x27887, x84626);
  nand n36757(x36757, x27947, x36670);
  nand n36758(x36758, x36757, x36756);
  nand n36759(x36759, x27947, x36673);
  nand n36760(x36760, x27947, x36676);
  nand n36761(x36761, x27947, x36679);
  nand n36762(x36762, x27947, x36682);
  nand n36763(x36763, x27947, x84623);
  nand n36764(x36764, x27947, x84624);
  nand n36765(x36765, x27947, x84625);
  nand n36766(x36766, x27947, x84626);
  nand n36767(x36767, x27889, x36737);
  nand n36768(x36768, x27948, x36689);
  nand n36769(x36769, x36768, x36767);
  nand n36770(x36770, x27889, x36740);
  nand n36771(x36771, x27948, x36692);
  nand n36772(x36772, x36771, x36770);
  nand n36773(x36773, x27889, x36743);
  nand n36774(x36774, x27948, x36695);
  nand n36775(x36775, x36774, x36773);
  nand n36776(x36776, x27889, x36746);
  nand n36777(x36777, x27948, x36698);
  nand n36778(x36778, x36777, x36776);
  nand n36779(x36779, x27889, x36749);
  nand n36780(x36780, x27948, x36701);
  nand n36781(x36781, x36780, x36779);
  nand n36782(x36782, x27889, x36752);
  nand n36783(x36783, x27948, x36704);
  nand n36784(x36784, x36783, x36782);
  nand n36785(x36785, x27889, x36755);
  nand n36786(x36786, x27948, x36707);
  nand n36787(x36787, x36786, x36785);
  nand n36788(x36788, x27889, x36758);
  nand n36789(x36789, x27948, x36710);
  nand n36790(x36790, x36789, x36788);
  nand n36791(x36791, x27889, x84627);
  nand n36792(x36792, x27948, x36713);
  nand n36793(x36793, x36792, x36791);
  nand n36794(x36794, x27889, x84628);
  nand n36795(x36795, x27948, x36716);
  nand n36796(x36796, x36795, x36794);
  nand n36797(x36797, x27889, x84629);
  nand n36798(x36798, x27948, x36719);
  nand n36799(x36799, x36798, x36797);
  nand n36800(x36800, x27889, x84630);
  nand n36801(x36801, x27948, x36722);
  nand n36802(x36802, x36801, x36800);
  nand n36803(x36803, x27889, x84631);
  nand n36804(x36804, x27948, x36725);
  nand n36805(x36805, x36804, x36803);
  nand n36806(x36806, x27889, x84632);
  nand n36807(x36807, x27948, x36728);
  nand n36808(x36808, x36807, x36806);
  nand n36809(x36809, x27889, x84633);
  nand n36810(x36810, x27948, x36731);
  nand n36811(x36811, x36810, x36809);
  nand n36812(x36812, x27889, x84634);
  nand n36813(x36813, x27948, x36734);
  nand n36814(x36814, x36813, x36812);
  nand n36815(x36815, x27948, x36737);
  nand n36816(x36816, x27948, x36740);
  nand n36817(x36817, x27948, x36743);
  nand n36818(x36818, x27948, x36746);
  nand n36819(x36819, x27948, x36749);
  nand n36820(x36820, x27948, x36752);
  nand n36821(x36821, x27948, x36755);
  nand n36822(x36822, x27948, x36758);
  nand n36823(x36823, x27948, x84627);
  nand n36824(x36824, x27948, x84628);
  nand n36825(x36825, x27948, x84629);
  nand n36826(x36826, x27948, x84630);
  nand n36827(x36827, x27948, x84631);
  nand n36828(x36828, x27948, x84632);
  nand n36829(x36829, x27948, x84633);
  nand n36830(x36830, x27948, x84634);
  nand n36831(x36831, x71977, x27881);
  nand n36832(x36832, x16876, x36769);
  nand n36833(x36833, x36832, x25733);
  nand n36834(x36834, x71977, x84604);
  nand n36835(x36835, x16876, x35960);
  nand n36836(x36836, x71977, x28848);
  nand n36837(x36837, x16876, x28848);
  nand n36838(x36838, x36837, x36836);
  nand n36839(x36839, x71977, x36026);
  nand n36840(x36840, x16876, x35993);
  nand n36841(x36841, x36840, x36839);
  nand n36842(x36842, x71977, x35960);
  nand n36843(x36843, x36832, x36842);
  nand n36844(x36844, x16876, x28074);
  nand n36845(x36845, x36844, x36842);
  nand n36846(x36846, x71977, x72537);
  nand n36847(x36847, x25749, x84651);
  nand n36848(x36848, x71982, x36833);
  nand n36849(x36849, x25749, x84652);
  nand n36850(x36850, x36849, x36848);
  nand n36851(x36851, x71982, x84653);
  nand n36852(x36852, x25749, x36838);
  nand n36853(x36853, x36852, x36851);
  nand n36854(x36854, x71982, x36841);
  nand n36855(x36855, x25749, x36843);
  nand n36856(x36856, x36855, x36854);
  nand n36857(x36857, x71982, x84652);
  nand n36858(x36858, x25749, x84653);
  nand n36859(x36859, x36858, x36857);
  nand n36860(x36860, x71982, x36838);
  nand n36861(x36861, x25749, x36841);
  nand n36862(x36862, x36861, x36860);
  nand n36863(x36863, x71982, x36845);
  nand n36864(x36864, x25749, x84654);
  nand n36865(x36865, x36864, x36863);
  nand n36866(x36866, x71987, x84655);
  nand n36867(x36867, x25772, x36850);
  nand n36868(x36868, x36867, x25771);
  nand n36869(x36869, x71987, x36853);
  nand n36870(x36870, x25772, x36856);
  nand n36871(x36871, x36870, x36869);
  nand n36872(x36872, x71987, x36859);
  nand n36873(x36873, x25772, x36862);
  nand n36874(x36874, x36873, x36872);
  nand n36875(x36875, x71987, x36865);
  nand n36876(x36876, x25782, x84656);
  nand n36877(x36877, x71992, x36868);
  nand n36878(x36878, x25782, x36871);
  nand n36879(x36879, x36878, x36877);
  nand n36880(x36880, x71992, x36874);
  nand n36881(x36881, x25782, x84657);
  nand n36882(x36882, x36881, x36880);
  nand n36883(x36883, x25790, x84658);
  nand n36884(x36884, x71997, x36879);
  nand n36885(x36885, x25790, x36882);
  nand n36886(x36886, x36885, x36884);
  nand n36887(x36887, x72002, x84659);
  nand n36888(x36888, x25796, x36886);
  nand n36889(x36889, x36888, x36887);
  nand n36890(x36890, x71977, x27883);
  nand n36891(x36891, x16876, x36772);
  nand n36892(x36892, x36891, x25801);
  nand n36893(x36893, x71977, x84605);
  nand n36894(x36894, x16876, x84557);
  nand n36895(x36895, x71977, x28853);
  nand n36896(x36896, x16876, x28853);
  nand n36897(x36897, x36896, x36895);
  nand n36898(x36898, x71977, x36028);
  nand n36899(x36899, x16876, x35994);
  nand n36900(x36900, x36899, x36898);
  nand n36901(x36901, x71977, x29012);
  nand n36902(x36902, x36891, x36901);
  nand n36903(x36903, x16876, x28080);
  nand n36904(x36904, x36903, x36901);
  nand n36905(x36905, x71977, x35839);
  nand n36906(x36906, x25749, x84660);
  nand n36907(x36907, x71982, x36892);
  nand n36908(x36908, x25749, x84661);
  nand n36909(x36909, x36908, x36907);
  nand n36910(x36910, x71982, x84662);
  nand n36911(x36911, x25749, x36897);
  nand n36912(x36912, x36911, x36910);
  nand n36913(x36913, x71982, x36900);
  nand n36914(x36914, x25749, x36902);
  nand n36915(x36915, x36914, x36913);
  nand n36916(x36916, x71982, x84661);
  nand n36917(x36917, x25749, x84662);
  nand n36918(x36918, x36917, x36916);
  nand n36919(x36919, x71982, x36897);
  nand n36920(x36920, x25749, x36900);
  nand n36921(x36921, x36920, x36919);
  nand n36922(x36922, x71982, x36904);
  nand n36923(x36923, x25749, x84663);
  nand n36924(x36924, x36923, x36922);
  nand n36925(x36925, x71987, x84664);
  nand n36926(x36926, x25772, x36909);
  nand n36927(x36927, x36926, x25838);
  nand n36928(x36928, x71987, x36912);
  nand n36929(x36929, x25772, x36915);
  nand n36930(x36930, x36929, x36928);
  nand n36931(x36931, x71987, x36918);
  nand n36932(x36932, x25772, x36921);
  nand n36933(x36933, x36932, x36931);
  nand n36934(x36934, x71987, x36924);
  nand n36935(x36935, x25782, x84665);
  nand n36936(x36936, x71992, x36927);
  nand n36937(x36937, x25782, x36930);
  nand n36938(x36938, x36937, x36936);
  nand n36939(x36939, x71992, x36933);
  nand n36940(x36940, x25782, x84666);
  nand n36941(x36941, x36940, x36939);
  nand n36942(x36942, x25790, x84667);
  nand n36943(x36943, x71997, x36938);
  nand n36944(x36944, x25790, x36941);
  nand n36945(x36945, x36944, x36943);
  nand n36946(x36946, x72002, x84668);
  nand n36947(x36947, x25796, x36945);
  nand n36948(x36948, x36947, x36946);
  nand n36949(x36949, x71977, x27885);
  nand n36950(x36950, x16876, x36775);
  nand n36951(x36951, x36950, x25864);
  nand n36952(x36952, x71977, x84606);
  nand n36953(x36953, x16876, x84558);
  nand n36954(x36954, x71977, x28858);
  nand n36955(x36955, x16876, x28858);
  nand n36956(x36956, x36955, x36954);
  nand n36957(x36957, x71977, x36030);
  nand n36958(x36958, x16876, x35995);
  nand n36959(x36959, x36958, x36957);
  nand n36960(x36960, x71977, x29027);
  nand n36961(x36961, x36950, x36960);
  nand n36962(x36962, x16876, x28086);
  nand n36963(x36963, x36962, x36960);
  nand n36964(x36964, x71977, x35843);
  nand n36965(x36965, x25749, x84669);
  nand n36966(x36966, x71982, x36951);
  nand n36967(x36967, x25749, x84670);
  nand n36968(x36968, x36967, x36966);
  nand n36969(x36969, x71982, x84671);
  nand n36970(x36970, x25749, x36956);
  nand n36971(x36971, x36970, x36969);
  nand n36972(x36972, x71982, x36959);
  nand n36973(x36973, x25749, x36961);
  nand n36974(x36974, x36973, x36972);
  nand n36975(x36975, x71982, x84670);
  nand n36976(x36976, x25749, x84671);
  nand n36977(x36977, x36976, x36975);
  nand n36978(x36978, x71982, x36956);
  nand n36979(x36979, x25749, x36959);
  nand n36980(x36980, x36979, x36978);
  nand n36981(x36981, x71982, x36963);
  nand n36982(x36982, x25749, x84672);
  nand n36983(x36983, x36982, x36981);
  nand n36984(x36984, x71987, x84673);
  nand n36985(x36985, x25772, x36968);
  nand n36986(x36986, x36985, x25901);
  nand n36987(x36987, x71987, x36971);
  nand n36988(x36988, x25772, x36974);
  nand n36989(x36989, x36988, x36987);
  nand n36990(x36990, x71987, x36977);
  nand n36991(x36991, x25772, x36980);
  nand n36992(x36992, x36991, x36990);
  nand n36993(x36993, x71987, x36983);
  nand n36994(x36994, x25782, x84674);
  nand n36995(x36995, x71992, x36986);
  nand n36996(x36996, x25782, x36989);
  nand n36997(x36997, x36996, x36995);
  nand n36998(x36998, x71992, x36992);
  nand n36999(x36999, x25782, x84675);
  nand n37000(x37000, x36999, x36998);
  nand n37001(x37001, x25790, x84676);
  nand n37002(x37002, x71997, x36997);
  nand n37003(x37003, x25790, x37000);
  nand n37004(x37004, x37003, x37002);
  nand n37005(x37005, x72002, x84677);
  nand n37006(x37006, x25796, x37004);
  nand n37007(x37007, x37006, x37005);
  nand n37008(x37008, x71977, x27887);
  nand n37009(x37009, x16876, x36778);
  nand n37010(x37010, x37009, x25927);
  nand n37011(x37011, x71977, x84607);
  nand n37012(x37012, x16876, x84559);
  nand n37013(x37013, x71977, x28863);
  nand n37014(x37014, x16876, x28863);
  nand n37015(x37015, x37014, x37013);
  nand n37016(x37016, x71977, x36032);
  nand n37017(x37017, x16876, x35996);
  nand n37018(x37018, x37017, x37016);
  nand n37019(x37019, x71977, x29051);
  nand n37020(x37020, x37009, x37019);
  nand n37021(x37021, x16876, x28092);
  nand n37022(x37022, x37021, x37019);
  nand n37023(x37023, x71977, x35847);
  nand n37024(x37024, x25749, x84678);
  nand n37025(x37025, x71982, x37010);
  nand n37026(x37026, x25749, x84679);
  nand n37027(x37027, x37026, x37025);
  nand n37028(x37028, x71982, x84680);
  nand n37029(x37029, x25749, x37015);
  nand n37030(x37030, x37029, x37028);
  nand n37031(x37031, x71982, x37018);
  nand n37032(x37032, x25749, x37020);
  nand n37033(x37033, x37032, x37031);
  nand n37034(x37034, x71982, x84679);
  nand n37035(x37035, x25749, x84680);
  nand n37036(x37036, x37035, x37034);
  nand n37037(x37037, x71982, x37015);
  nand n37038(x37038, x25749, x37018);
  nand n37039(x37039, x37038, x37037);
  nand n37040(x37040, x71982, x37022);
  nand n37041(x37041, x25749, x84681);
  nand n37042(x37042, x37041, x37040);
  nand n37043(x37043, x71987, x84682);
  nand n37044(x37044, x25772, x37027);
  nand n37045(x37045, x37044, x25964);
  nand n37046(x37046, x71987, x37030);
  nand n37047(x37047, x25772, x37033);
  nand n37048(x37048, x37047, x37046);
  nand n37049(x37049, x71987, x37036);
  nand n37050(x37050, x25772, x37039);
  nand n37051(x37051, x37050, x37049);
  nand n37052(x37052, x71987, x37042);
  nand n37053(x37053, x25782, x84683);
  nand n37054(x37054, x71992, x37045);
  nand n37055(x37055, x25782, x37048);
  nand n37056(x37056, x37055, x37054);
  nand n37057(x37057, x71992, x37051);
  nand n37058(x37058, x25782, x84684);
  nand n37059(x37059, x37058, x37057);
  nand n37060(x37060, x25790, x84685);
  nand n37061(x37061, x71997, x37056);
  nand n37062(x37062, x25790, x37059);
  nand n37063(x37063, x37062, x37061);
  nand n37064(x37064, x72002, x84686);
  nand n37065(x37065, x25796, x37063);
  nand n37066(x37066, x37065, x37064);
  nand n37067(x37067, x71977, x27889);
  nand n37068(x37068, x16876, x36781);
  nand n37069(x37069, x37068, x25990);
  nand n37070(x37070, x71977, x84608);
  nand n37071(x37071, x16876, x84560);
  nand n37072(x37072, x71977, x28868);
  nand n37073(x37073, x16876, x28868);
  nand n37074(x37074, x37073, x37072);
  nand n37075(x37075, x71977, x36034);
  nand n37076(x37076, x16876, x35997);
  nand n37077(x37077, x37076, x37075);
  nand n37078(x37078, x71977, x29082);
  nand n37079(x37079, x37068, x37078);
  nand n37080(x37080, x16876, x28098);
  nand n37081(x37081, x37080, x37078);
  nand n37082(x37082, x71977, x35851);
  nand n37083(x37083, x25749, x84687);
  nand n37084(x37084, x71982, x37069);
  nand n37085(x37085, x25749, x84688);
  nand n37086(x37086, x37085, x37084);
  nand n37087(x37087, x71982, x84689);
  nand n37088(x37088, x25749, x37074);
  nand n37089(x37089, x37088, x37087);
  nand n37090(x37090, x71982, x37077);
  nand n37091(x37091, x25749, x37079);
  nand n37092(x37092, x37091, x37090);
  nand n37093(x37093, x71982, x84688);
  nand n37094(x37094, x25749, x84689);
  nand n37095(x37095, x37094, x37093);
  nand n37096(x37096, x71982, x37074);
  nand n37097(x37097, x25749, x37077);
  nand n37098(x37098, x37097, x37096);
  nand n37099(x37099, x71982, x37081);
  nand n37100(x37100, x25749, x84690);
  nand n37101(x37101, x37100, x37099);
  nand n37102(x37102, x71987, x84691);
  nand n37103(x37103, x25772, x37086);
  nand n37104(x37104, x37103, x26027);
  nand n37105(x37105, x71987, x37089);
  nand n37106(x37106, x25772, x37092);
  nand n37107(x37107, x37106, x37105);
  nand n37108(x37108, x71987, x37095);
  nand n37109(x37109, x25772, x37098);
  nand n37110(x37110, x37109, x37108);
  nand n37111(x37111, x71987, x37101);
  nand n37112(x37112, x25782, x84692);
  nand n37113(x37113, x71992, x37104);
  nand n37114(x37114, x25782, x37107);
  nand n37115(x37115, x37114, x37113);
  nand n37116(x37116, x71992, x37110);
  nand n37117(x37117, x25782, x84693);
  nand n37118(x37118, x37117, x37116);
  nand n37119(x37119, x25790, x84694);
  nand n37120(x37120, x71997, x37115);
  nand n37121(x37121, x25790, x37118);
  nand n37122(x37122, x37121, x37120);
  nand n37123(x37123, x72002, x84695);
  nand n37124(x37124, x25796, x37122);
  nand n37125(x37125, x37124, x37123);
  nand n37126(x37126, x71977, x27891);
  nand n37127(x37127, x16876, x36784);
  nand n37128(x37128, x37127, x26053);
  nand n37129(x37129, x71977, x84609);
  nand n37130(x37130, x16876, x84561);
  nand n37131(x37131, x71977, x28873);
  nand n37132(x37132, x16876, x28873);
  nand n37133(x37133, x37132, x37131);
  nand n37134(x37134, x71977, x36036);
  nand n37135(x37135, x16876, x35998);
  nand n37136(x37136, x37135, x37134);
  nand n37137(x37137, x71977, x29121);
  nand n37138(x37138, x37127, x37137);
  nand n37139(x37139, x16876, x28104);
  nand n37140(x37140, x37139, x37137);
  nand n37141(x37141, x71977, x35855);
  nand n37142(x37142, x25749, x84696);
  nand n37143(x37143, x71982, x37128);
  nand n37144(x37144, x25749, x84697);
  nand n37145(x37145, x37144, x37143);
  nand n37146(x37146, x71982, x84698);
  nand n37147(x37147, x25749, x37133);
  nand n37148(x37148, x37147, x37146);
  nand n37149(x37149, x71982, x37136);
  nand n37150(x37150, x25749, x37138);
  nand n37151(x37151, x37150, x37149);
  nand n37152(x37152, x71982, x84697);
  nand n37153(x37153, x25749, x84698);
  nand n37154(x37154, x37153, x37152);
  nand n37155(x37155, x71982, x37133);
  nand n37156(x37156, x25749, x37136);
  nand n37157(x37157, x37156, x37155);
  nand n37158(x37158, x71982, x37140);
  nand n37159(x37159, x25749, x84699);
  nand n37160(x37160, x37159, x37158);
  nand n37161(x37161, x71987, x84700);
  nand n37162(x37162, x25772, x37145);
  nand n37163(x37163, x37162, x26090);
  nand n37164(x37164, x71987, x37148);
  nand n37165(x37165, x25772, x37151);
  nand n37166(x37166, x37165, x37164);
  nand n37167(x37167, x71987, x37154);
  nand n37168(x37168, x25772, x37157);
  nand n37169(x37169, x37168, x37167);
  nand n37170(x37170, x71987, x37160);
  nand n37171(x37171, x25782, x84701);
  nand n37172(x37172, x71992, x37163);
  nand n37173(x37173, x25782, x37166);
  nand n37174(x37174, x37173, x37172);
  nand n37175(x37175, x71992, x37169);
  nand n37176(x37176, x25782, x84702);
  nand n37177(x37177, x37176, x37175);
  nand n37178(x37178, x25790, x84703);
  nand n37179(x37179, x71997, x37174);
  nand n37180(x37180, x25790, x37177);
  nand n37181(x37181, x37180, x37179);
  nand n37182(x37182, x72002, x84704);
  nand n37183(x37183, x25796, x37181);
  nand n37184(x37184, x37183, x37182);
  nand n37185(x37185, x71977, x27893);
  nand n37186(x37186, x16876, x36787);
  nand n37187(x37187, x37186, x26116);
  nand n37188(x37188, x71977, x84610);
  nand n37189(x37189, x16876, x35503);
  nand n37190(x37190, x71977, x28878);
  nand n37191(x37191, x16876, x28878);
  nand n37192(x37192, x37191, x37190);
  nand n37193(x37193, x71977, x36038);
  nand n37194(x37194, x16876, x35999);
  nand n37195(x37195, x37194, x37193);
  nand n37196(x37196, x71977, x29169);
  nand n37197(x37197, x37186, x37196);
  nand n37198(x37198, x16876, x28110);
  nand n37199(x37199, x37198, x37196);
  nand n37200(x37200, x71977, x35859);
  nand n37201(x37201, x25749, x84705);
  nand n37202(x37202, x71982, x37187);
  nand n37203(x37203, x25749, x84706);
  nand n37204(x37204, x37203, x37202);
  nand n37205(x37205, x71982, x84707);
  nand n37206(x37206, x25749, x37192);
  nand n37207(x37207, x37206, x37205);
  nand n37208(x37208, x71982, x37195);
  nand n37209(x37209, x25749, x37197);
  nand n37210(x37210, x37209, x37208);
  nand n37211(x37211, x71982, x84706);
  nand n37212(x37212, x25749, x84707);
  nand n37213(x37213, x37212, x37211);
  nand n37214(x37214, x71982, x37192);
  nand n37215(x37215, x25749, x37195);
  nand n37216(x37216, x37215, x37214);
  nand n37217(x37217, x71982, x37199);
  nand n37218(x37218, x25749, x84708);
  nand n37219(x37219, x37218, x37217);
  nand n37220(x37220, x71987, x84709);
  nand n37221(x37221, x25772, x37204);
  nand n37222(x37222, x37221, x26153);
  nand n37223(x37223, x71987, x37207);
  nand n37224(x37224, x25772, x37210);
  nand n37225(x37225, x37224, x37223);
  nand n37226(x37226, x71987, x37213);
  nand n37227(x37227, x25772, x37216);
  nand n37228(x37228, x37227, x37226);
  nand n37229(x37229, x71987, x37219);
  nand n37230(x37230, x25782, x84710);
  nand n37231(x37231, x71992, x37222);
  nand n37232(x37232, x25782, x37225);
  nand n37233(x37233, x37232, x37231);
  nand n37234(x37234, x71992, x37228);
  nand n37235(x37235, x25782, x84711);
  nand n37236(x37236, x37235, x37234);
  nand n37237(x37237, x25790, x84712);
  nand n37238(x37238, x71997, x37233);
  nand n37239(x37239, x25790, x37236);
  nand n37240(x37240, x37239, x37238);
  nand n37241(x37241, x72002, x84713);
  nand n37242(x37242, x25796, x37240);
  nand n37243(x37243, x37242, x37241);
  nand n37244(x37244, x71977, x27895);
  nand n37245(x37245, x16876, x36790);
  nand n37246(x37246, x37245, x26179);
  nand n37247(x37247, x71977, x84611);
  nand n37248(x37248, x16876, x35507);
  nand n37249(x37249, x71977, x28883);
  nand n37250(x37250, x16876, x28883);
  nand n37251(x37251, x37250, x37249);
  nand n37252(x37252, x71977, x36040);
  nand n37253(x37253, x16876, x36000);
  nand n37254(x37254, x37253, x37252);
  nand n37255(x37255, x71977, x29224);
  nand n37256(x37256, x37245, x37255);
  nand n37257(x37257, x16876, x28116);
  nand n37258(x37258, x37257, x37255);
  nand n37259(x37259, x71977, x35863);
  nand n37260(x37260, x25749, x84714);
  nand n37261(x37261, x71982, x37246);
  nand n37262(x37262, x25749, x84715);
  nand n37263(x37263, x37262, x37261);
  nand n37264(x37264, x71982, x84716);
  nand n37265(x37265, x25749, x37251);
  nand n37266(x37266, x37265, x37264);
  nand n37267(x37267, x71982, x37254);
  nand n37268(x37268, x25749, x37256);
  nand n37269(x37269, x37268, x37267);
  nand n37270(x37270, x71982, x84715);
  nand n37271(x37271, x25749, x84716);
  nand n37272(x37272, x37271, x37270);
  nand n37273(x37273, x71982, x37251);
  nand n37274(x37274, x25749, x37254);
  nand n37275(x37275, x37274, x37273);
  nand n37276(x37276, x71982, x37258);
  nand n37277(x37277, x25749, x84717);
  nand n37278(x37278, x37277, x37276);
  nand n37279(x37279, x71987, x84718);
  nand n37280(x37280, x25772, x37263);
  nand n37281(x37281, x37280, x26216);
  nand n37282(x37282, x71987, x37266);
  nand n37283(x37283, x25772, x37269);
  nand n37284(x37284, x37283, x37282);
  nand n37285(x37285, x71987, x37272);
  nand n37286(x37286, x25772, x37275);
  nand n37287(x37287, x37286, x37285);
  nand n37288(x37288, x71987, x37278);
  nand n37289(x37289, x25782, x84719);
  nand n37290(x37290, x71992, x37281);
  nand n37291(x37291, x25782, x37284);
  nand n37292(x37292, x37291, x37290);
  nand n37293(x37293, x71992, x37287);
  nand n37294(x37294, x25782, x84720);
  nand n37295(x37295, x37294, x37293);
  nand n37296(x37296, x25790, x84721);
  nand n37297(x37297, x71997, x37292);
  nand n37298(x37298, x25790, x37295);
  nand n37299(x37299, x37298, x37297);
  nand n37300(x37300, x72002, x84722);
  nand n37301(x37301, x25796, x37299);
  nand n37302(x37302, x37301, x37300);
  nand n37303(x37303, x71977, x27897);
  nand n37304(x37304, x16876, x36793);
  nand n37305(x37305, x37304, x26242);
  nand n37306(x37306, x71977, x84612);
  nand n37307(x37307, x16876, x35511);
  nand n37308(x37308, x71977, x28888);
  nand n37309(x37309, x16876, x28888);
  nand n37310(x37310, x37309, x37308);
  nand n37311(x37311, x71977, x36042);
  nand n37312(x37312, x16876, x36001);
  nand n37313(x37313, x37312, x37311);
  nand n37314(x37314, x71977, x29287);
  nand n37315(x37315, x37304, x37314);
  nand n37316(x37316, x16876, x28122);
  nand n37317(x37317, x37316, x37314);
  nand n37318(x37318, x71977, x35867);
  nand n37319(x37319, x25749, x84723);
  nand n37320(x37320, x71982, x37305);
  nand n37321(x37321, x25749, x84724);
  nand n37322(x37322, x37321, x37320);
  nand n37323(x37323, x71982, x84725);
  nand n37324(x37324, x25749, x37310);
  nand n37325(x37325, x37324, x37323);
  nand n37326(x37326, x71982, x37313);
  nand n37327(x37327, x25749, x37315);
  nand n37328(x37328, x37327, x37326);
  nand n37329(x37329, x71982, x84724);
  nand n37330(x37330, x25749, x84725);
  nand n37331(x37331, x37330, x37329);
  nand n37332(x37332, x71982, x37310);
  nand n37333(x37333, x25749, x37313);
  nand n37334(x37334, x37333, x37332);
  nand n37335(x37335, x71982, x37317);
  nand n37336(x37336, x25749, x84726);
  nand n37337(x37337, x37336, x37335);
  nand n37338(x37338, x71987, x84727);
  nand n37339(x37339, x25772, x37322);
  nand n37340(x37340, x37339, x26279);
  nand n37341(x37341, x71987, x37325);
  nand n37342(x37342, x25772, x37328);
  nand n37343(x37343, x37342, x37341);
  nand n37344(x37344, x71987, x37331);
  nand n37345(x37345, x25772, x37334);
  nand n37346(x37346, x37345, x37344);
  nand n37347(x37347, x71987, x37337);
  nand n37348(x37348, x25782, x84728);
  nand n37349(x37349, x71992, x37340);
  nand n37350(x37350, x25782, x37343);
  nand n37351(x37351, x37350, x37349);
  nand n37352(x37352, x71992, x37346);
  nand n37353(x37353, x25782, x84729);
  nand n37354(x37354, x37353, x37352);
  nand n37355(x37355, x25790, x84730);
  nand n37356(x37356, x71997, x37351);
  nand n37357(x37357, x25790, x37354);
  nand n37358(x37358, x37357, x37356);
  nand n37359(x37359, x72002, x84731);
  nand n37360(x37360, x25796, x37358);
  nand n37361(x37361, x37360, x37359);
  nand n37362(x37362, x71977, x27899);
  nand n37363(x37363, x16876, x36796);
  nand n37364(x37364, x37363, x26305);
  nand n37365(x37365, x71977, x84613);
  nand n37366(x37366, x16876, x35515);
  nand n37367(x37367, x71977, x28893);
  nand n37368(x37368, x16876, x28893);
  nand n37369(x37369, x37368, x37367);
  nand n37370(x37370, x71977, x36044);
  nand n37371(x37371, x16876, x36002);
  nand n37372(x37372, x37371, x37370);
  nand n37373(x37373, x71977, x29359);
  nand n37374(x37374, x37363, x37373);
  nand n37375(x37375, x16876, x28128);
  nand n37376(x37376, x37375, x37373);
  nand n37377(x37377, x71977, x35871);
  nand n37378(x37378, x25749, x84732);
  nand n37379(x37379, x71982, x37364);
  nand n37380(x37380, x25749, x84733);
  nand n37381(x37381, x37380, x37379);
  nand n37382(x37382, x71982, x84734);
  nand n37383(x37383, x25749, x37369);
  nand n37384(x37384, x37383, x37382);
  nand n37385(x37385, x71982, x37372);
  nand n37386(x37386, x25749, x37374);
  nand n37387(x37387, x37386, x37385);
  nand n37388(x37388, x71982, x84733);
  nand n37389(x37389, x25749, x84734);
  nand n37390(x37390, x37389, x37388);
  nand n37391(x37391, x71982, x37369);
  nand n37392(x37392, x25749, x37372);
  nand n37393(x37393, x37392, x37391);
  nand n37394(x37394, x71982, x37376);
  nand n37395(x37395, x25749, x84735);
  nand n37396(x37396, x37395, x37394);
  nand n37397(x37397, x71987, x84736);
  nand n37398(x37398, x25772, x37381);
  nand n37399(x37399, x37398, x26342);
  nand n37400(x37400, x71987, x37384);
  nand n37401(x37401, x25772, x37387);
  nand n37402(x37402, x37401, x37400);
  nand n37403(x37403, x71987, x37390);
  nand n37404(x37404, x25772, x37393);
  nand n37405(x37405, x37404, x37403);
  nand n37406(x37406, x71987, x37396);
  nand n37407(x37407, x25782, x84737);
  nand n37408(x37408, x71992, x37399);
  nand n37409(x37409, x25782, x37402);
  nand n37410(x37410, x37409, x37408);
  nand n37411(x37411, x71992, x37405);
  nand n37412(x37412, x25782, x84738);
  nand n37413(x37413, x37412, x37411);
  nand n37414(x37414, x25790, x84739);
  nand n37415(x37415, x71997, x37410);
  nand n37416(x37416, x25790, x37413);
  nand n37417(x37417, x37416, x37415);
  nand n37418(x37418, x72002, x84740);
  nand n37419(x37419, x25796, x37417);
  nand n37420(x37420, x37419, x37418);
  nand n37421(x37421, x71977, x27901);
  nand n37422(x37422, x16876, x36799);
  nand n37423(x37423, x37422, x26368);
  nand n37424(x37424, x71977, x84614);
  nand n37425(x37425, x16876, x35519);
  nand n37426(x37426, x71977, x28898);
  nand n37427(x37427, x16876, x28898);
  nand n37428(x37428, x37427, x37426);
  nand n37429(x37429, x71977, x36046);
  nand n37430(x37430, x16876, x36003);
  nand n37431(x37431, x37430, x37429);
  nand n37432(x37432, x71977, x29438);
  nand n37433(x37433, x37422, x37432);
  nand n37434(x37434, x16876, x28134);
  nand n37435(x37435, x37434, x37432);
  nand n37436(x37436, x71977, x35875);
  nand n37437(x37437, x25749, x84741);
  nand n37438(x37438, x71982, x37423);
  nand n37439(x37439, x25749, x84742);
  nand n37440(x37440, x37439, x37438);
  nand n37441(x37441, x71982, x84743);
  nand n37442(x37442, x25749, x37428);
  nand n37443(x37443, x37442, x37441);
  nand n37444(x37444, x71982, x37431);
  nand n37445(x37445, x25749, x37433);
  nand n37446(x37446, x37445, x37444);
  nand n37447(x37447, x71982, x84742);
  nand n37448(x37448, x25749, x84743);
  nand n37449(x37449, x37448, x37447);
  nand n37450(x37450, x71982, x37428);
  nand n37451(x37451, x25749, x37431);
  nand n37452(x37452, x37451, x37450);
  nand n37453(x37453, x71982, x37435);
  nand n37454(x37454, x25749, x84744);
  nand n37455(x37455, x37454, x37453);
  nand n37456(x37456, x71987, x84745);
  nand n37457(x37457, x25772, x37440);
  nand n37458(x37458, x37457, x26405);
  nand n37459(x37459, x71987, x37443);
  nand n37460(x37460, x25772, x37446);
  nand n37461(x37461, x37460, x37459);
  nand n37462(x37462, x71987, x37449);
  nand n37463(x37463, x25772, x37452);
  nand n37464(x37464, x37463, x37462);
  nand n37465(x37465, x71987, x37455);
  nand n37466(x37466, x25782, x84746);
  nand n37467(x37467, x71992, x37458);
  nand n37468(x37468, x25782, x37461);
  nand n37469(x37469, x37468, x37467);
  nand n37470(x37470, x71992, x37464);
  nand n37471(x37471, x25782, x84747);
  nand n37472(x37472, x37471, x37470);
  nand n37473(x37473, x25790, x84748);
  nand n37474(x37474, x71997, x37469);
  nand n37475(x37475, x25790, x37472);
  nand n37476(x37476, x37475, x37474);
  nand n37477(x37477, x72002, x84749);
  nand n37478(x37478, x25796, x37476);
  nand n37479(x37479, x37478, x37477);
  nand n37480(x37480, x71977, x27903);
  nand n37481(x37481, x16876, x36802);
  nand n37482(x37482, x37481, x26431);
  nand n37483(x37483, x71977, x84615);
  nand n37484(x37484, x16876, x35523);
  nand n37485(x37485, x71977, x28903);
  nand n37486(x37486, x16876, x28903);
  nand n37487(x37487, x37486, x37485);
  nand n37488(x37488, x71977, x36048);
  nand n37489(x37489, x16876, x36004);
  nand n37490(x37490, x37489, x37488);
  nand n37491(x37491, x71977, x29525);
  nand n37492(x37492, x37481, x37491);
  nand n37493(x37493, x16876, x28140);
  nand n37494(x37494, x37493, x37491);
  nand n37495(x37495, x71977, x35879);
  nand n37496(x37496, x25749, x84750);
  nand n37497(x37497, x71982, x37482);
  nand n37498(x37498, x25749, x84751);
  nand n37499(x37499, x37498, x37497);
  nand n37500(x37500, x71982, x84752);
  nand n37501(x37501, x25749, x37487);
  nand n37502(x37502, x37501, x37500);
  nand n37503(x37503, x71982, x37490);
  nand n37504(x37504, x25749, x37492);
  nand n37505(x37505, x37504, x37503);
  nand n37506(x37506, x71982, x84751);
  nand n37507(x37507, x25749, x84752);
  nand n37508(x37508, x37507, x37506);
  nand n37509(x37509, x71982, x37487);
  nand n37510(x37510, x25749, x37490);
  nand n37511(x37511, x37510, x37509);
  nand n37512(x37512, x71982, x37494);
  nand n37513(x37513, x25749, x84753);
  nand n37514(x37514, x37513, x37512);
  nand n37515(x37515, x71987, x84754);
  nand n37516(x37516, x25772, x37499);
  nand n37517(x37517, x37516, x26468);
  nand n37518(x37518, x71987, x37502);
  nand n37519(x37519, x25772, x37505);
  nand n37520(x37520, x37519, x37518);
  nand n37521(x37521, x71987, x37508);
  nand n37522(x37522, x25772, x37511);
  nand n37523(x37523, x37522, x37521);
  nand n37524(x37524, x71987, x37514);
  nand n37525(x37525, x25782, x84755);
  nand n37526(x37526, x71992, x37517);
  nand n37527(x37527, x25782, x37520);
  nand n37528(x37528, x37527, x37526);
  nand n37529(x37529, x71992, x37523);
  nand n37530(x37530, x25782, x84756);
  nand n37531(x37531, x37530, x37529);
  nand n37532(x37532, x25790, x84757);
  nand n37533(x37533, x71997, x37528);
  nand n37534(x37534, x25790, x37531);
  nand n37535(x37535, x37534, x37533);
  nand n37536(x37536, x72002, x84758);
  nand n37537(x37537, x25796, x37535);
  nand n37538(x37538, x37537, x37536);
  nand n37539(x37539, x71977, x27905);
  nand n37540(x37540, x16876, x36805);
  nand n37541(x37541, x37540, x26494);
  nand n37542(x37542, x71977, x84616);
  nand n37543(x37543, x16876, x35527);
  nand n37544(x37544, x71977, x28908);
  nand n37545(x37545, x16876, x28908);
  nand n37546(x37546, x37545, x37544);
  nand n37547(x37547, x71977, x36050);
  nand n37548(x37548, x16876, x36005);
  nand n37549(x37549, x37548, x37547);
  nand n37550(x37550, x71977, x29621);
  nand n37551(x37551, x37540, x37550);
  nand n37552(x37552, x16876, x28146);
  nand n37553(x37553, x37552, x37550);
  nand n37554(x37554, x71977, x35883);
  nand n37555(x37555, x25749, x84759);
  nand n37556(x37556, x71982, x37541);
  nand n37557(x37557, x25749, x84760);
  nand n37558(x37558, x37557, x37556);
  nand n37559(x37559, x71982, x84761);
  nand n37560(x37560, x25749, x37546);
  nand n37561(x37561, x37560, x37559);
  nand n37562(x37562, x71982, x37549);
  nand n37563(x37563, x25749, x37551);
  nand n37564(x37564, x37563, x37562);
  nand n37565(x37565, x71982, x84760);
  nand n37566(x37566, x25749, x84761);
  nand n37567(x37567, x37566, x37565);
  nand n37568(x37568, x71982, x37546);
  nand n37569(x37569, x25749, x37549);
  nand n37570(x37570, x37569, x37568);
  nand n37571(x37571, x71982, x37553);
  nand n37572(x37572, x25749, x84762);
  nand n37573(x37573, x37572, x37571);
  nand n37574(x37574, x71987, x84763);
  nand n37575(x37575, x25772, x37558);
  nand n37576(x37576, x37575, x26531);
  nand n37577(x37577, x71987, x37561);
  nand n37578(x37578, x25772, x37564);
  nand n37579(x37579, x37578, x37577);
  nand n37580(x37580, x71987, x37567);
  nand n37581(x37581, x25772, x37570);
  nand n37582(x37582, x37581, x37580);
  nand n37583(x37583, x71987, x37573);
  nand n37584(x37584, x25782, x84764);
  nand n37585(x37585, x71992, x37576);
  nand n37586(x37586, x25782, x37579);
  nand n37587(x37587, x37586, x37585);
  nand n37588(x37588, x71992, x37582);
  nand n37589(x37589, x25782, x84765);
  nand n37590(x37590, x37589, x37588);
  nand n37591(x37591, x25790, x84766);
  nand n37592(x37592, x71997, x37587);
  nand n37593(x37593, x25790, x37590);
  nand n37594(x37594, x37593, x37592);
  nand n37595(x37595, x72002, x84767);
  nand n37596(x37596, x25796, x37594);
  nand n37597(x37597, x37596, x37595);
  nand n37598(x37598, x71977, x27907);
  nand n37599(x37599, x16876, x36808);
  nand n37600(x37600, x37599, x26557);
  nand n37601(x37601, x71977, x84617);
  nand n37602(x37602, x16876, x35531);
  nand n37603(x37603, x71977, x28913);
  nand n37604(x37604, x16876, x28913);
  nand n37605(x37605, x37604, x37603);
  nand n37606(x37606, x71977, x36052);
  nand n37607(x37607, x16876, x36006);
  nand n37608(x37608, x37607, x37606);
  nand n37609(x37609, x71977, x29724);
  nand n37610(x37610, x37599, x37609);
  nand n37611(x37611, x16876, x28152);
  nand n37612(x37612, x37611, x37609);
  nand n37613(x37613, x71977, x35887);
  nand n37614(x37614, x25749, x84768);
  nand n37615(x37615, x71982, x37600);
  nand n37616(x37616, x25749, x84769);
  nand n37617(x37617, x37616, x37615);
  nand n37618(x37618, x71982, x84770);
  nand n37619(x37619, x25749, x37605);
  nand n37620(x37620, x37619, x37618);
  nand n37621(x37621, x71982, x37608);
  nand n37622(x37622, x25749, x37610);
  nand n37623(x37623, x37622, x37621);
  nand n37624(x37624, x71982, x84769);
  nand n37625(x37625, x25749, x84770);
  nand n37626(x37626, x37625, x37624);
  nand n37627(x37627, x71982, x37605);
  nand n37628(x37628, x25749, x37608);
  nand n37629(x37629, x37628, x37627);
  nand n37630(x37630, x71982, x37612);
  nand n37631(x37631, x25749, x84771);
  nand n37632(x37632, x37631, x37630);
  nand n37633(x37633, x71987, x84772);
  nand n37634(x37634, x25772, x37617);
  nand n37635(x37635, x37634, x26594);
  nand n37636(x37636, x71987, x37620);
  nand n37637(x37637, x25772, x37623);
  nand n37638(x37638, x37637, x37636);
  nand n37639(x37639, x71987, x37626);
  nand n37640(x37640, x25772, x37629);
  nand n37641(x37641, x37640, x37639);
  nand n37642(x37642, x71987, x37632);
  nand n37643(x37643, x25782, x84773);
  nand n37644(x37644, x71992, x37635);
  nand n37645(x37645, x25782, x37638);
  nand n37646(x37646, x37645, x37644);
  nand n37647(x37647, x71992, x37641);
  nand n37648(x37648, x25782, x84774);
  nand n37649(x37649, x37648, x37647);
  nand n37650(x37650, x25790, x84775);
  nand n37651(x37651, x71997, x37646);
  nand n37652(x37652, x25790, x37649);
  nand n37653(x37653, x37652, x37651);
  nand n37654(x37654, x72002, x84776);
  nand n37655(x37655, x25796, x37653);
  nand n37656(x37656, x37655, x37654);
  nand n37657(x37657, x71977, x27909);
  nand n37658(x37658, x16876, x36811);
  nand n37659(x37659, x37658, x26620);
  nand n37660(x37660, x71977, x84618);
  nand n37661(x37661, x16876, x35536);
  nand n37662(x37662, x71977, x28918);
  nand n37663(x37663, x16876, x28918);
  nand n37664(x37664, x37663, x37662);
  nand n37665(x37665, x71977, x36054);
  nand n37666(x37666, x16876, x36007);
  nand n37667(x37667, x37666, x37665);
  nand n37668(x37668, x71977, x29835);
  nand n37669(x37669, x37658, x37668);
  nand n37670(x37670, x16876, x28158);
  nand n37671(x37671, x37670, x37668);
  nand n37672(x37672, x71977, x35891);
  nand n37673(x37673, x25749, x84777);
  nand n37674(x37674, x71982, x37659);
  nand n37675(x37675, x25749, x84778);
  nand n37676(x37676, x37675, x37674);
  nand n37677(x37677, x71982, x84779);
  nand n37678(x37678, x25749, x37664);
  nand n37679(x37679, x37678, x37677);
  nand n37680(x37680, x71982, x37667);
  nand n37681(x37681, x25749, x37669);
  nand n37682(x37682, x37681, x37680);
  nand n37683(x37683, x71982, x84778);
  nand n37684(x37684, x25749, x84779);
  nand n37685(x37685, x37684, x37683);
  nand n37686(x37686, x71982, x37664);
  nand n37687(x37687, x25749, x37667);
  nand n37688(x37688, x37687, x37686);
  nand n37689(x37689, x71982, x37671);
  nand n37690(x37690, x25749, x84780);
  nand n37691(x37691, x37690, x37689);
  nand n37692(x37692, x71987, x84781);
  nand n37693(x37693, x25772, x37676);
  nand n37694(x37694, x37693, x26657);
  nand n37695(x37695, x71987, x37679);
  nand n37696(x37696, x25772, x37682);
  nand n37697(x37697, x37696, x37695);
  nand n37698(x37698, x71987, x37685);
  nand n37699(x37699, x25772, x37688);
  nand n37700(x37700, x37699, x37698);
  nand n37701(x37701, x71987, x37691);
  nand n37702(x37702, x25782, x84782);
  nand n37703(x37703, x71992, x37694);
  nand n37704(x37704, x25782, x37697);
  nand n37705(x37705, x37704, x37703);
  nand n37706(x37706, x71992, x37700);
  nand n37707(x37707, x25782, x84783);
  nand n37708(x37708, x37707, x37706);
  nand n37709(x37709, x25790, x84784);
  nand n37710(x37710, x71997, x37705);
  nand n37711(x37711, x25790, x37708);
  nand n37712(x37712, x37711, x37710);
  nand n37713(x37713, x72002, x84785);
  nand n37714(x37714, x25796, x37712);
  nand n37715(x37715, x37714, x37713);
  nand n37716(x37716, x71977, x27911);
  nand n37717(x37717, x16876, x36814);
  nand n37718(x37718, x37717, x26683);
  nand n37719(x37719, x71977, x84619);
  nand n37720(x37720, x16876, x35541);
  nand n37721(x37721, x71977, x28923);
  nand n37722(x37722, x16876, x28923);
  nand n37723(x37723, x37722, x37721);
  nand n37724(x37724, x71977, x36056);
  nand n37725(x37725, x16876, x36008);
  nand n37726(x37726, x37725, x37724);
  nand n37727(x37727, x71977, x29955);
  nand n37728(x37728, x37717, x37727);
  nand n37729(x37729, x16876, x28164);
  nand n37730(x37730, x37729, x37727);
  nand n37731(x37731, x71977, x35895);
  nand n37732(x37732, x25749, x84786);
  nand n37733(x37733, x71982, x37718);
  nand n37734(x37734, x25749, x84787);
  nand n37735(x37735, x37734, x37733);
  nand n37736(x37736, x71982, x84788);
  nand n37737(x37737, x25749, x37723);
  nand n37738(x37738, x37737, x37736);
  nand n37739(x37739, x71982, x37726);
  nand n37740(x37740, x25749, x37728);
  nand n37741(x37741, x37740, x37739);
  nand n37742(x37742, x71982, x84787);
  nand n37743(x37743, x25749, x84788);
  nand n37744(x37744, x37743, x37742);
  nand n37745(x37745, x71982, x37723);
  nand n37746(x37746, x25749, x37726);
  nand n37747(x37747, x37746, x37745);
  nand n37748(x37748, x71982, x37730);
  nand n37749(x37749, x25749, x84789);
  nand n37750(x37750, x37749, x37748);
  nand n37751(x37751, x71987, x84790);
  nand n37752(x37752, x25772, x37735);
  nand n37753(x37753, x37752, x26720);
  nand n37754(x37754, x71987, x37738);
  nand n37755(x37755, x25772, x37741);
  nand n37756(x37756, x37755, x37754);
  nand n37757(x37757, x71987, x37744);
  nand n37758(x37758, x25772, x37747);
  nand n37759(x37759, x37758, x37757);
  nand n37760(x37760, x71987, x37750);
  nand n37761(x37761, x25782, x84791);
  nand n37762(x37762, x71992, x37753);
  nand n37763(x37763, x25782, x37756);
  nand n37764(x37764, x37763, x37762);
  nand n37765(x37765, x71992, x37759);
  nand n37766(x37766, x25782, x84792);
  nand n37767(x37767, x37766, x37765);
  nand n37768(x37768, x25790, x84793);
  nand n37769(x37769, x71997, x37764);
  nand n37770(x37770, x25790, x37767);
  nand n37771(x37771, x37770, x37769);
  nand n37772(x37772, x72002, x84794);
  nand n37773(x37773, x25796, x37771);
  nand n37774(x37774, x37773, x37772);
  nand n37775(x37775, x71977, x27913);
  nand n37776(x37776, x16876, x84635);
  nand n37777(x37777, x37776, x26746);
  nand n37778(x37778, x71977, x36430);
  nand n37779(x37779, x16876, x35545);
  nand n37780(x37780, x71977, x28928);
  nand n37781(x37781, x16876, x28928);
  nand n37782(x37782, x37781, x37780);
  nand n37783(x37783, x71977, x36058);
  nand n37784(x37784, x16876, x36009);
  nand n37785(x37785, x37784, x37783);
  nand n37786(x37786, x71977, x35962);
  nand n37787(x37787, x37776, x37786);
  nand n37788(x37788, x16876, x28170);
  nand n37789(x37789, x37788, x37786);
  nand n37790(x37790, x71977, x35899);
  nand n37791(x37791, x25749, x84795);
  nand n37792(x37792, x71982, x37777);
  nand n37793(x37793, x25749, x84796);
  nand n37794(x37794, x37793, x37792);
  nand n37795(x37795, x71982, x84797);
  nand n37796(x37796, x25749, x37782);
  nand n37797(x37797, x37796, x37795);
  nand n37798(x37798, x71982, x37785);
  nand n37799(x37799, x25749, x37787);
  nand n37800(x37800, x37799, x37798);
  nand n37801(x37801, x71982, x84796);
  nand n37802(x37802, x25749, x84797);
  nand n37803(x37803, x37802, x37801);
  nand n37804(x37804, x71982, x37782);
  nand n37805(x37805, x25749, x37785);
  nand n37806(x37806, x37805, x37804);
  nand n37807(x37807, x71982, x37789);
  nand n37808(x37808, x25749, x84798);
  nand n37809(x37809, x37808, x37807);
  nand n37810(x37810, x71987, x84799);
  nand n37811(x37811, x25772, x37794);
  nand n37812(x37812, x37811, x26783);
  nand n37813(x37813, x71987, x37797);
  nand n37814(x37814, x25772, x37800);
  nand n37815(x37815, x37814, x37813);
  nand n37816(x37816, x71987, x37803);
  nand n37817(x37817, x25772, x37806);
  nand n37818(x37818, x37817, x37816);
  nand n37819(x37819, x71987, x37809);
  nand n37820(x37820, x25782, x84800);
  nand n37821(x37821, x71992, x37812);
  nand n37822(x37822, x25782, x37815);
  nand n37823(x37823, x37822, x37821);
  nand n37824(x37824, x71992, x37818);
  nand n37825(x37825, x25782, x84801);
  nand n37826(x37826, x37825, x37824);
  nand n37827(x37827, x25790, x84802);
  nand n37828(x37828, x71997, x37823);
  nand n37829(x37829, x25790, x37826);
  nand n37830(x37830, x37829, x37828);
  nand n37831(x37831, x72002, x84803);
  nand n37832(x37832, x25796, x37830);
  nand n37833(x37833, x37832, x37831);
  nand n37834(x37834, x71977, x27915);
  nand n37835(x37835, x16876, x84636);
  nand n37836(x37836, x37835, x26809);
  nand n37837(x37837, x71977, x36433);
  nand n37838(x37838, x16876, x35549);
  nand n37839(x37839, x71977, x28933);
  nand n37840(x37840, x16876, x28933);
  nand n37841(x37841, x37840, x37839);
  nand n37842(x37842, x71977, x36060);
  nand n37843(x37843, x16876, x36010);
  nand n37844(x37844, x37843, x37842);
  nand n37845(x37845, x71977, x35964);
  nand n37846(x37846, x37835, x37845);
  nand n37847(x37847, x16876, x28176);
  nand n37848(x37848, x37847, x37845);
  nand n37849(x37849, x71977, x35903);
  nand n37850(x37850, x25749, x84804);
  nand n37851(x37851, x71982, x37836);
  nand n37852(x37852, x25749, x84805);
  nand n37853(x37853, x37852, x37851);
  nand n37854(x37854, x71982, x84806);
  nand n37855(x37855, x25749, x37841);
  nand n37856(x37856, x37855, x37854);
  nand n37857(x37857, x71982, x37844);
  nand n37858(x37858, x25749, x37846);
  nand n37859(x37859, x37858, x37857);
  nand n37860(x37860, x71982, x84805);
  nand n37861(x37861, x25749, x84806);
  nand n37862(x37862, x37861, x37860);
  nand n37863(x37863, x71982, x37841);
  nand n37864(x37864, x25749, x37844);
  nand n37865(x37865, x37864, x37863);
  nand n37866(x37866, x71982, x37848);
  nand n37867(x37867, x25749, x84807);
  nand n37868(x37868, x37867, x37866);
  nand n37869(x37869, x71987, x84808);
  nand n37870(x37870, x25772, x37853);
  nand n37871(x37871, x37870, x26846);
  nand n37872(x37872, x71987, x37856);
  nand n37873(x37873, x25772, x37859);
  nand n37874(x37874, x37873, x37872);
  nand n37875(x37875, x71987, x37862);
  nand n37876(x37876, x25772, x37865);
  nand n37877(x37877, x37876, x37875);
  nand n37878(x37878, x71987, x37868);
  nand n37879(x37879, x25782, x84809);
  nand n37880(x37880, x71992, x37871);
  nand n37881(x37881, x25782, x37874);
  nand n37882(x37882, x37881, x37880);
  nand n37883(x37883, x71992, x37877);
  nand n37884(x37884, x25782, x84810);
  nand n37885(x37885, x37884, x37883);
  nand n37886(x37886, x25790, x84811);
  nand n37887(x37887, x71997, x37882);
  nand n37888(x37888, x25790, x37885);
  nand n37889(x37889, x37888, x37887);
  nand n37890(x37890, x72002, x84812);
  nand n37891(x37891, x25796, x37889);
  nand n37892(x37892, x37891, x37890);
  nand n37893(x37893, x71977, x27917);
  nand n37894(x37894, x16876, x84637);
  nand n37895(x37895, x37894, x26872);
  nand n37896(x37896, x71977, x36436);
  nand n37897(x37897, x16876, x35553);
  nand n37898(x37898, x71977, x28938);
  nand n37899(x37899, x16876, x28938);
  nand n37900(x37900, x37899, x37898);
  nand n37901(x37901, x71977, x36062);
  nand n37902(x37902, x16876, x36011);
  nand n37903(x37903, x37902, x37901);
  nand n37904(x37904, x71977, x35966);
  nand n37905(x37905, x37894, x37904);
  nand n37906(x37906, x16876, x28182);
  nand n37907(x37907, x37906, x37904);
  nand n37908(x37908, x71977, x35907);
  nand n37909(x37909, x25749, x84813);
  nand n37910(x37910, x71982, x37895);
  nand n37911(x37911, x25749, x84814);
  nand n37912(x37912, x37911, x37910);
  nand n37913(x37913, x71982, x84815);
  nand n37914(x37914, x25749, x37900);
  nand n37915(x37915, x37914, x37913);
  nand n37916(x37916, x71982, x37903);
  nand n37917(x37917, x25749, x37905);
  nand n37918(x37918, x37917, x37916);
  nand n37919(x37919, x71982, x84814);
  nand n37920(x37920, x25749, x84815);
  nand n37921(x37921, x37920, x37919);
  nand n37922(x37922, x71982, x37900);
  nand n37923(x37923, x25749, x37903);
  nand n37924(x37924, x37923, x37922);
  nand n37925(x37925, x71982, x37907);
  nand n37926(x37926, x25749, x84816);
  nand n37927(x37927, x37926, x37925);
  nand n37928(x37928, x71987, x84817);
  nand n37929(x37929, x25772, x37912);
  nand n37930(x37930, x37929, x26909);
  nand n37931(x37931, x71987, x37915);
  nand n37932(x37932, x25772, x37918);
  nand n37933(x37933, x37932, x37931);
  nand n37934(x37934, x71987, x37921);
  nand n37935(x37935, x25772, x37924);
  nand n37936(x37936, x37935, x37934);
  nand n37937(x37937, x71987, x37927);
  nand n37938(x37938, x25782, x84818);
  nand n37939(x37939, x71992, x37930);
  nand n37940(x37940, x25782, x37933);
  nand n37941(x37941, x37940, x37939);
  nand n37942(x37942, x71992, x37936);
  nand n37943(x37943, x25782, x84819);
  nand n37944(x37944, x37943, x37942);
  nand n37945(x37945, x25790, x84820);
  nand n37946(x37946, x71997, x37941);
  nand n37947(x37947, x25790, x37944);
  nand n37948(x37948, x37947, x37946);
  nand n37949(x37949, x72002, x84821);
  nand n37950(x37950, x25796, x37948);
  nand n37951(x37951, x37950, x37949);
  nand n37952(x37952, x71977, x27919);
  nand n37953(x37953, x16876, x84638);
  nand n37954(x37954, x37953, x26935);
  nand n37955(x37955, x71977, x36439);
  nand n37956(x37956, x16876, x35557);
  nand n37957(x37957, x71977, x28943);
  nand n37958(x37958, x16876, x28943);
  nand n37959(x37959, x37958, x37957);
  nand n37960(x37960, x71977, x36064);
  nand n37961(x37961, x16876, x36012);
  nand n37962(x37962, x37961, x37960);
  nand n37963(x37963, x71977, x35968);
  nand n37964(x37964, x37953, x37963);
  nand n37965(x37965, x16876, x28188);
  nand n37966(x37966, x37965, x37963);
  nand n37967(x37967, x71977, x35911);
  nand n37968(x37968, x25749, x84822);
  nand n37969(x37969, x71982, x37954);
  nand n37970(x37970, x25749, x84823);
  nand n37971(x37971, x37970, x37969);
  nand n37972(x37972, x71982, x84824);
  nand n37973(x37973, x25749, x37959);
  nand n37974(x37974, x37973, x37972);
  nand n37975(x37975, x71982, x37962);
  nand n37976(x37976, x25749, x37964);
  nand n37977(x37977, x37976, x37975);
  nand n37978(x37978, x71982, x84823);
  nand n37979(x37979, x25749, x84824);
  nand n37980(x37980, x37979, x37978);
  nand n37981(x37981, x71982, x37959);
  nand n37982(x37982, x25749, x37962);
  nand n37983(x37983, x37982, x37981);
  nand n37984(x37984, x71982, x37966);
  nand n37985(x37985, x25749, x84825);
  nand n37986(x37986, x37985, x37984);
  nand n37987(x37987, x71987, x84826);
  nand n37988(x37988, x25772, x37971);
  nand n37989(x37989, x37988, x26972);
  nand n37990(x37990, x71987, x37974);
  nand n37991(x37991, x25772, x37977);
  nand n37992(x37992, x37991, x37990);
  nand n37993(x37993, x71987, x37980);
  nand n37994(x37994, x25772, x37983);
  nand n37995(x37995, x37994, x37993);
  nand n37996(x37996, x71987, x37986);
  nand n37997(x37997, x25782, x84827);
  nand n37998(x37998, x71992, x37989);
  nand n37999(x37999, x25782, x37992);
  nand n38000(x38000, x37999, x37998);
  nand n38001(x38001, x71992, x37995);
  nand n38002(x38002, x25782, x84828);
  nand n38003(x38003, x38002, x38001);
  nand n38004(x38004, x25790, x84829);
  nand n38005(x38005, x71997, x38000);
  nand n38006(x38006, x25790, x38003);
  nand n38007(x38007, x38006, x38005);
  nand n38008(x38008, x72002, x84830);
  nand n38009(x38009, x25796, x38007);
  nand n38010(x38010, x38009, x38008);
  nand n38011(x38011, x71977, x27921);
  nand n38012(x38012, x16876, x84639);
  nand n38013(x38013, x38012, x26998);
  nand n38014(x38014, x71977, x36442);
  nand n38015(x38015, x16876, x35561);
  nand n38016(x38016, x71977, x28948);
  nand n38017(x38017, x16876, x28948);
  nand n38018(x38018, x38017, x38016);
  nand n38019(x38019, x71977, x36066);
  nand n38020(x38020, x16876, x36013);
  nand n38021(x38021, x38020, x38019);
  nand n38022(x38022, x71977, x35970);
  nand n38023(x38023, x38012, x38022);
  nand n38024(x38024, x16876, x28194);
  nand n38025(x38025, x38024, x38022);
  nand n38026(x38026, x71977, x35915);
  nand n38027(x38027, x25749, x84831);
  nand n38028(x38028, x71982, x38013);
  nand n38029(x38029, x25749, x84832);
  nand n38030(x38030, x38029, x38028);
  nand n38031(x38031, x71982, x84833);
  nand n38032(x38032, x25749, x38018);
  nand n38033(x38033, x38032, x38031);
  nand n38034(x38034, x71982, x38021);
  nand n38035(x38035, x25749, x38023);
  nand n38036(x38036, x38035, x38034);
  nand n38037(x38037, x71982, x84832);
  nand n38038(x38038, x25749, x84833);
  nand n38039(x38039, x38038, x38037);
  nand n38040(x38040, x71982, x38018);
  nand n38041(x38041, x25749, x38021);
  nand n38042(x38042, x38041, x38040);
  nand n38043(x38043, x71982, x38025);
  nand n38044(x38044, x25749, x84834);
  nand n38045(x38045, x38044, x38043);
  nand n38046(x38046, x71987, x84835);
  nand n38047(x38047, x25772, x38030);
  nand n38048(x38048, x38047, x27035);
  nand n38049(x38049, x71987, x38033);
  nand n38050(x38050, x25772, x38036);
  nand n38051(x38051, x38050, x38049);
  nand n38052(x38052, x71987, x38039);
  nand n38053(x38053, x25772, x38042);
  nand n38054(x38054, x38053, x38052);
  nand n38055(x38055, x71987, x38045);
  nand n38056(x38056, x25782, x84836);
  nand n38057(x38057, x71992, x38048);
  nand n38058(x38058, x25782, x38051);
  nand n38059(x38059, x38058, x38057);
  nand n38060(x38060, x71992, x38054);
  nand n38061(x38061, x25782, x84837);
  nand n38062(x38062, x38061, x38060);
  nand n38063(x38063, x25790, x84838);
  nand n38064(x38064, x71997, x38059);
  nand n38065(x38065, x25790, x38062);
  nand n38066(x38066, x38065, x38064);
  nand n38067(x38067, x72002, x84839);
  nand n38068(x38068, x25796, x38066);
  nand n38069(x38069, x38068, x38067);
  nand n38070(x38070, x71977, x27923);
  nand n38071(x38071, x16876, x84640);
  nand n38072(x38072, x38071, x27061);
  nand n38073(x38073, x71977, x36445);
  nand n38074(x38074, x16876, x35565);
  nand n38075(x38075, x71977, x28953);
  nand n38076(x38076, x16876, x28953);
  nand n38077(x38077, x38076, x38075);
  nand n38078(x38078, x71977, x36068);
  nand n38079(x38079, x16876, x36014);
  nand n38080(x38080, x38079, x38078);
  nand n38081(x38081, x71977, x35972);
  nand n38082(x38082, x38071, x38081);
  nand n38083(x38083, x16876, x28200);
  nand n38084(x38084, x38083, x38081);
  nand n38085(x38085, x71977, x35919);
  nand n38086(x38086, x25749, x84840);
  nand n38087(x38087, x71982, x38072);
  nand n38088(x38088, x25749, x84841);
  nand n38089(x38089, x38088, x38087);
  nand n38090(x38090, x71982, x84842);
  nand n38091(x38091, x25749, x38077);
  nand n38092(x38092, x38091, x38090);
  nand n38093(x38093, x71982, x38080);
  nand n38094(x38094, x25749, x38082);
  nand n38095(x38095, x38094, x38093);
  nand n38096(x38096, x71982, x84841);
  nand n38097(x38097, x25749, x84842);
  nand n38098(x38098, x38097, x38096);
  nand n38099(x38099, x71982, x38077);
  nand n38100(x38100, x25749, x38080);
  nand n38101(x38101, x38100, x38099);
  nand n38102(x38102, x71982, x38084);
  nand n38103(x38103, x25749, x84843);
  nand n38104(x38104, x38103, x38102);
  nand n38105(x38105, x71987, x84844);
  nand n38106(x38106, x25772, x38089);
  nand n38107(x38107, x38106, x27098);
  nand n38108(x38108, x71987, x38092);
  nand n38109(x38109, x25772, x38095);
  nand n38110(x38110, x38109, x38108);
  nand n38111(x38111, x71987, x38098);
  nand n38112(x38112, x25772, x38101);
  nand n38113(x38113, x38112, x38111);
  nand n38114(x38114, x71987, x38104);
  nand n38115(x38115, x25782, x84845);
  nand n38116(x38116, x71992, x38107);
  nand n38117(x38117, x25782, x38110);
  nand n38118(x38118, x38117, x38116);
  nand n38119(x38119, x71992, x38113);
  nand n38120(x38120, x25782, x84846);
  nand n38121(x38121, x38120, x38119);
  nand n38122(x38122, x25790, x84847);
  nand n38123(x38123, x71997, x38118);
  nand n38124(x38124, x25790, x38121);
  nand n38125(x38125, x38124, x38123);
  nand n38126(x38126, x72002, x84848);
  nand n38127(x38127, x25796, x38125);
  nand n38128(x38128, x38127, x38126);
  nand n38129(x38129, x71977, x27925);
  nand n38130(x38130, x16876, x84641);
  nand n38131(x38131, x38130, x27124);
  nand n38132(x38132, x71977, x36448);
  nand n38133(x38133, x16876, x35570);
  nand n38134(x38134, x71977, x28958);
  nand n38135(x38135, x16876, x28958);
  nand n38136(x38136, x38135, x38134);
  nand n38137(x38137, x71977, x36070);
  nand n38138(x38138, x16876, x36015);
  nand n38139(x38139, x38138, x38137);
  nand n38140(x38140, x71977, x35974);
  nand n38141(x38141, x38130, x38140);
  nand n38142(x38142, x16876, x28206);
  nand n38143(x38143, x38142, x38140);
  nand n38144(x38144, x71977, x35923);
  nand n38145(x38145, x25749, x84849);
  nand n38146(x38146, x71982, x38131);
  nand n38147(x38147, x25749, x84850);
  nand n38148(x38148, x38147, x38146);
  nand n38149(x38149, x71982, x84851);
  nand n38150(x38150, x25749, x38136);
  nand n38151(x38151, x38150, x38149);
  nand n38152(x38152, x71982, x38139);
  nand n38153(x38153, x25749, x38141);
  nand n38154(x38154, x38153, x38152);
  nand n38155(x38155, x71982, x84850);
  nand n38156(x38156, x25749, x84851);
  nand n38157(x38157, x38156, x38155);
  nand n38158(x38158, x71982, x38136);
  nand n38159(x38159, x25749, x38139);
  nand n38160(x38160, x38159, x38158);
  nand n38161(x38161, x71982, x38143);
  nand n38162(x38162, x25749, x84852);
  nand n38163(x38163, x38162, x38161);
  nand n38164(x38164, x71987, x84853);
  nand n38165(x38165, x25772, x38148);
  nand n38166(x38166, x38165, x27161);
  nand n38167(x38167, x71987, x38151);
  nand n38168(x38168, x25772, x38154);
  nand n38169(x38169, x38168, x38167);
  nand n38170(x38170, x71987, x38157);
  nand n38171(x38171, x25772, x38160);
  nand n38172(x38172, x38171, x38170);
  nand n38173(x38173, x71987, x38163);
  nand n38174(x38174, x25782, x84854);
  nand n38175(x38175, x71992, x38166);
  nand n38176(x38176, x25782, x38169);
  nand n38177(x38177, x38176, x38175);
  nand n38178(x38178, x71992, x38172);
  nand n38179(x38179, x25782, x84855);
  nand n38180(x38180, x38179, x38178);
  nand n38181(x38181, x25790, x84856);
  nand n38182(x38182, x71997, x38177);
  nand n38183(x38183, x25790, x38180);
  nand n38184(x38184, x38183, x38182);
  nand n38185(x38185, x72002, x84857);
  nand n38186(x38186, x25796, x38184);
  nand n38187(x38187, x38186, x38185);
  nand n38188(x38188, x71977, x27927);
  nand n38189(x38189, x16876, x84642);
  nand n38190(x38190, x38189, x27187);
  nand n38191(x38191, x71977, x36451);
  nand n38192(x38192, x16876, x35575);
  nand n38193(x38193, x71977, x28963);
  nand n38194(x38194, x16876, x28963);
  nand n38195(x38195, x38194, x38193);
  nand n38196(x38196, x71977, x36072);
  nand n38197(x38197, x16876, x36016);
  nand n38198(x38198, x38197, x38196);
  nand n38199(x38199, x71977, x35976);
  nand n38200(x38200, x38189, x38199);
  nand n38201(x38201, x16876, x28212);
  nand n38202(x38202, x38201, x38199);
  nand n38203(x38203, x71977, x35927);
  nand n38204(x38204, x25749, x84858);
  nand n38205(x38205, x71982, x38190);
  nand n38206(x38206, x25749, x84859);
  nand n38207(x38207, x38206, x38205);
  nand n38208(x38208, x71982, x84860);
  nand n38209(x38209, x25749, x38195);
  nand n38210(x38210, x38209, x38208);
  nand n38211(x38211, x71982, x38198);
  nand n38212(x38212, x25749, x38200);
  nand n38213(x38213, x38212, x38211);
  nand n38214(x38214, x71982, x84859);
  nand n38215(x38215, x25749, x84860);
  nand n38216(x38216, x38215, x38214);
  nand n38217(x38217, x71982, x38195);
  nand n38218(x38218, x25749, x38198);
  nand n38219(x38219, x38218, x38217);
  nand n38220(x38220, x71982, x38202);
  nand n38221(x38221, x25749, x84861);
  nand n38222(x38222, x38221, x38220);
  nand n38223(x38223, x71987, x84862);
  nand n38224(x38224, x25772, x38207);
  nand n38225(x38225, x38224, x27224);
  nand n38226(x38226, x71987, x38210);
  nand n38227(x38227, x25772, x38213);
  nand n38228(x38228, x38227, x38226);
  nand n38229(x38229, x71987, x38216);
  nand n38230(x38230, x25772, x38219);
  nand n38231(x38231, x38230, x38229);
  nand n38232(x38232, x71987, x38222);
  nand n38233(x38233, x25782, x84863);
  nand n38234(x38234, x71992, x38225);
  nand n38235(x38235, x25782, x38228);
  nand n38236(x38236, x38235, x38234);
  nand n38237(x38237, x71992, x38231);
  nand n38238(x38238, x25782, x84864);
  nand n38239(x38239, x38238, x38237);
  nand n38240(x38240, x25790, x84865);
  nand n38241(x38241, x71997, x38236);
  nand n38242(x38242, x25790, x38239);
  nand n38243(x38243, x38242, x38241);
  nand n38244(x38244, x72002, x84866);
  nand n38245(x38245, x25796, x38243);
  nand n38246(x38246, x38245, x38244);
  nand n38247(x38247, x71977, x27929);
  nand n38248(x38248, x16876, x84643);
  nand n38249(x38249, x38248, x27250);
  nand n38250(x38250, x71977, x36454);
  nand n38251(x38251, x16876, x35580);
  nand n38252(x38252, x71977, x28968);
  nand n38253(x38253, x16876, x28968);
  nand n38254(x38254, x38253, x38252);
  nand n38255(x38255, x71977, x36074);
  nand n38256(x38256, x16876, x36017);
  nand n38257(x38257, x38256, x38255);
  nand n38258(x38258, x71977, x35978);
  nand n38259(x38259, x38248, x38258);
  nand n38260(x38260, x16876, x28218);
  nand n38261(x38261, x38260, x38258);
  nand n38262(x38262, x71977, x35931);
  nand n38263(x38263, x25749, x84867);
  nand n38264(x38264, x71982, x38249);
  nand n38265(x38265, x25749, x84868);
  nand n38266(x38266, x38265, x38264);
  nand n38267(x38267, x71982, x84869);
  nand n38268(x38268, x25749, x38254);
  nand n38269(x38269, x38268, x38267);
  nand n38270(x38270, x71982, x38257);
  nand n38271(x38271, x25749, x38259);
  nand n38272(x38272, x38271, x38270);
  nand n38273(x38273, x71982, x84868);
  nand n38274(x38274, x25749, x84869);
  nand n38275(x38275, x38274, x38273);
  nand n38276(x38276, x71982, x38254);
  nand n38277(x38277, x25749, x38257);
  nand n38278(x38278, x38277, x38276);
  nand n38279(x38279, x71982, x38261);
  nand n38280(x38280, x25749, x84870);
  nand n38281(x38281, x38280, x38279);
  nand n38282(x38282, x71987, x84871);
  nand n38283(x38283, x25772, x38266);
  nand n38284(x38284, x38283, x27287);
  nand n38285(x38285, x71987, x38269);
  nand n38286(x38286, x25772, x38272);
  nand n38287(x38287, x38286, x38285);
  nand n38288(x38288, x71987, x38275);
  nand n38289(x38289, x25772, x38278);
  nand n38290(x38290, x38289, x38288);
  nand n38291(x38291, x71987, x38281);
  nand n38292(x38292, x25782, x84872);
  nand n38293(x38293, x71992, x38284);
  nand n38294(x38294, x25782, x38287);
  nand n38295(x38295, x38294, x38293);
  nand n38296(x38296, x71992, x38290);
  nand n38297(x38297, x25782, x84873);
  nand n38298(x38298, x38297, x38296);
  nand n38299(x38299, x25790, x84874);
  nand n38300(x38300, x71997, x38295);
  nand n38301(x38301, x25790, x38298);
  nand n38302(x38302, x38301, x38300);
  nand n38303(x38303, x72002, x84875);
  nand n38304(x38304, x25796, x38302);
  nand n38305(x38305, x38304, x38303);
  nand n38306(x38306, x71977, x27931);
  nand n38307(x38307, x16876, x84644);
  nand n38308(x38308, x38307, x27313);
  nand n38309(x38309, x71977, x36457);
  nand n38310(x38310, x16876, x35585);
  nand n38311(x38311, x71977, x28973);
  nand n38312(x38312, x16876, x28973);
  nand n38313(x38313, x38312, x38311);
  nand n38314(x38314, x71977, x36076);
  nand n38315(x38315, x16876, x36018);
  nand n38316(x38316, x38315, x38314);
  nand n38317(x38317, x71977, x35980);
  nand n38318(x38318, x38307, x38317);
  nand n38319(x38319, x16876, x28224);
  nand n38320(x38320, x38319, x38317);
  nand n38321(x38321, x71977, x35935);
  nand n38322(x38322, x25749, x84876);
  nand n38323(x38323, x71982, x38308);
  nand n38324(x38324, x25749, x84877);
  nand n38325(x38325, x38324, x38323);
  nand n38326(x38326, x71982, x84878);
  nand n38327(x38327, x25749, x38313);
  nand n38328(x38328, x38327, x38326);
  nand n38329(x38329, x71982, x38316);
  nand n38330(x38330, x25749, x38318);
  nand n38331(x38331, x38330, x38329);
  nand n38332(x38332, x71982, x84877);
  nand n38333(x38333, x25749, x84878);
  nand n38334(x38334, x38333, x38332);
  nand n38335(x38335, x71982, x38313);
  nand n38336(x38336, x25749, x38316);
  nand n38337(x38337, x38336, x38335);
  nand n38338(x38338, x71982, x38320);
  nand n38339(x38339, x25749, x84879);
  nand n38340(x38340, x38339, x38338);
  nand n38341(x38341, x71987, x84880);
  nand n38342(x38342, x25772, x38325);
  nand n38343(x38343, x38342, x27350);
  nand n38344(x38344, x71987, x38328);
  nand n38345(x38345, x25772, x38331);
  nand n38346(x38346, x38345, x38344);
  nand n38347(x38347, x71987, x38334);
  nand n38348(x38348, x25772, x38337);
  nand n38349(x38349, x38348, x38347);
  nand n38350(x38350, x71987, x38340);
  nand n38351(x38351, x25782, x84881);
  nand n38352(x38352, x71992, x38343);
  nand n38353(x38353, x25782, x38346);
  nand n38354(x38354, x38353, x38352);
  nand n38355(x38355, x71992, x38349);
  nand n38356(x38356, x25782, x84882);
  nand n38357(x38357, x38356, x38355);
  nand n38358(x38358, x25790, x84883);
  nand n38359(x38359, x71997, x38354);
  nand n38360(x38360, x25790, x38357);
  nand n38361(x38361, x38360, x38359);
  nand n38362(x38362, x72002, x84884);
  nand n38363(x38363, x25796, x38361);
  nand n38364(x38364, x38363, x38362);
  nand n38365(x38365, x71977, x27933);
  nand n38366(x38366, x16876, x84645);
  nand n38367(x38367, x38366, x27376);
  nand n38368(x38368, x71977, x36460);
  nand n38369(x38369, x16876, x35590);
  nand n38370(x38370, x71977, x28978);
  nand n38371(x38371, x16876, x28978);
  nand n38372(x38372, x38371, x38370);
  nand n38373(x38373, x71977, x36078);
  nand n38374(x38374, x16876, x36019);
  nand n38375(x38375, x38374, x38373);
  nand n38376(x38376, x71977, x35982);
  nand n38377(x38377, x38366, x38376);
  nand n38378(x38378, x16876, x28230);
  nand n38379(x38379, x38378, x38376);
  nand n38380(x38380, x71977, x35939);
  nand n38381(x38381, x25749, x84885);
  nand n38382(x38382, x71982, x38367);
  nand n38383(x38383, x25749, x84886);
  nand n38384(x38384, x38383, x38382);
  nand n38385(x38385, x71982, x84887);
  nand n38386(x38386, x25749, x38372);
  nand n38387(x38387, x38386, x38385);
  nand n38388(x38388, x71982, x38375);
  nand n38389(x38389, x25749, x38377);
  nand n38390(x38390, x38389, x38388);
  nand n38391(x38391, x71982, x84886);
  nand n38392(x38392, x25749, x84887);
  nand n38393(x38393, x38392, x38391);
  nand n38394(x38394, x71982, x38372);
  nand n38395(x38395, x25749, x38375);
  nand n38396(x38396, x38395, x38394);
  nand n38397(x38397, x71982, x38379);
  nand n38398(x38398, x25749, x84888);
  nand n38399(x38399, x38398, x38397);
  nand n38400(x38400, x71987, x84889);
  nand n38401(x38401, x25772, x38384);
  nand n38402(x38402, x38401, x27413);
  nand n38403(x38403, x71987, x38387);
  nand n38404(x38404, x25772, x38390);
  nand n38405(x38405, x38404, x38403);
  nand n38406(x38406, x71987, x38393);
  nand n38407(x38407, x25772, x38396);
  nand n38408(x38408, x38407, x38406);
  nand n38409(x38409, x71987, x38399);
  nand n38410(x38410, x25782, x84890);
  nand n38411(x38411, x71992, x38402);
  nand n38412(x38412, x25782, x38405);
  nand n38413(x38413, x38412, x38411);
  nand n38414(x38414, x71992, x38408);
  nand n38415(x38415, x25782, x84891);
  nand n38416(x38416, x38415, x38414);
  nand n38417(x38417, x25790, x84892);
  nand n38418(x38418, x71997, x38413);
  nand n38419(x38419, x25790, x38416);
  nand n38420(x38420, x38419, x38418);
  nand n38421(x38421, x72002, x84893);
  nand n38422(x38422, x25796, x38420);
  nand n38423(x38423, x38422, x38421);
  nand n38424(x38424, x71977, x27935);
  nand n38425(x38425, x16876, x84646);
  nand n38426(x38426, x38425, x27439);
  nand n38427(x38427, x71977, x36463);
  nand n38428(x38428, x16876, x35595);
  nand n38429(x38429, x71977, x28983);
  nand n38430(x38430, x16876, x28983);
  nand n38431(x38431, x38430, x38429);
  nand n38432(x38432, x71977, x36080);
  nand n38433(x38433, x16876, x36020);
  nand n38434(x38434, x38433, x38432);
  nand n38435(x38435, x71977, x35984);
  nand n38436(x38436, x38425, x38435);
  nand n38437(x38437, x16876, x28236);
  nand n38438(x38438, x38437, x38435);
  nand n38439(x38439, x71977, x35943);
  nand n38440(x38440, x25749, x84894);
  nand n38441(x38441, x71982, x38426);
  nand n38442(x38442, x25749, x84895);
  nand n38443(x38443, x38442, x38441);
  nand n38444(x38444, x71982, x84896);
  nand n38445(x38445, x25749, x38431);
  nand n38446(x38446, x38445, x38444);
  nand n38447(x38447, x71982, x38434);
  nand n38448(x38448, x25749, x38436);
  nand n38449(x38449, x38448, x38447);
  nand n38450(x38450, x71982, x84895);
  nand n38451(x38451, x25749, x84896);
  nand n38452(x38452, x38451, x38450);
  nand n38453(x38453, x71982, x38431);
  nand n38454(x38454, x25749, x38434);
  nand n38455(x38455, x38454, x38453);
  nand n38456(x38456, x71982, x38438);
  nand n38457(x38457, x25749, x84897);
  nand n38458(x38458, x38457, x38456);
  nand n38459(x38459, x71987, x84898);
  nand n38460(x38460, x25772, x38443);
  nand n38461(x38461, x38460, x27476);
  nand n38462(x38462, x71987, x38446);
  nand n38463(x38463, x25772, x38449);
  nand n38464(x38464, x38463, x38462);
  nand n38465(x38465, x71987, x38452);
  nand n38466(x38466, x25772, x38455);
  nand n38467(x38467, x38466, x38465);
  nand n38468(x38468, x71987, x38458);
  nand n38469(x38469, x25782, x84899);
  nand n38470(x38470, x71992, x38461);
  nand n38471(x38471, x25782, x38464);
  nand n38472(x38472, x38471, x38470);
  nand n38473(x38473, x71992, x38467);
  nand n38474(x38474, x25782, x84900);
  nand n38475(x38475, x38474, x38473);
  nand n38476(x38476, x25790, x84901);
  nand n38477(x38477, x71997, x38472);
  nand n38478(x38478, x25790, x38475);
  nand n38479(x38479, x38478, x38477);
  nand n38480(x38480, x72002, x84902);
  nand n38481(x38481, x25796, x38479);
  nand n38482(x38482, x38481, x38480);
  nand n38483(x38483, x71977, x27937);
  nand n38484(x38484, x16876, x84647);
  nand n38485(x38485, x38484, x27502);
  nand n38486(x38486, x71977, x36466);
  nand n38487(x38487, x16876, x35600);
  nand n38488(x38488, x71977, x28988);
  nand n38489(x38489, x16876, x28988);
  nand n38490(x38490, x38489, x38488);
  nand n38491(x38491, x71977, x36082);
  nand n38492(x38492, x16876, x36021);
  nand n38493(x38493, x38492, x38491);
  nand n38494(x38494, x71977, x35986);
  nand n38495(x38495, x38484, x38494);
  nand n38496(x38496, x16876, x28242);
  nand n38497(x38497, x38496, x38494);
  nand n38498(x38498, x71977, x35947);
  nand n38499(x38499, x25749, x84903);
  nand n38500(x38500, x71982, x38485);
  nand n38501(x38501, x25749, x84904);
  nand n38502(x38502, x38501, x38500);
  nand n38503(x38503, x71982, x84905);
  nand n38504(x38504, x25749, x38490);
  nand n38505(x38505, x38504, x38503);
  nand n38506(x38506, x71982, x38493);
  nand n38507(x38507, x25749, x38495);
  nand n38508(x38508, x38507, x38506);
  nand n38509(x38509, x71982, x84904);
  nand n38510(x38510, x25749, x84905);
  nand n38511(x38511, x38510, x38509);
  nand n38512(x38512, x71982, x38490);
  nand n38513(x38513, x25749, x38493);
  nand n38514(x38514, x38513, x38512);
  nand n38515(x38515, x71982, x38497);
  nand n38516(x38516, x25749, x84906);
  nand n38517(x38517, x38516, x38515);
  nand n38518(x38518, x71987, x84907);
  nand n38519(x38519, x25772, x38502);
  nand n38520(x38520, x38519, x27539);
  nand n38521(x38521, x71987, x38505);
  nand n38522(x38522, x25772, x38508);
  nand n38523(x38523, x38522, x38521);
  nand n38524(x38524, x71987, x38511);
  nand n38525(x38525, x25772, x38514);
  nand n38526(x38526, x38525, x38524);
  nand n38527(x38527, x71987, x38517);
  nand n38528(x38528, x25782, x84908);
  nand n38529(x38529, x71992, x38520);
  nand n38530(x38530, x25782, x38523);
  nand n38531(x38531, x38530, x38529);
  nand n38532(x38532, x71992, x38526);
  nand n38533(x38533, x25782, x84909);
  nand n38534(x38534, x38533, x38532);
  nand n38535(x38535, x25790, x84910);
  nand n38536(x38536, x71997, x38531);
  nand n38537(x38537, x25790, x38534);
  nand n38538(x38538, x38537, x38536);
  nand n38539(x38539, x72002, x84911);
  nand n38540(x38540, x25796, x38538);
  nand n38541(x38541, x38540, x38539);
  nand n38542(x38542, x71977, x27939);
  nand n38543(x38543, x16876, x84648);
  nand n38544(x38544, x38543, x27565);
  nand n38545(x38545, x71977, x36469);
  nand n38546(x38546, x16876, x35605);
  nand n38547(x38547, x71977, x28993);
  nand n38548(x38548, x16876, x28993);
  nand n38549(x38549, x38548, x38547);
  nand n38550(x38550, x71977, x36084);
  nand n38551(x38551, x16876, x36022);
  nand n38552(x38552, x38551, x38550);
  nand n38553(x38553, x71977, x35988);
  nand n38554(x38554, x38543, x38553);
  nand n38555(x38555, x16876, x28248);
  nand n38556(x38556, x38555, x38553);
  nand n38557(x38557, x71977, x35951);
  nand n38558(x38558, x25749, x84912);
  nand n38559(x38559, x71982, x38544);
  nand n38560(x38560, x25749, x84913);
  nand n38561(x38561, x38560, x38559);
  nand n38562(x38562, x71982, x84914);
  nand n38563(x38563, x25749, x38549);
  nand n38564(x38564, x38563, x38562);
  nand n38565(x38565, x71982, x38552);
  nand n38566(x38566, x25749, x38554);
  nand n38567(x38567, x38566, x38565);
  nand n38568(x38568, x71982, x84913);
  nand n38569(x38569, x25749, x84914);
  nand n38570(x38570, x38569, x38568);
  nand n38571(x38571, x71982, x38549);
  nand n38572(x38572, x25749, x38552);
  nand n38573(x38573, x38572, x38571);
  nand n38574(x38574, x71982, x38556);
  nand n38575(x38575, x25749, x84915);
  nand n38576(x38576, x38575, x38574);
  nand n38577(x38577, x71987, x84916);
  nand n38578(x38578, x25772, x38561);
  nand n38579(x38579, x38578, x27602);
  nand n38580(x38580, x71987, x38564);
  nand n38581(x38581, x25772, x38567);
  nand n38582(x38582, x38581, x38580);
  nand n38583(x38583, x71987, x38570);
  nand n38584(x38584, x25772, x38573);
  nand n38585(x38585, x38584, x38583);
  nand n38586(x38586, x71987, x38576);
  nand n38587(x38587, x25782, x84917);
  nand n38588(x38588, x71992, x38579);
  nand n38589(x38589, x25782, x38582);
  nand n38590(x38590, x38589, x38588);
  nand n38591(x38591, x71992, x38585);
  nand n38592(x38592, x25782, x84918);
  nand n38593(x38593, x38592, x38591);
  nand n38594(x38594, x25790, x84919);
  nand n38595(x38595, x71997, x38590);
  nand n38596(x38596, x25790, x38593);
  nand n38597(x38597, x38596, x38595);
  nand n38598(x38598, x72002, x84920);
  nand n38599(x38599, x25796, x38597);
  nand n38600(x38600, x38599, x38598);
  nand n38601(x38601, x71977, x27941);
  nand n38602(x38602, x16876, x84649);
  nand n38603(x38603, x38602, x27628);
  nand n38604(x38604, x71977, x36472);
  nand n38605(x38605, x16876, x35610);
  nand n38606(x38606, x71977, x28998);
  nand n38607(x38607, x16876, x28998);
  nand n38608(x38608, x38607, x38606);
  nand n38609(x38609, x71977, x36086);
  nand n38610(x38610, x16876, x36023);
  nand n38611(x38611, x38610, x38609);
  nand n38612(x38612, x71977, x35990);
  nand n38613(x38613, x38602, x38612);
  nand n38614(x38614, x16876, x28254);
  nand n38615(x38615, x38614, x38612);
  nand n38616(x38616, x71977, x35955);
  nand n38617(x38617, x25749, x84921);
  nand n38618(x38618, x71982, x38603);
  nand n38619(x38619, x25749, x84922);
  nand n38620(x38620, x38619, x38618);
  nand n38621(x38621, x71982, x84923);
  nand n38622(x38622, x25749, x38608);
  nand n38623(x38623, x38622, x38621);
  nand n38624(x38624, x71982, x38611);
  nand n38625(x38625, x25749, x38613);
  nand n38626(x38626, x38625, x38624);
  nand n38627(x38627, x71982, x84922);
  nand n38628(x38628, x25749, x84923);
  nand n38629(x38629, x38628, x38627);
  nand n38630(x38630, x71982, x38608);
  nand n38631(x38631, x25749, x38611);
  nand n38632(x38632, x38631, x38630);
  nand n38633(x38633, x71982, x38615);
  nand n38634(x38634, x25749, x84924);
  nand n38635(x38635, x38634, x38633);
  nand n38636(x38636, x71987, x84925);
  nand n38637(x38637, x25772, x38620);
  nand n38638(x38638, x38637, x27665);
  nand n38639(x38639, x71987, x38623);
  nand n38640(x38640, x25772, x38626);
  nand n38641(x38641, x38640, x38639);
  nand n38642(x38642, x71987, x38629);
  nand n38643(x38643, x25772, x38632);
  nand n38644(x38644, x38643, x38642);
  nand n38645(x38645, x71987, x38635);
  nand n38646(x38646, x25782, x84926);
  nand n38647(x38647, x71992, x38638);
  nand n38648(x38648, x25782, x38641);
  nand n38649(x38649, x38648, x38647);
  nand n38650(x38650, x71992, x38644);
  nand n38651(x38651, x25782, x84927);
  nand n38652(x38652, x38651, x38650);
  nand n38653(x38653, x25790, x84928);
  nand n38654(x38654, x71997, x38649);
  nand n38655(x38655, x25790, x38652);
  nand n38656(x38656, x38655, x38654);
  nand n38657(x38657, x72002, x84929);
  nand n38658(x38658, x25796, x38656);
  nand n38659(x38659, x38658, x38657);
  nand n38660(x38660, x71977, x27943);
  nand n38661(x38661, x16876, x84650);
  nand n38662(x38662, x38661, x27691);
  nand n38663(x38663, x71977, x36475);
  nand n38664(x38664, x16876, x35615);
  nand n38665(x38665, x71977, x29003);
  nand n38666(x38666, x16876, x29003);
  nand n38667(x38667, x38666, x38665);
  nand n38668(x38668, x71977, x36088);
  nand n38669(x38669, x16876, x36024);
  nand n38670(x38670, x38669, x38668);
  nand n38671(x38671, x71977, x35992);
  nand n38672(x38672, x38661, x38671);
  nand n38673(x38673, x16876, x28260);
  nand n38674(x38674, x38673, x38671);
  nand n38675(x38675, x71977, x35959);
  nand n38676(x38676, x25749, x84930);
  nand n38677(x38677, x71982, x38662);
  nand n38678(x38678, x25749, x84931);
  nand n38679(x38679, x38678, x38677);
  nand n38680(x38680, x71982, x84932);
  nand n38681(x38681, x25749, x38667);
  nand n38682(x38682, x38681, x38680);
  nand n38683(x38683, x71982, x38670);
  nand n38684(x38684, x25749, x38672);
  nand n38685(x38685, x38684, x38683);
  nand n38686(x38686, x71982, x84931);
  nand n38687(x38687, x25749, x84932);
  nand n38688(x38688, x38687, x38686);
  nand n38689(x38689, x71982, x38667);
  nand n38690(x38690, x25749, x38670);
  nand n38691(x38691, x38690, x38689);
  nand n38692(x38692, x71982, x38674);
  nand n38693(x38693, x25749, x84933);
  nand n38694(x38694, x38693, x38692);
  nand n38695(x38695, x71987, x84934);
  nand n38696(x38696, x25772, x38679);
  nand n38697(x38697, x38696, x27728);
  nand n38698(x38698, x71987, x38682);
  nand n38699(x38699, x25772, x38685);
  nand n38700(x38700, x38699, x38698);
  nand n38701(x38701, x71987, x38688);
  nand n38702(x38702, x25772, x38691);
  nand n38703(x38703, x38702, x38701);
  nand n38704(x38704, x71987, x38694);
  nand n38705(x38705, x25782, x84935);
  nand n38706(x38706, x71992, x38697);
  nand n38707(x38707, x25782, x38700);
  nand n38708(x38708, x38707, x38706);
  nand n38709(x38709, x71992, x38703);
  nand n38710(x38710, x25782, x84936);
  nand n38711(x38711, x38710, x38709);
  nand n38712(x38712, x25790, x84937);
  nand n38713(x38713, x71997, x38708);
  nand n38714(x38714, x25790, x38711);
  nand n38715(x38715, x38714, x38713);
  nand n38716(x38716, x72002, x84938);
  nand n38717(x38717, x25796, x38715);
  nand n38718(x38718, x38717, x38716);
  nand n38719(x38719, x16745, x36889);
  nand n38720(x38720, x68738, x38722);
  nand n38721(x38721, x38720, x38719);
  nand n38723(x38723, x16745, x36948);
  nand n38724(x38724, x68738, x38726);
  nand n38725(x38725, x38724, x38723);
  nand n38727(x38727, x16745, x37007);
  nand n38728(x38728, x68738, x38730);
  nand n38729(x38729, x38728, x38727);
  nand n38731(x38731, x16745, x37066);
  nand n38732(x38732, x68738, x38734);
  nand n38733(x38733, x38732, x38731);
  nand n38735(x38735, x16745, x37125);
  nand n38736(x38736, x68738, x38738);
  nand n38737(x38737, x38736, x38735);
  nand n38739(x38739, x16745, x37184);
  nand n38740(x38740, x68738, x38742);
  nand n38741(x38741, x38740, x38739);
  nand n38743(x38743, x16745, x37243);
  nand n38744(x38744, x68738, x38746);
  nand n38745(x38745, x38744, x38743);
  nand n38747(x38747, x16745, x37302);
  nand n38748(x38748, x68738, x38750);
  nand n38749(x38749, x38748, x38747);
  nand n38751(x38751, x16745, x37361);
  nand n38752(x38752, x68738, x38754);
  nand n38753(x38753, x38752, x38751);
  nand n38755(x38755, x16745, x37420);
  nand n38756(x38756, x68738, x38758);
  nand n38757(x38757, x38756, x38755);
  nand n38759(x38759, x16745, x37479);
  nand n38760(x38760, x68738, x38762);
  nand n38761(x38761, x38760, x38759);
  nand n38763(x38763, x16745, x37538);
  nand n38764(x38764, x68738, x38766);
  nand n38765(x38765, x38764, x38763);
  nand n38767(x38767, x16745, x37597);
  nand n38768(x38768, x68738, x38770);
  nand n38769(x38769, x38768, x38767);
  nand n38771(x38771, x16745, x37656);
  nand n38772(x38772, x68738, x38774);
  nand n38773(x38773, x38772, x38771);
  nand n38775(x38775, x16745, x37715);
  nand n38776(x38776, x68738, x38778);
  nand n38777(x38777, x38776, x38775);
  nand n38779(x38779, x16745, x37774);
  nand n38780(x38780, x68738, x38782);
  nand n38781(x38781, x38780, x38779);
  nand n38783(x38783, x16745, x37833);
  nand n38784(x38784, x68738, x38786);
  nand n38785(x38785, x38784, x38783);
  nand n38787(x38787, x16745, x37892);
  nand n38788(x38788, x68738, x38790);
  nand n38789(x38789, x38788, x38787);
  nand n38791(x38791, x16745, x37951);
  nand n38792(x38792, x68738, x38794);
  nand n38793(x38793, x38792, x38791);
  nand n38795(x38795, x16745, x38010);
  nand n38796(x38796, x68738, x38798);
  nand n38797(x38797, x38796, x38795);
  nand n38799(x38799, x16745, x38069);
  nand n38800(x38800, x68738, x38802);
  nand n38801(x38801, x38800, x38799);
  nand n38803(x38803, x16745, x38128);
  nand n38804(x38804, x68738, x38806);
  nand n38805(x38805, x38804, x38803);
  nand n38807(x38807, x16745, x38187);
  nand n38808(x38808, x68738, x38810);
  nand n38809(x38809, x38808, x38807);
  nand n38811(x38811, x16745, x38246);
  nand n38812(x38812, x68738, x38814);
  nand n38813(x38813, x38812, x38811);
  nand n38815(x38815, x16745, x38305);
  nand n38816(x38816, x68738, x38818);
  nand n38817(x38817, x38816, x38815);
  nand n38819(x38819, x16745, x38364);
  nand n38820(x38820, x68738, x38822);
  nand n38821(x38821, x38820, x38819);
  nand n38823(x38823, x16745, x38423);
  nand n38824(x38824, x68738, x38826);
  nand n38825(x38825, x38824, x38823);
  nand n38827(x38827, x16745, x38482);
  nand n38828(x38828, x68738, x38830);
  nand n38829(x38829, x38828, x38827);
  nand n38831(x38831, x16745, x38541);
  nand n38832(x38832, x68738, x38834);
  nand n38833(x38833, x38832, x38831);
  nand n38835(x38835, x16745, x38600);
  nand n38836(x38836, x68738, x38838);
  nand n38837(x38837, x38836, x38835);
  nand n38839(x38839, x16745, x38659);
  nand n38840(x38840, x68738, x38842);
  nand n38841(x38841, x38840, x38839);
  nand n38843(x38843, x16745, x38718);
  nand n38844(x38844, x68738, x38846);
  nand n38845(x38845, x38844, x38843);
  nand n38847(x38847, x16747, x73187);
  nand n38848(x38848, x38847, x16746);
  nand n38849(x38849, x16747, x73192);
  nand n38850(x38850, x38849, x16750);
  nand n38851(x38851, x16747, x73197);
  nand n38852(x38852, x38851, x16753);
  nand n38853(x38853, x16747, x73202);
  nand n38854(x38854, x38853, x16756);
  nand n38855(x38855, x16747, x73207);
  nand n38856(x38856, x38855, x16759);
  nand n38857(x38857, x16747, x73212);
  nand n38858(x38858, x38857, x16762);
  nand n38859(x38859, x16747, x73217);
  nand n38860(x38860, x38859, x16765);
  nand n38861(x38861, x16747, x73222);
  nand n38862(x38862, x38861, x16768);
  nand n38863(x38863, x16747, x73227);
  nand n38864(x38864, x38863, x16771);
  nand n38865(x38865, x16747, x73232);
  nand n38866(x38866, x38865, x16774);
  nand n38867(x38867, x16747, x73237);
  nand n38868(x38868, x38867, x16777);
  nand n38869(x38869, x16747, x73242);
  nand n38870(x38870, x38869, x16780);
  nand n38871(x38871, x16747, x73247);
  nand n38872(x38872, x38871, x16783);
  nand n38873(x38873, x16747, x73252);
  nand n38874(x38874, x38873, x16786);
  nand n38875(x38875, x16747, x73257);
  nand n38876(x38876, x38875, x16789);
  nand n38877(x38877, x16747, x73262);
  nand n38878(x38878, x38877, x16792);
  nand n38879(x38879, x16747, x73267);
  nand n38880(x38880, x38879, x16795);
  nand n38881(x38881, x16747, x73272);
  nand n38882(x38882, x38881, x16798);
  nand n38883(x38883, x16747, x73277);
  nand n38884(x38884, x38883, x16801);
  nand n38885(x38885, x16747, x73282);
  nand n38886(x38886, x38885, x16804);
  nand n38887(x38887, x16747, x73287);
  nand n38888(x38888, x38887, x16807);
  nand n38889(x38889, x16747, x73292);
  nand n38890(x38890, x38889, x16810);
  nand n38891(x38891, x16747, x73297);
  nand n38892(x38892, x38891, x16813);
  nand n38893(x38893, x16747, x73302);
  nand n38894(x38894, x38893, x16816);
  nand n38895(x38895, x16747, x73307);
  nand n38896(x38896, x38895, x16819);
  nand n38897(x38897, x16747, x73312);
  nand n38898(x38898, x38897, x16822);
  nand n38899(x38899, x16747, x73317);
  nand n38900(x38900, x38899, x16825);
  nand n38901(x38901, x16747, x73322);
  nand n38902(x38902, x38901, x16828);
  nand n38903(x38903, x16747, x73327);
  nand n38904(x38904, x38903, x16831);
  nand n38905(x38905, x16747, x73332);
  nand n38906(x38906, x38905, x16834);
  nand n38907(x38907, x16747, x73337);
  nand n38908(x38908, x38907, x16837);
  nand n38909(x38909, x16747, x73342);
  nand n38910(x38910, x38909, x16840);
  nand n38943(x38943, x71977, x38911);
  nand n38944(x38944, x16876, x38848);
  nand n38945(x38945, x38944, x38943);
  nand n38946(x38946, x71977, x38912);
  nand n38947(x38947, x16876, x38850);
  nand n38948(x38948, x38947, x38946);
  nand n38949(x38949, x71977, x38913);
  nand n38950(x38950, x16876, x38852);
  nand n38951(x38951, x38950, x38949);
  nand n38952(x38952, x71977, x38914);
  nand n38953(x38953, x16876, x38854);
  nand n38954(x38954, x38953, x38952);
  nand n38955(x38955, x71977, x38915);
  nand n38956(x38956, x16876, x38856);
  nand n38957(x38957, x38956, x38955);
  nand n38958(x38958, x71977, x38916);
  nand n38959(x38959, x16876, x38858);
  nand n38960(x38960, x38959, x38958);
  nand n38961(x38961, x71977, x38917);
  nand n38962(x38962, x16876, x38860);
  nand n38963(x38963, x38962, x38961);
  nand n38964(x38964, x71977, x38918);
  nand n38965(x38965, x16876, x38862);
  nand n38966(x38966, x38965, x38964);
  nand n38967(x38967, x71977, x38919);
  nand n38968(x38968, x16876, x38864);
  nand n38969(x38969, x38968, x38967);
  nand n38970(x38970, x71977, x38920);
  nand n38971(x38971, x16876, x38866);
  nand n38972(x38972, x38971, x38970);
  nand n38973(x38973, x71977, x38921);
  nand n38974(x38974, x16876, x38868);
  nand n38975(x38975, x38974, x38973);
  nand n38976(x38976, x71977, x38922);
  nand n38977(x38977, x16876, x38870);
  nand n38978(x38978, x38977, x38976);
  nand n38979(x38979, x71977, x38923);
  nand n38980(x38980, x16876, x38872);
  nand n38981(x38981, x38980, x38979);
  nand n38982(x38982, x71977, x38924);
  nand n38983(x38983, x16876, x38874);
  nand n38984(x38984, x38983, x38982);
  nand n38985(x38985, x71977, x38925);
  nand n38986(x38986, x16876, x38876);
  nand n38987(x38987, x38986, x38985);
  nand n38988(x38988, x71977, x38926);
  nand n38989(x38989, x16876, x38878);
  nand n38990(x38990, x38989, x38988);
  nand n38991(x38991, x71977, x38927);
  nand n38992(x38992, x16876, x38880);
  nand n38993(x38993, x38992, x38991);
  nand n38994(x38994, x71977, x38928);
  nand n38995(x38995, x16876, x38882);
  nand n38996(x38996, x38995, x38994);
  nand n38997(x38997, x71977, x38929);
  nand n38998(x38998, x16876, x38884);
  nand n38999(x38999, x38998, x38997);
  nand n39000(x39000, x71977, x38930);
  nand n39001(x39001, x16876, x38886);
  nand n39002(x39002, x39001, x39000);
  nand n39003(x39003, x71977, x38931);
  nand n39004(x39004, x16876, x38888);
  nand n39005(x39005, x39004, x39003);
  nand n39006(x39006, x71977, x38932);
  nand n39007(x39007, x16876, x38890);
  nand n39008(x39008, x39007, x39006);
  nand n39009(x39009, x71977, x38933);
  nand n39010(x39010, x16876, x38892);
  nand n39011(x39011, x39010, x39009);
  nand n39012(x39012, x71977, x38934);
  nand n39013(x39013, x16876, x38894);
  nand n39014(x39014, x39013, x39012);
  nand n39015(x39015, x71977, x38935);
  nand n39016(x39016, x16876, x38896);
  nand n39017(x39017, x39016, x39015);
  nand n39018(x39018, x71977, x38936);
  nand n39019(x39019, x16876, x38898);
  nand n39020(x39020, x39019, x39018);
  nand n39021(x39021, x71977, x38937);
  nand n39022(x39022, x16876, x38900);
  nand n39023(x39023, x39022, x39021);
  nand n39024(x39024, x71977, x38938);
  nand n39025(x39025, x16876, x38902);
  nand n39026(x39026, x39025, x39024);
  nand n39027(x39027, x71977, x38939);
  nand n39028(x39028, x16876, x38904);
  nand n39029(x39029, x39028, x39027);
  nand n39030(x39030, x71977, x38940);
  nand n39031(x39031, x16876, x38906);
  nand n39032(x39032, x39031, x39030);
  nand n39033(x39033, x71977, x38941);
  nand n39034(x39034, x16876, x38908);
  nand n39035(x39035, x39034, x39033);
  nand n39036(x39036, x71977, x38942);
  nand n39037(x39037, x16876, x38910);
  nand n39038(x39038, x39037, x39036);
  nand n39039(x39039, x73027, x38945);
  nand n39042(x39042, x39041, x39040);
  nand n39043(x39043, x39042, x39039);
  nand n39045(x39045, x73032, x38948);
  nand n39048(x39048, x39047, x39046);
  nand n39049(x39049, x39048, x39045);
  nand n39051(x39051, x73037, x38951);
  nand n39054(x39054, x39053, x39052);
  nand n39055(x39055, x39054, x39051);
  nand n39057(x39057, x73042, x38954);
  nand n39060(x39060, x39059, x39058);
  nand n39061(x39061, x39060, x39057);
  nand n39063(x39063, x73047, x38957);
  nand n39066(x39066, x39065, x39064);
  nand n39067(x39067, x39066, x39063);
  nand n39069(x39069, x73052, x38960);
  nand n39072(x39072, x39071, x39070);
  nand n39073(x39073, x39072, x39069);
  nand n39075(x39075, x73057, x38963);
  nand n39078(x39078, x39077, x39076);
  nand n39079(x39079, x39078, x39075);
  nand n39081(x39081, x73062, x38966);
  nand n39084(x39084, x39083, x39082);
  nand n39085(x39085, x39084, x39081);
  nand n39087(x39087, x73067, x38969);
  nand n39090(x39090, x39089, x39088);
  nand n39091(x39091, x39090, x39087);
  nand n39093(x39093, x73072, x38972);
  nand n39096(x39096, x39095, x39094);
  nand n39097(x39097, x39096, x39093);
  nand n39099(x39099, x73077, x38975);
  nand n39102(x39102, x39101, x39100);
  nand n39103(x39103, x39102, x39099);
  nand n39105(x39105, x73082, x38978);
  nand n39108(x39108, x39107, x39106);
  nand n39109(x39109, x39108, x39105);
  nand n39111(x39111, x73087, x38981);
  nand n39114(x39114, x39113, x39112);
  nand n39115(x39115, x39114, x39111);
  nand n39117(x39117, x73092, x38984);
  nand n39120(x39120, x39119, x39118);
  nand n39121(x39121, x39120, x39117);
  nand n39123(x39123, x73097, x38987);
  nand n39126(x39126, x39125, x39124);
  nand n39127(x39127, x39126, x39123);
  nand n39129(x39129, x73102, x38990);
  nand n39132(x39132, x39131, x39130);
  nand n39133(x39133, x39132, x39129);
  nand n39135(x39135, x73107, x38993);
  nand n39138(x39138, x39137, x39136);
  nand n39139(x39139, x39138, x39135);
  nand n39141(x39141, x73112, x38996);
  nand n39144(x39144, x39143, x39142);
  nand n39145(x39145, x39144, x39141);
  nand n39147(x39147, x73117, x38999);
  nand n39150(x39150, x39149, x39148);
  nand n39151(x39151, x39150, x39147);
  nand n39153(x39153, x73122, x39002);
  nand n39156(x39156, x39155, x39154);
  nand n39157(x39157, x39156, x39153);
  nand n39159(x39159, x73127, x39005);
  nand n39162(x39162, x39161, x39160);
  nand n39163(x39163, x39162, x39159);
  nand n39165(x39165, x73132, x39008);
  nand n39168(x39168, x39167, x39166);
  nand n39169(x39169, x39168, x39165);
  nand n39171(x39171, x73137, x39011);
  nand n39174(x39174, x39173, x39172);
  nand n39175(x39175, x39174, x39171);
  nand n39177(x39177, x73142, x39014);
  nand n39180(x39180, x39179, x39178);
  nand n39181(x39181, x39180, x39177);
  nand n39183(x39183, x73147, x39017);
  nand n39186(x39186, x39185, x39184);
  nand n39187(x39187, x39186, x39183);
  nand n39189(x39189, x73152, x39020);
  nand n39192(x39192, x39191, x39190);
  nand n39193(x39193, x39192, x39189);
  nand n39195(x39195, x73157, x39023);
  nand n39198(x39198, x39197, x39196);
  nand n39199(x39199, x39198, x39195);
  nand n39201(x39201, x73162, x39026);
  nand n39204(x39204, x39203, x39202);
  nand n39205(x39205, x39204, x39201);
  nand n39207(x39207, x73167, x39029);
  nand n39210(x39210, x39209, x39208);
  nand n39211(x39211, x39210, x39207);
  nand n39213(x39213, x73172, x39032);
  nand n39216(x39216, x39215, x39214);
  nand n39217(x39217, x39216, x39213);
  nand n39219(x39219, x73177, x39035);
  nand n39222(x39222, x39221, x39220);
  nand n39223(x39223, x39222, x39219);
  nand n39225(x39225, x73182, x39038);
  nand n39228(x39228, x39227, x39226);
  nand n39229(x39229, x39228, x39225);
  nand n39261(x39261, x39044, x71977);
  nand n39262(x39262, x39261, x39039);
  nand n39263(x39263, x39050, x39231);
  nand n39264(x39264, x39263, x39045);
  nand n39265(x39265, x39050, x39044);
  nand n39267(x39267, x39056, x39232);
  nand n39268(x39268, x39267, x39051);
  nand n39269(x39269, x39056, x39050);
  nand n39271(x39271, x39062, x39233);
  nand n39272(x39272, x39271, x39057);
  nand n39273(x39273, x39062, x39056);
  nand n39275(x39275, x39068, x39234);
  nand n39276(x39276, x39275, x39063);
  nand n39277(x39277, x39068, x39062);
  nand n39279(x39279, x39074, x39235);
  nand n39280(x39280, x39279, x39069);
  nand n39281(x39281, x39074, x39068);
  nand n39283(x39283, x39080, x39236);
  nand n39284(x39284, x39283, x39075);
  nand n39285(x39285, x39080, x39074);
  nand n39287(x39287, x39086, x39237);
  nand n39288(x39288, x39287, x39081);
  nand n39289(x39289, x39086, x39080);
  nand n39291(x39291, x39092, x39238);
  nand n39292(x39292, x39291, x39087);
  nand n39293(x39293, x39092, x39086);
  nand n39295(x39295, x39098, x39239);
  nand n39296(x39296, x39295, x39093);
  nand n39297(x39297, x39098, x39092);
  nand n39299(x39299, x39104, x39240);
  nand n39300(x39300, x39299, x39099);
  nand n39301(x39301, x39104, x39098);
  nand n39303(x39303, x39110, x39241);
  nand n39304(x39304, x39303, x39105);
  nand n39305(x39305, x39110, x39104);
  nand n39307(x39307, x39116, x39242);
  nand n39308(x39308, x39307, x39111);
  nand n39309(x39309, x39116, x39110);
  nand n39311(x39311, x39122, x39243);
  nand n39312(x39312, x39311, x39117);
  nand n39313(x39313, x39122, x39116);
  nand n39315(x39315, x39128, x39244);
  nand n39316(x39316, x39315, x39123);
  nand n39317(x39317, x39128, x39122);
  nand n39319(x39319, x39134, x39245);
  nand n39320(x39320, x39319, x39129);
  nand n39321(x39321, x39134, x39128);
  nand n39323(x39323, x39140, x39246);
  nand n39324(x39324, x39323, x39135);
  nand n39325(x39325, x39140, x39134);
  nand n39327(x39327, x39146, x39247);
  nand n39328(x39328, x39327, x39141);
  nand n39329(x39329, x39146, x39140);
  nand n39331(x39331, x39152, x39248);
  nand n39332(x39332, x39331, x39147);
  nand n39333(x39333, x39152, x39146);
  nand n39335(x39335, x39158, x39249);
  nand n39336(x39336, x39335, x39153);
  nand n39337(x39337, x39158, x39152);
  nand n39339(x39339, x39164, x39250);
  nand n39340(x39340, x39339, x39159);
  nand n39341(x39341, x39164, x39158);
  nand n39343(x39343, x39170, x39251);
  nand n39344(x39344, x39343, x39165);
  nand n39345(x39345, x39170, x39164);
  nand n39347(x39347, x39176, x39252);
  nand n39348(x39348, x39347, x39171);
  nand n39349(x39349, x39176, x39170);
  nand n39351(x39351, x39182, x39253);
  nand n39352(x39352, x39351, x39177);
  nand n39353(x39353, x39182, x39176);
  nand n39355(x39355, x39188, x39254);
  nand n39356(x39356, x39355, x39183);
  nand n39357(x39357, x39188, x39182);
  nand n39359(x39359, x39194, x39255);
  nand n39360(x39360, x39359, x39189);
  nand n39361(x39361, x39194, x39188);
  nand n39363(x39363, x39200, x39256);
  nand n39364(x39364, x39363, x39195);
  nand n39365(x39365, x39200, x39194);
  nand n39367(x39367, x39206, x39257);
  nand n39368(x39368, x39367, x39201);
  nand n39369(x39369, x39206, x39200);
  nand n39371(x39371, x39212, x39258);
  nand n39372(x39372, x39371, x39207);
  nand n39373(x39373, x39212, x39206);
  nand n39375(x39375, x39218, x39259);
  nand n39376(x39376, x39375, x39213);
  nand n39377(x39377, x39218, x39212);
  nand n39379(x39379, x39224, x39260);
  nand n39380(x39380, x39379, x39219);
  nand n39381(x39381, x39224, x39218);
  nand n39383(x39383, x39266, x71977);
  nand n39385(x39385, x39383, x39384);
  nand n39386(x39386, x39270, x39262);
  nand n39388(x39388, x39386, x39387);
  nand n39389(x39389, x39274, x39264);
  nand n39391(x39391, x39389, x39390);
  nand n39392(x39392, x39274, x39266);
  nand n39394(x39394, x39278, x39268);
  nand n39396(x39396, x39394, x39395);
  nand n39397(x39397, x39278, x39270);
  nand n39399(x39399, x39282, x39272);
  nand n39401(x39401, x39399, x39400);
  nand n39402(x39402, x39282, x39274);
  nand n39404(x39404, x39286, x39276);
  nand n39406(x39406, x39404, x39405);
  nand n39407(x39407, x39286, x39278);
  nand n39409(x39409, x39290, x39280);
  nand n39411(x39411, x39409, x39410);
  nand n39412(x39412, x39290, x39282);
  nand n39414(x39414, x39294, x39284);
  nand n39416(x39416, x39414, x39415);
  nand n39417(x39417, x39294, x39286);
  nand n39419(x39419, x39298, x39288);
  nand n39421(x39421, x39419, x39420);
  nand n39422(x39422, x39298, x39290);
  nand n39424(x39424, x39302, x39292);
  nand n39426(x39426, x39424, x39425);
  nand n39427(x39427, x39302, x39294);
  nand n39429(x39429, x39306, x39296);
  nand n39431(x39431, x39429, x39430);
  nand n39432(x39432, x39306, x39298);
  nand n39434(x39434, x39310, x39300);
  nand n39436(x39436, x39434, x39435);
  nand n39437(x39437, x39310, x39302);
  nand n39439(x39439, x39314, x39304);
  nand n39441(x39441, x39439, x39440);
  nand n39442(x39442, x39314, x39306);
  nand n39444(x39444, x39318, x39308);
  nand n39446(x39446, x39444, x39445);
  nand n39447(x39447, x39318, x39310);
  nand n39449(x39449, x39322, x39312);
  nand n39451(x39451, x39449, x39450);
  nand n39452(x39452, x39322, x39314);
  nand n39454(x39454, x39326, x39316);
  nand n39456(x39456, x39454, x39455);
  nand n39457(x39457, x39326, x39318);
  nand n39459(x39459, x39330, x39320);
  nand n39461(x39461, x39459, x39460);
  nand n39462(x39462, x39330, x39322);
  nand n39464(x39464, x39334, x39324);
  nand n39466(x39466, x39464, x39465);
  nand n39467(x39467, x39334, x39326);
  nand n39469(x39469, x39338, x39328);
  nand n39471(x39471, x39469, x39470);
  nand n39472(x39472, x39338, x39330);
  nand n39474(x39474, x39342, x39332);
  nand n39476(x39476, x39474, x39475);
  nand n39477(x39477, x39342, x39334);
  nand n39479(x39479, x39346, x39336);
  nand n39481(x39481, x39479, x39480);
  nand n39482(x39482, x39346, x39338);
  nand n39484(x39484, x39350, x39340);
  nand n39486(x39486, x39484, x39485);
  nand n39487(x39487, x39350, x39342);
  nand n39489(x39489, x39354, x39344);
  nand n39491(x39491, x39489, x39490);
  nand n39492(x39492, x39354, x39346);
  nand n39494(x39494, x39358, x39348);
  nand n39496(x39496, x39494, x39495);
  nand n39497(x39497, x39358, x39350);
  nand n39499(x39499, x39362, x39352);
  nand n39501(x39501, x39499, x39500);
  nand n39502(x39502, x39362, x39354);
  nand n39504(x39504, x39366, x39356);
  nand n39506(x39506, x39504, x39505);
  nand n39507(x39507, x39366, x39358);
  nand n39509(x39509, x39370, x39360);
  nand n39511(x39511, x39509, x39510);
  nand n39512(x39512, x39370, x39362);
  nand n39514(x39514, x39374, x39364);
  nand n39516(x39516, x39514, x39515);
  nand n39517(x39517, x39374, x39366);
  nand n39519(x39519, x39378, x39368);
  nand n39521(x39521, x39519, x39520);
  nand n39522(x39522, x39378, x39370);
  nand n39524(x39524, x39382, x39372);
  nand n39526(x39526, x39524, x39525);
  nand n39527(x39527, x39382, x39374);
  nand n39529(x39529, x39393, x71977);
  nand n39531(x39531, x39529, x39530);
  nand n39532(x39532, x39398, x39262);
  nand n39534(x39534, x39532, x39533);
  nand n39535(x39535, x39403, x39385);
  nand n39537(x39537, x39535, x39536);
  nand n39538(x39538, x39408, x39388);
  nand n39540(x39540, x39538, x39539);
  nand n39541(x39541, x39413, x39391);
  nand n39543(x39543, x39541, x39542);
  nand n39544(x39544, x39413, x39393);
  nand n39546(x39546, x39418, x39396);
  nand n39548(x39548, x39546, x39547);
  nand n39549(x39549, x39418, x39398);
  nand n39551(x39551, x39423, x39401);
  nand n39553(x39553, x39551, x39552);
  nand n39554(x39554, x39423, x39403);
  nand n39556(x39556, x39428, x39406);
  nand n39558(x39558, x39556, x39557);
  nand n39559(x39559, x39428, x39408);
  nand n39561(x39561, x39433, x39411);
  nand n39563(x39563, x39561, x39562);
  nand n39564(x39564, x39433, x39413);
  nand n39566(x39566, x39438, x39416);
  nand n39568(x39568, x39566, x39567);
  nand n39569(x39569, x39438, x39418);
  nand n39571(x39571, x39443, x39421);
  nand n39573(x39573, x39571, x39572);
  nand n39574(x39574, x39443, x39423);
  nand n39576(x39576, x39448, x39426);
  nand n39578(x39578, x39576, x39577);
  nand n39579(x39579, x39448, x39428);
  nand n39581(x39581, x39453, x39431);
  nand n39583(x39583, x39581, x39582);
  nand n39584(x39584, x39453, x39433);
  nand n39586(x39586, x39458, x39436);
  nand n39588(x39588, x39586, x39587);
  nand n39589(x39589, x39458, x39438);
  nand n39591(x39591, x39463, x39441);
  nand n39593(x39593, x39591, x39592);
  nand n39594(x39594, x39463, x39443);
  nand n39596(x39596, x39468, x39446);
  nand n39598(x39598, x39596, x39597);
  nand n39599(x39599, x39468, x39448);
  nand n39601(x39601, x39473, x39451);
  nand n39603(x39603, x39601, x39602);
  nand n39604(x39604, x39473, x39453);
  nand n39606(x39606, x39478, x39456);
  nand n39608(x39608, x39606, x39607);
  nand n39609(x39609, x39478, x39458);
  nand n39611(x39611, x39483, x39461);
  nand n39613(x39613, x39611, x39612);
  nand n39614(x39614, x39483, x39463);
  nand n39616(x39616, x39488, x39466);
  nand n39618(x39618, x39616, x39617);
  nand n39619(x39619, x39488, x39468);
  nand n39621(x39621, x39493, x39471);
  nand n39623(x39623, x39621, x39622);
  nand n39624(x39624, x39493, x39473);
  nand n39626(x39626, x39498, x39476);
  nand n39628(x39628, x39626, x39627);
  nand n39629(x39629, x39498, x39478);
  nand n39631(x39631, x39503, x39481);
  nand n39633(x39633, x39631, x39632);
  nand n39634(x39634, x39503, x39483);
  nand n39636(x39636, x39508, x39486);
  nand n39638(x39638, x39636, x39637);
  nand n39639(x39639, x39508, x39488);
  nand n39641(x39641, x39513, x39491);
  nand n39643(x39643, x39641, x39642);
  nand n39644(x39644, x39513, x39493);
  nand n39646(x39646, x39518, x39496);
  nand n39648(x39648, x39646, x39647);
  nand n39649(x39649, x39518, x39498);
  nand n39651(x39651, x39523, x39501);
  nand n39653(x39653, x39651, x39652);
  nand n39654(x39654, x39523, x39503);
  nand n39656(x39656, x39528, x39506);
  nand n39658(x39658, x39656, x39657);
  nand n39659(x39659, x39528, x39508);
  nand n39661(x39661, x39545, x71977);
  nand n39663(x39663, x39661, x39662);
  nand n39664(x39664, x39550, x39262);
  nand n39666(x39666, x39664, x39665);
  nand n39667(x39667, x39555, x39385);
  nand n39669(x39669, x39667, x39668);
  nand n39670(x39670, x39560, x39388);
  nand n39672(x39672, x39670, x39671);
  nand n39673(x39673, x39565, x39531);
  nand n39675(x39675, x39673, x39674);
  nand n39676(x39676, x39570, x39534);
  nand n39678(x39678, x39676, x39677);
  nand n39679(x39679, x39575, x39537);
  nand n39681(x39681, x39679, x39680);
  nand n39682(x39682, x39580, x39540);
  nand n39684(x39684, x39682, x39683);
  nand n39685(x39685, x39585, x39543);
  nand n39687(x39687, x39685, x39686);
  nand n39688(x39688, x39585, x39545);
  nand n39690(x39690, x39590, x39548);
  nand n39692(x39692, x39690, x39691);
  nand n39693(x39693, x39590, x39550);
  nand n39695(x39695, x39595, x39553);
  nand n39697(x39697, x39695, x39696);
  nand n39698(x39698, x39595, x39555);
  nand n39700(x39700, x39600, x39558);
  nand n39702(x39702, x39700, x39701);
  nand n39703(x39703, x39600, x39560);
  nand n39705(x39705, x39605, x39563);
  nand n39707(x39707, x39705, x39706);
  nand n39708(x39708, x39605, x39565);
  nand n39710(x39710, x39610, x39568);
  nand n39712(x39712, x39710, x39711);
  nand n39713(x39713, x39610, x39570);
  nand n39715(x39715, x39615, x39573);
  nand n39717(x39717, x39715, x39716);
  nand n39718(x39718, x39615, x39575);
  nand n39720(x39720, x39620, x39578);
  nand n39722(x39722, x39720, x39721);
  nand n39723(x39723, x39620, x39580);
  nand n39725(x39725, x39625, x39583);
  nand n39727(x39727, x39725, x39726);
  nand n39728(x39728, x39625, x39585);
  nand n39730(x39730, x39630, x39588);
  nand n39732(x39732, x39730, x39731);
  nand n39733(x39733, x39630, x39590);
  nand n39735(x39735, x39635, x39593);
  nand n39737(x39737, x39735, x39736);
  nand n39738(x39738, x39635, x39595);
  nand n39740(x39740, x39640, x39598);
  nand n39742(x39742, x39740, x39741);
  nand n39743(x39743, x39640, x39600);
  nand n39745(x39745, x39645, x39603);
  nand n39747(x39747, x39745, x39746);
  nand n39748(x39748, x39645, x39605);
  nand n39750(x39750, x39650, x39608);
  nand n39752(x39752, x39750, x39751);
  nand n39753(x39753, x39650, x39610);
  nand n39755(x39755, x39655, x39613);
  nand n39757(x39757, x39755, x39756);
  nand n39758(x39758, x39655, x39615);
  nand n39760(x39760, x39660, x39618);
  nand n39762(x39762, x39760, x39761);
  nand n39763(x39763, x39660, x39620);
  nand n39765(x39765, x39689, x71977);
  nand n39767(x39767, x39765, x39766);
  nand n39768(x39768, x39694, x39262);
  nand n39770(x39770, x39768, x39769);
  nand n39771(x39771, x39699, x39385);
  nand n39773(x39773, x39771, x39772);
  nand n39774(x39774, x39704, x39388);
  nand n39776(x39776, x39774, x39775);
  nand n39777(x39777, x39709, x39531);
  nand n39779(x39779, x39777, x39778);
  nand n39780(x39780, x39714, x39534);
  nand n39782(x39782, x39780, x39781);
  nand n39783(x39783, x39719, x39537);
  nand n39785(x39785, x39783, x39784);
  nand n39786(x39786, x39724, x39540);
  nand n39788(x39788, x39786, x39787);
  nand n39789(x39789, x39729, x39663);
  nand n39791(x39791, x39789, x39790);
  nand n39792(x39792, x39734, x39666);
  nand n39794(x39794, x39792, x39793);
  nand n39795(x39795, x39739, x39669);
  nand n39797(x39797, x39795, x39796);
  nand n39798(x39798, x39744, x39672);
  nand n39800(x39800, x39798, x39799);
  nand n39801(x39801, x39749, x39675);
  nand n39803(x39803, x39801, x39802);
  nand n39804(x39804, x39754, x39678);
  nand n39806(x39806, x39804, x39805);
  nand n39807(x39807, x39759, x39681);
  nand n39809(x39809, x39807, x39808);
  nand n39810(x39810, x39764, x39684);
  nand n39812(x39812, x39810, x39811);
  nand n39813(x39813, x39043, x16876);
  nand n39814(x39814, x39813, x39261);
  nand n39816(x39816, x39050, x39262);
  nand n39818(x39818, x39049, x39817);
  nand n39819(x39819, x39818, x39816);
  nand n39821(x39821, x39056, x39385);
  nand n39823(x39823, x39055, x39822);
  nand n39824(x39824, x39823, x39821);
  nand n39826(x39826, x39062, x39388);
  nand n39828(x39828, x39061, x39827);
  nand n39829(x39829, x39828, x39826);
  nand n39831(x39831, x39068, x39531);
  nand n39833(x39833, x39067, x39832);
  nand n39834(x39834, x39833, x39831);
  nand n39836(x39836, x39074, x39534);
  nand n39838(x39838, x39073, x39837);
  nand n39839(x39839, x39838, x39836);
  nand n39841(x39841, x39080, x39537);
  nand n39843(x39843, x39079, x39842);
  nand n39844(x39844, x39843, x39841);
  nand n39846(x39846, x39086, x39540);
  nand n39848(x39848, x39085, x39847);
  nand n39849(x39849, x39848, x39846);
  nand n39851(x39851, x39092, x39663);
  nand n39853(x39853, x39091, x39852);
  nand n39854(x39854, x39853, x39851);
  nand n39856(x39856, x39098, x39666);
  nand n39858(x39858, x39097, x39857);
  nand n39859(x39859, x39858, x39856);
  nand n39861(x39861, x39104, x39669);
  nand n39863(x39863, x39103, x39862);
  nand n39864(x39864, x39863, x39861);
  nand n39866(x39866, x39110, x39672);
  nand n39868(x39868, x39109, x39867);
  nand n39869(x39869, x39868, x39866);
  nand n39871(x39871, x39116, x39675);
  nand n39873(x39873, x39115, x39872);
  nand n39874(x39874, x39873, x39871);
  nand n39876(x39876, x39122, x39678);
  nand n39878(x39878, x39121, x39877);
  nand n39879(x39879, x39878, x39876);
  nand n39881(x39881, x39128, x39681);
  nand n39883(x39883, x39127, x39882);
  nand n39884(x39884, x39883, x39881);
  nand n39886(x39886, x39134, x39684);
  nand n39888(x39888, x39133, x39887);
  nand n39889(x39889, x39888, x39886);
  nand n39891(x39891, x39140, x39767);
  nand n39893(x39893, x39139, x39892);
  nand n39894(x39894, x39893, x39891);
  nand n39896(x39896, x39146, x39770);
  nand n39898(x39898, x39145, x39897);
  nand n39899(x39899, x39898, x39896);
  nand n39901(x39901, x39152, x39773);
  nand n39903(x39903, x39151, x39902);
  nand n39904(x39904, x39903, x39901);
  nand n39906(x39906, x39158, x39776);
  nand n39908(x39908, x39157, x39907);
  nand n39909(x39909, x39908, x39906);
  nand n39911(x39911, x39164, x39779);
  nand n39913(x39913, x39163, x39912);
  nand n39914(x39914, x39913, x39911);
  nand n39916(x39916, x39170, x39782);
  nand n39918(x39918, x39169, x39917);
  nand n39919(x39919, x39918, x39916);
  nand n39921(x39921, x39176, x39785);
  nand n39923(x39923, x39175, x39922);
  nand n39924(x39924, x39923, x39921);
  nand n39926(x39926, x39182, x39788);
  nand n39928(x39928, x39181, x39927);
  nand n39929(x39929, x39928, x39926);
  nand n39931(x39931, x39188, x39791);
  nand n39933(x39933, x39187, x39932);
  nand n39934(x39934, x39933, x39931);
  nand n39936(x39936, x39194, x39794);
  nand n39938(x39938, x39193, x39937);
  nand n39939(x39939, x39938, x39936);
  nand n39941(x39941, x39200, x39797);
  nand n39943(x39943, x39199, x39942);
  nand n39944(x39944, x39943, x39941);
  nand n39946(x39946, x39206, x39800);
  nand n39948(x39948, x39205, x39947);
  nand n39949(x39949, x39948, x39946);
  nand n39951(x39951, x39212, x39803);
  nand n39953(x39953, x39211, x39952);
  nand n39954(x39954, x39953, x39951);
  nand n39956(x39956, x39218, x39806);
  nand n39958(x39958, x39217, x39957);
  nand n39959(x39959, x39958, x39956);
  nand n39961(x39961, x39224, x39809);
  nand n39963(x39963, x39223, x39962);
  nand n39964(x39964, x39963, x39961);
  nand n39966(x39966, x39230, x39812);
  nand n39968(x39968, x39229, x39967);
  nand n39969(x39969, x39968, x39966);
  nand n39971(x39971, x73027, x38848);
  nand n39972(x39972, x73032, x38848);
  nand n39974(x39974, x73027, x38850);
  nand n39976(x39976, x73037, x38848);
  nand n39978(x39978, x73032, x38850);
  nand n39980(x39980, x73027, x38852);
  nand n39982(x39982, x73042, x38848);
  nand n39984(x39984, x73037, x38850);
  nand n39986(x39986, x73032, x38852);
  nand n39988(x39988, x73027, x38854);
  nand n39989(x39989, x73047, x38848);
  nand n39991(x39991, x73042, x38850);
  nand n39993(x39993, x73037, x38852);
  nand n39995(x39995, x73032, x38854);
  nand n39997(x39997, x73027, x38856);
  nand n39999(x39999, x73052, x38848);
  nand n40001(x40001, x73047, x38850);
  nand n40003(x40003, x73042, x38852);
  nand n40005(x40005, x73037, x38854);
  nand n40007(x40007, x73032, x38856);
  nand n40009(x40009, x73027, x38858);
  nand n40011(x40011, x73057, x38848);
  nand n40013(x40013, x73052, x38850);
  nand n40015(x40015, x73047, x38852);
  nand n40017(x40017, x73042, x38854);
  nand n40019(x40019, x73037, x38856);
  nand n40021(x40021, x73032, x38858);
  nand n40023(x40023, x73027, x38860);
  nand n40024(x40024, x73062, x38848);
  nand n40026(x40026, x73057, x38850);
  nand n40028(x40028, x73052, x38852);
  nand n40030(x40030, x73047, x38854);
  nand n40032(x40032, x73042, x38856);
  nand n40034(x40034, x73037, x38858);
  nand n40036(x40036, x73032, x38860);
  nand n40038(x40038, x73027, x38862);
  nand n40040(x40040, x73067, x38848);
  nand n40042(x40042, x73062, x38850);
  nand n40044(x40044, x73057, x38852);
  nand n40046(x40046, x73052, x38854);
  nand n40048(x40048, x73047, x38856);
  nand n40050(x40050, x73042, x38858);
  nand n40052(x40052, x73037, x38860);
  nand n40054(x40054, x73032, x38862);
  nand n40056(x40056, x73027, x38864);
  nand n40058(x40058, x73072, x38848);
  nand n40060(x40060, x73067, x38850);
  nand n40062(x40062, x73062, x38852);
  nand n40064(x40064, x73057, x38854);
  nand n40066(x40066, x73052, x38856);
  nand n40068(x40068, x73047, x38858);
  nand n40070(x40070, x73042, x38860);
  nand n40072(x40072, x73037, x38862);
  nand n40074(x40074, x73032, x38864);
  nand n40076(x40076, x73027, x38866);
  nand n40077(x40077, x73077, x38848);
  nand n40079(x40079, x73072, x38850);
  nand n40081(x40081, x73067, x38852);
  nand n40083(x40083, x73062, x38854);
  nand n40085(x40085, x73057, x38856);
  nand n40087(x40087, x73052, x38858);
  nand n40089(x40089, x73047, x38860);
  nand n40091(x40091, x73042, x38862);
  nand n40093(x40093, x73037, x38864);
  nand n40095(x40095, x73032, x38866);
  nand n40097(x40097, x73027, x38868);
  nand n40099(x40099, x73082, x38848);
  nand n40101(x40101, x73077, x38850);
  nand n40103(x40103, x73072, x38852);
  nand n40105(x40105, x73067, x38854);
  nand n40107(x40107, x73062, x38856);
  nand n40109(x40109, x73057, x38858);
  nand n40111(x40111, x73052, x38860);
  nand n40113(x40113, x73047, x38862);
  nand n40115(x40115, x73042, x38864);
  nand n40117(x40117, x73037, x38866);
  nand n40119(x40119, x73032, x38868);
  nand n40121(x40121, x73027, x38870);
  nand n40123(x40123, x73087, x38848);
  nand n40125(x40125, x73082, x38850);
  nand n40127(x40127, x73077, x38852);
  nand n40129(x40129, x73072, x38854);
  nand n40131(x40131, x73067, x38856);
  nand n40133(x40133, x73062, x38858);
  nand n40135(x40135, x73057, x38860);
  nand n40137(x40137, x73052, x38862);
  nand n40139(x40139, x73047, x38864);
  nand n40141(x40141, x73042, x38866);
  nand n40143(x40143, x73037, x38868);
  nand n40145(x40145, x73032, x38870);
  nand n40147(x40147, x73027, x38872);
  nand n40148(x40148, x73092, x38848);
  nand n40150(x40150, x73087, x38850);
  nand n40152(x40152, x73082, x38852);
  nand n40154(x40154, x73077, x38854);
  nand n40156(x40156, x73072, x38856);
  nand n40158(x40158, x73067, x38858);
  nand n40160(x40160, x73062, x38860);
  nand n40162(x40162, x73057, x38862);
  nand n40164(x40164, x73052, x38864);
  nand n40166(x40166, x73047, x38866);
  nand n40168(x40168, x73042, x38868);
  nand n40170(x40170, x73037, x38870);
  nand n40172(x40172, x73032, x38872);
  nand n40174(x40174, x73027, x38874);
  nand n40176(x40176, x73097, x38848);
  nand n40178(x40178, x73092, x38850);
  nand n40180(x40180, x73087, x38852);
  nand n40182(x40182, x73082, x38854);
  nand n40184(x40184, x73077, x38856);
  nand n40186(x40186, x73072, x38858);
  nand n40188(x40188, x73067, x38860);
  nand n40190(x40190, x73062, x38862);
  nand n40192(x40192, x73057, x38864);
  nand n40194(x40194, x73052, x38866);
  nand n40196(x40196, x73047, x38868);
  nand n40198(x40198, x73042, x38870);
  nand n40200(x40200, x73037, x38872);
  nand n40202(x40202, x73032, x38874);
  nand n40204(x40204, x73027, x38876);
  nand n40206(x40206, x73102, x38848);
  nand n40208(x40208, x73097, x38850);
  nand n40210(x40210, x73092, x38852);
  nand n40212(x40212, x73087, x38854);
  nand n40214(x40214, x73082, x38856);
  nand n40216(x40216, x73077, x38858);
  nand n40218(x40218, x73072, x38860);
  nand n40220(x40220, x73067, x38862);
  nand n40222(x40222, x73062, x38864);
  nand n40224(x40224, x73057, x38866);
  nand n40226(x40226, x73052, x38868);
  nand n40228(x40228, x73047, x38870);
  nand n40230(x40230, x73042, x38872);
  nand n40232(x40232, x73037, x38874);
  nand n40234(x40234, x73032, x38876);
  nand n40236(x40236, x73027, x38878);
  nand n40237(x40237, x73107, x38848);
  nand n40239(x40239, x73102, x38850);
  nand n40241(x40241, x73097, x38852);
  nand n40243(x40243, x73092, x38854);
  nand n40245(x40245, x73087, x38856);
  nand n40247(x40247, x73082, x38858);
  nand n40249(x40249, x73077, x38860);
  nand n40251(x40251, x73072, x38862);
  nand n40253(x40253, x73067, x38864);
  nand n40255(x40255, x73062, x38866);
  nand n40257(x40257, x73057, x38868);
  nand n40259(x40259, x73052, x38870);
  nand n40261(x40261, x73047, x38872);
  nand n40263(x40263, x73042, x38874);
  nand n40265(x40265, x73037, x38876);
  nand n40267(x40267, x73032, x38878);
  nand n40269(x40269, x73027, x38880);
  nand n40271(x40271, x73112, x38848);
  nand n40273(x40273, x73107, x38850);
  nand n40275(x40275, x73102, x38852);
  nand n40277(x40277, x73097, x38854);
  nand n40279(x40279, x73092, x38856);
  nand n40281(x40281, x73087, x38858);
  nand n40283(x40283, x73082, x38860);
  nand n40285(x40285, x73077, x38862);
  nand n40287(x40287, x73072, x38864);
  nand n40289(x40289, x73067, x38866);
  nand n40291(x40291, x73062, x38868);
  nand n40293(x40293, x73057, x38870);
  nand n40295(x40295, x73052, x38872);
  nand n40297(x40297, x73047, x38874);
  nand n40299(x40299, x73042, x38876);
  nand n40301(x40301, x73037, x38878);
  nand n40303(x40303, x73032, x38880);
  nand n40305(x40305, x73027, x38882);
  nand n40307(x40307, x73117, x38848);
  nand n40309(x40309, x73112, x38850);
  nand n40311(x40311, x73107, x38852);
  nand n40313(x40313, x73102, x38854);
  nand n40315(x40315, x73097, x38856);
  nand n40317(x40317, x73092, x38858);
  nand n40319(x40319, x73087, x38860);
  nand n40321(x40321, x73082, x38862);
  nand n40323(x40323, x73077, x38864);
  nand n40325(x40325, x73072, x38866);
  nand n40327(x40327, x73067, x38868);
  nand n40329(x40329, x73062, x38870);
  nand n40331(x40331, x73057, x38872);
  nand n40333(x40333, x73052, x38874);
  nand n40335(x40335, x73047, x38876);
  nand n40337(x40337, x73042, x38878);
  nand n40339(x40339, x73037, x38880);
  nand n40341(x40341, x73032, x38882);
  nand n40343(x40343, x73027, x38884);
  nand n40344(x40344, x73122, x38848);
  nand n40346(x40346, x73117, x38850);
  nand n40348(x40348, x73112, x38852);
  nand n40350(x40350, x73107, x38854);
  nand n40352(x40352, x73102, x38856);
  nand n40354(x40354, x73097, x38858);
  nand n40356(x40356, x73092, x38860);
  nand n40358(x40358, x73087, x38862);
  nand n40360(x40360, x73082, x38864);
  nand n40362(x40362, x73077, x38866);
  nand n40364(x40364, x73072, x38868);
  nand n40366(x40366, x73067, x38870);
  nand n40368(x40368, x73062, x38872);
  nand n40370(x40370, x73057, x38874);
  nand n40372(x40372, x73052, x38876);
  nand n40374(x40374, x73047, x38878);
  nand n40376(x40376, x73042, x38880);
  nand n40378(x40378, x73037, x38882);
  nand n40380(x40380, x73032, x38884);
  nand n40382(x40382, x73027, x38886);
  nand n40384(x40384, x73127, x38848);
  nand n40386(x40386, x73122, x38850);
  nand n40388(x40388, x73117, x38852);
  nand n40390(x40390, x73112, x38854);
  nand n40392(x40392, x73107, x38856);
  nand n40394(x40394, x73102, x38858);
  nand n40396(x40396, x73097, x38860);
  nand n40398(x40398, x73092, x38862);
  nand n40400(x40400, x73087, x38864);
  nand n40402(x40402, x73082, x38866);
  nand n40404(x40404, x73077, x38868);
  nand n40406(x40406, x73072, x38870);
  nand n40408(x40408, x73067, x38872);
  nand n40410(x40410, x73062, x38874);
  nand n40412(x40412, x73057, x38876);
  nand n40414(x40414, x73052, x38878);
  nand n40416(x40416, x73047, x38880);
  nand n40418(x40418, x73042, x38882);
  nand n40420(x40420, x73037, x38884);
  nand n40422(x40422, x73032, x38886);
  nand n40424(x40424, x73027, x38888);
  nand n40426(x40426, x73132, x38848);
  nand n40428(x40428, x73127, x38850);
  nand n40430(x40430, x73122, x38852);
  nand n40432(x40432, x73117, x38854);
  nand n40434(x40434, x73112, x38856);
  nand n40436(x40436, x73107, x38858);
  nand n40438(x40438, x73102, x38860);
  nand n40440(x40440, x73097, x38862);
  nand n40442(x40442, x73092, x38864);
  nand n40444(x40444, x73087, x38866);
  nand n40446(x40446, x73082, x38868);
  nand n40448(x40448, x73077, x38870);
  nand n40450(x40450, x73072, x38872);
  nand n40452(x40452, x73067, x38874);
  nand n40454(x40454, x73062, x38876);
  nand n40456(x40456, x73057, x38878);
  nand n40458(x40458, x73052, x38880);
  nand n40460(x40460, x73047, x38882);
  nand n40462(x40462, x73042, x38884);
  nand n40464(x40464, x73037, x38886);
  nand n40466(x40466, x73032, x38888);
  nand n40468(x40468, x73027, x38890);
  nand n40469(x40469, x73137, x38848);
  nand n40471(x40471, x73132, x38850);
  nand n40473(x40473, x73127, x38852);
  nand n40475(x40475, x73122, x38854);
  nand n40477(x40477, x73117, x38856);
  nand n40479(x40479, x73112, x38858);
  nand n40481(x40481, x73107, x38860);
  nand n40483(x40483, x73102, x38862);
  nand n40485(x40485, x73097, x38864);
  nand n40487(x40487, x73092, x38866);
  nand n40489(x40489, x73087, x38868);
  nand n40491(x40491, x73082, x38870);
  nand n40493(x40493, x73077, x38872);
  nand n40495(x40495, x73072, x38874);
  nand n40497(x40497, x73067, x38876);
  nand n40499(x40499, x73062, x38878);
  nand n40501(x40501, x73057, x38880);
  nand n40503(x40503, x73052, x38882);
  nand n40505(x40505, x73047, x38884);
  nand n40507(x40507, x73042, x38886);
  nand n40509(x40509, x73037, x38888);
  nand n40511(x40511, x73032, x38890);
  nand n40513(x40513, x73027, x38892);
  nand n40515(x40515, x73142, x38848);
  nand n40517(x40517, x73137, x38850);
  nand n40519(x40519, x73132, x38852);
  nand n40521(x40521, x73127, x38854);
  nand n40523(x40523, x73122, x38856);
  nand n40525(x40525, x73117, x38858);
  nand n40527(x40527, x73112, x38860);
  nand n40529(x40529, x73107, x38862);
  nand n40531(x40531, x73102, x38864);
  nand n40533(x40533, x73097, x38866);
  nand n40535(x40535, x73092, x38868);
  nand n40537(x40537, x73087, x38870);
  nand n40539(x40539, x73082, x38872);
  nand n40541(x40541, x73077, x38874);
  nand n40543(x40543, x73072, x38876);
  nand n40545(x40545, x73067, x38878);
  nand n40547(x40547, x73062, x38880);
  nand n40549(x40549, x73057, x38882);
  nand n40551(x40551, x73052, x38884);
  nand n40553(x40553, x73047, x38886);
  nand n40555(x40555, x73042, x38888);
  nand n40557(x40557, x73037, x38890);
  nand n40559(x40559, x73032, x38892);
  nand n40561(x40561, x73027, x38894);
  nand n40563(x40563, x73147, x38848);
  nand n40565(x40565, x73142, x38850);
  nand n40567(x40567, x73137, x38852);
  nand n40569(x40569, x73132, x38854);
  nand n40571(x40571, x73127, x38856);
  nand n40573(x40573, x73122, x38858);
  nand n40575(x40575, x73117, x38860);
  nand n40577(x40577, x73112, x38862);
  nand n40579(x40579, x73107, x38864);
  nand n40581(x40581, x73102, x38866);
  nand n40583(x40583, x73097, x38868);
  nand n40585(x40585, x73092, x38870);
  nand n40587(x40587, x73087, x38872);
  nand n40589(x40589, x73082, x38874);
  nand n40591(x40591, x73077, x38876);
  nand n40593(x40593, x73072, x38878);
  nand n40595(x40595, x73067, x38880);
  nand n40597(x40597, x73062, x38882);
  nand n40599(x40599, x73057, x38884);
  nand n40601(x40601, x73052, x38886);
  nand n40603(x40603, x73047, x38888);
  nand n40605(x40605, x73042, x38890);
  nand n40607(x40607, x73037, x38892);
  nand n40609(x40609, x73032, x38894);
  nand n40611(x40611, x73027, x38896);
  nand n40612(x40612, x73152, x38848);
  nand n40614(x40614, x73147, x38850);
  nand n40616(x40616, x73142, x38852);
  nand n40618(x40618, x73137, x38854);
  nand n40620(x40620, x73132, x38856);
  nand n40622(x40622, x73127, x38858);
  nand n40624(x40624, x73122, x38860);
  nand n40626(x40626, x73117, x38862);
  nand n40628(x40628, x73112, x38864);
  nand n40630(x40630, x73107, x38866);
  nand n40632(x40632, x73102, x38868);
  nand n40634(x40634, x73097, x38870);
  nand n40636(x40636, x73092, x38872);
  nand n40638(x40638, x73087, x38874);
  nand n40640(x40640, x73082, x38876);
  nand n40642(x40642, x73077, x38878);
  nand n40644(x40644, x73072, x38880);
  nand n40646(x40646, x73067, x38882);
  nand n40648(x40648, x73062, x38884);
  nand n40650(x40650, x73057, x38886);
  nand n40652(x40652, x73052, x38888);
  nand n40654(x40654, x73047, x38890);
  nand n40656(x40656, x73042, x38892);
  nand n40658(x40658, x73037, x38894);
  nand n40660(x40660, x73032, x38896);
  nand n40662(x40662, x73027, x38898);
  nand n40664(x40664, x73157, x38848);
  nand n40666(x40666, x73152, x38850);
  nand n40668(x40668, x73147, x38852);
  nand n40670(x40670, x73142, x38854);
  nand n40672(x40672, x73137, x38856);
  nand n40674(x40674, x73132, x38858);
  nand n40676(x40676, x73127, x38860);
  nand n40678(x40678, x73122, x38862);
  nand n40680(x40680, x73117, x38864);
  nand n40682(x40682, x73112, x38866);
  nand n40684(x40684, x73107, x38868);
  nand n40686(x40686, x73102, x38870);
  nand n40688(x40688, x73097, x38872);
  nand n40690(x40690, x73092, x38874);
  nand n40692(x40692, x73087, x38876);
  nand n40694(x40694, x73082, x38878);
  nand n40696(x40696, x73077, x38880);
  nand n40698(x40698, x73072, x38882);
  nand n40700(x40700, x73067, x38884);
  nand n40702(x40702, x73062, x38886);
  nand n40704(x40704, x73057, x38888);
  nand n40706(x40706, x73052, x38890);
  nand n40708(x40708, x73047, x38892);
  nand n40710(x40710, x73042, x38894);
  nand n40712(x40712, x73037, x38896);
  nand n40714(x40714, x73032, x38898);
  nand n40716(x40716, x73027, x38900);
  nand n40718(x40718, x73162, x38848);
  nand n40720(x40720, x73157, x38850);
  nand n40722(x40722, x73152, x38852);
  nand n40724(x40724, x73147, x38854);
  nand n40726(x40726, x73142, x38856);
  nand n40728(x40728, x73137, x38858);
  nand n40730(x40730, x73132, x38860);
  nand n40732(x40732, x73127, x38862);
  nand n40734(x40734, x73122, x38864);
  nand n40736(x40736, x73117, x38866);
  nand n40738(x40738, x73112, x38868);
  nand n40740(x40740, x73107, x38870);
  nand n40742(x40742, x73102, x38872);
  nand n40744(x40744, x73097, x38874);
  nand n40746(x40746, x73092, x38876);
  nand n40748(x40748, x73087, x38878);
  nand n40750(x40750, x73082, x38880);
  nand n40752(x40752, x73077, x38882);
  nand n40754(x40754, x73072, x38884);
  nand n40756(x40756, x73067, x38886);
  nand n40758(x40758, x73062, x38888);
  nand n40760(x40760, x73057, x38890);
  nand n40762(x40762, x73052, x38892);
  nand n40764(x40764, x73047, x38894);
  nand n40766(x40766, x73042, x38896);
  nand n40768(x40768, x73037, x38898);
  nand n40770(x40770, x73032, x38900);
  nand n40772(x40772, x73027, x38902);
  nand n40773(x40773, x73167, x38848);
  nand n40775(x40775, x73162, x38850);
  nand n40777(x40777, x73157, x38852);
  nand n40779(x40779, x73152, x38854);
  nand n40781(x40781, x73147, x38856);
  nand n40783(x40783, x73142, x38858);
  nand n40785(x40785, x73137, x38860);
  nand n40787(x40787, x73132, x38862);
  nand n40789(x40789, x73127, x38864);
  nand n40791(x40791, x73122, x38866);
  nand n40793(x40793, x73117, x38868);
  nand n40795(x40795, x73112, x38870);
  nand n40797(x40797, x73107, x38872);
  nand n40799(x40799, x73102, x38874);
  nand n40801(x40801, x73097, x38876);
  nand n40803(x40803, x73092, x38878);
  nand n40805(x40805, x73087, x38880);
  nand n40807(x40807, x73082, x38882);
  nand n40809(x40809, x73077, x38884);
  nand n40811(x40811, x73072, x38886);
  nand n40813(x40813, x73067, x38888);
  nand n40815(x40815, x73062, x38890);
  nand n40817(x40817, x73057, x38892);
  nand n40819(x40819, x73052, x38894);
  nand n40821(x40821, x73047, x38896);
  nand n40823(x40823, x73042, x38898);
  nand n40825(x40825, x73037, x38900);
  nand n40827(x40827, x73032, x38902);
  nand n40829(x40829, x73027, x38904);
  nand n40831(x40831, x73172, x38848);
  nand n40833(x40833, x73167, x38850);
  nand n40835(x40835, x73162, x38852);
  nand n40837(x40837, x73157, x38854);
  nand n40839(x40839, x73152, x38856);
  nand n40841(x40841, x73147, x38858);
  nand n40843(x40843, x73142, x38860);
  nand n40845(x40845, x73137, x38862);
  nand n40847(x40847, x73132, x38864);
  nand n40849(x40849, x73127, x38866);
  nand n40851(x40851, x73122, x38868);
  nand n40853(x40853, x73117, x38870);
  nand n40855(x40855, x73112, x38872);
  nand n40857(x40857, x73107, x38874);
  nand n40859(x40859, x73102, x38876);
  nand n40861(x40861, x73097, x38878);
  nand n40863(x40863, x73092, x38880);
  nand n40865(x40865, x73087, x38882);
  nand n40867(x40867, x73082, x38884);
  nand n40869(x40869, x73077, x38886);
  nand n40871(x40871, x73072, x38888);
  nand n40873(x40873, x73067, x38890);
  nand n40875(x40875, x73062, x38892);
  nand n40877(x40877, x73057, x38894);
  nand n40879(x40879, x73052, x38896);
  nand n40881(x40881, x73047, x38898);
  nand n40883(x40883, x73042, x38900);
  nand n40885(x40885, x73037, x38902);
  nand n40887(x40887, x73032, x38904);
  nand n40889(x40889, x73027, x38906);
  nand n40891(x40891, x73177, x38848);
  nand n40893(x40893, x73172, x38850);
  nand n40895(x40895, x73167, x38852);
  nand n40897(x40897, x73162, x38854);
  nand n40899(x40899, x73157, x38856);
  nand n40901(x40901, x73152, x38858);
  nand n40903(x40903, x73147, x38860);
  nand n40905(x40905, x73142, x38862);
  nand n40907(x40907, x73137, x38864);
  nand n40909(x40909, x73132, x38866);
  nand n40911(x40911, x73127, x38868);
  nand n40913(x40913, x73122, x38870);
  nand n40915(x40915, x73117, x38872);
  nand n40917(x40917, x73112, x38874);
  nand n40919(x40919, x73107, x38876);
  nand n40921(x40921, x73102, x38878);
  nand n40923(x40923, x73097, x38880);
  nand n40925(x40925, x73092, x38882);
  nand n40927(x40927, x73087, x38884);
  nand n40929(x40929, x73082, x38886);
  nand n40931(x40931, x73077, x38888);
  nand n40933(x40933, x73072, x38890);
  nand n40935(x40935, x73067, x38892);
  nand n40937(x40937, x73062, x38894);
  nand n40939(x40939, x73057, x38896);
  nand n40941(x40941, x73052, x38898);
  nand n40943(x40943, x73047, x38900);
  nand n40945(x40945, x73042, x38902);
  nand n40947(x40947, x73037, x38904);
  nand n40949(x40949, x73032, x38906);
  nand n40951(x40951, x73027, x38908);
  nand n40952(x40952, x73182, x38848);
  nand n40954(x40954, x73177, x38850);
  nand n40956(x40956, x73172, x38852);
  nand n40958(x40958, x73167, x38854);
  nand n40960(x40960, x73162, x38856);
  nand n40962(x40962, x73157, x38858);
  nand n40964(x40964, x73152, x38860);
  nand n40966(x40966, x73147, x38862);
  nand n40968(x40968, x73142, x38864);
  nand n40970(x40970, x73137, x38866);
  nand n40972(x40972, x73132, x38868);
  nand n40974(x40974, x73127, x38870);
  nand n40976(x40976, x73122, x38872);
  nand n40978(x40978, x73117, x38874);
  nand n40980(x40980, x73112, x38876);
  nand n40982(x40982, x73107, x38878);
  nand n40984(x40984, x73102, x38880);
  nand n40986(x40986, x73097, x38882);
  nand n40988(x40988, x73092, x38884);
  nand n40990(x40990, x73087, x38886);
  nand n40992(x40992, x73082, x38888);
  nand n40994(x40994, x73077, x38890);
  nand n40996(x40996, x73072, x38892);
  nand n40998(x40998, x73067, x38894);
  nand n41000(x41000, x73062, x38896);
  nand n41002(x41002, x73057, x38898);
  nand n41004(x41004, x73052, x38900);
  nand n41006(x41006, x73047, x38902);
  nand n41008(x41008, x73042, x38904);
  nand n41010(x41010, x73037, x38906);
  nand n41012(x41012, x73032, x38908);
  nand n41014(x41014, x73027, x38910);
  nand n41016(x41016, x39973, x39975);
  nand n41017(x41017, x39972, x39974);
  nand n41018(x41018, x41017, x41016);
  nand n41019(x41019, x39977, x39979);
  nand n41020(x41020, x39976, x39978);
  nand n41021(x41021, x41020, x41019);
  nand n41023(x41023, x39981, x41022);
  nand n41024(x41024, x39980, x41021);
  nand n41025(x41025, x41024, x41023);
  nand n41026(x41026, x41019, x41023);
  nand n41027(x41027, x39983, x39985);
  nand n41028(x41028, x39982, x39984);
  nand n41029(x41029, x41028, x41027);
  nand n41031(x41031, x39987, x41030);
  nand n41032(x41032, x39986, x41029);
  nand n41033(x41033, x41032, x41031);
  nand n41034(x41034, x41027, x41031);
  nand n41035(x41035, x39990, x39992);
  nand n41036(x41036, x39989, x39991);
  nand n41037(x41037, x41036, x41035);
  nand n41039(x41039, x39994, x41038);
  nand n41040(x41040, x39993, x41037);
  nand n41041(x41041, x41040, x41039);
  nand n41042(x41042, x41035, x41039);
  nand n41043(x41043, x39996, x39998);
  nand n41044(x41044, x39995, x39997);
  nand n41045(x41045, x41044, x41043);
  nand n41046(x41046, x40000, x40002);
  nand n41047(x41047, x39999, x40001);
  nand n41048(x41048, x41047, x41046);
  nand n41050(x41050, x40004, x41049);
  nand n41051(x41051, x40003, x41048);
  nand n41052(x41052, x41051, x41050);
  nand n41053(x41053, x41046, x41050);
  nand n41054(x41054, x40006, x40008);
  nand n41055(x41055, x40005, x40007);
  nand n41056(x41056, x41055, x41054);
  nand n41058(x41058, x40010, x41057);
  nand n41059(x41059, x40009, x41056);
  nand n41060(x41060, x41059, x41058);
  nand n41061(x41061, x41054, x41058);
  nand n41062(x41062, x40012, x40014);
  nand n41063(x41063, x40011, x40013);
  nand n41064(x41064, x41063, x41062);
  nand n41066(x41066, x40016, x41065);
  nand n41067(x41067, x40015, x41064);
  nand n41068(x41068, x41067, x41066);
  nand n41069(x41069, x41062, x41066);
  nand n41070(x41070, x40018, x40020);
  nand n41071(x41071, x40017, x40019);
  nand n41072(x41072, x41071, x41070);
  nand n41074(x41074, x40022, x41073);
  nand n41075(x41075, x40021, x41072);
  nand n41076(x41076, x41075, x41074);
  nand n41078(x41078, x41070, x41074);
  nand n41079(x41079, x40025, x40027);
  nand n41080(x41080, x40024, x40026);
  nand n41081(x41081, x41080, x41079);
  nand n41083(x41083, x40029, x41082);
  nand n41084(x41084, x40028, x41081);
  nand n41085(x41085, x41084, x41083);
  nand n41086(x41086, x41079, x41083);
  nand n41087(x41087, x40031, x40033);
  nand n41088(x41088, x40030, x40032);
  nand n41089(x41089, x41088, x41087);
  nand n41091(x41091, x40035, x41090);
  nand n41092(x41092, x40034, x41089);
  nand n41093(x41093, x41092, x41091);
  nand n41095(x41095, x41087, x41091);
  nand n41096(x41096, x40037, x40039);
  nand n41097(x41097, x40036, x40038);
  nand n41098(x41098, x41097, x41096);
  nand n41099(x41099, x40041, x40043);
  nand n41100(x41100, x40040, x40042);
  nand n41101(x41101, x41100, x41099);
  nand n41103(x41103, x40045, x41102);
  nand n41104(x41104, x40044, x41101);
  nand n41105(x41105, x41104, x41103);
  nand n41106(x41106, x41099, x41103);
  nand n41107(x41107, x40047, x40049);
  nand n41108(x41108, x40046, x40048);
  nand n41109(x41109, x41108, x41107);
  nand n41111(x41111, x40051, x41110);
  nand n41112(x41112, x40050, x41109);
  nand n41113(x41113, x41112, x41111);
  nand n41115(x41115, x41107, x41111);
  nand n41116(x41116, x40053, x40055);
  nand n41117(x41117, x40052, x40054);
  nand n41118(x41118, x41117, x41116);
  nand n41120(x41120, x40057, x41119);
  nand n41121(x41121, x40056, x41118);
  nand n41122(x41122, x41121, x41120);
  nand n41124(x41124, x41116, x41120);
  nand n41125(x41125, x40059, x40061);
  nand n41126(x41126, x40058, x40060);
  nand n41127(x41127, x41126, x41125);
  nand n41129(x41129, x40063, x41128);
  nand n41130(x41130, x40062, x41127);
  nand n41131(x41131, x41130, x41129);
  nand n41132(x41132, x41125, x41129);
  nand n41133(x41133, x40065, x40067);
  nand n41134(x41134, x40064, x40066);
  nand n41135(x41135, x41134, x41133);
  nand n41137(x41137, x40069, x41136);
  nand n41138(x41138, x40068, x41135);
  nand n41139(x41139, x41138, x41137);
  nand n41141(x41141, x41133, x41137);
  nand n41142(x41142, x40071, x40073);
  nand n41143(x41143, x40070, x40072);
  nand n41144(x41144, x41143, x41142);
  nand n41146(x41146, x40075, x41145);
  nand n41147(x41147, x40074, x41144);
  nand n41148(x41148, x41147, x41146);
  nand n41150(x41150, x41142, x41146);
  nand n41151(x41151, x40078, x40080);
  nand n41152(x41152, x40077, x40079);
  nand n41153(x41153, x41152, x41151);
  nand n41155(x41155, x40082, x41154);
  nand n41156(x41156, x40081, x41153);
  nand n41157(x41157, x41156, x41155);
  nand n41158(x41158, x41151, x41155);
  nand n41159(x41159, x40084, x40086);
  nand n41160(x41160, x40083, x40085);
  nand n41161(x41161, x41160, x41159);
  nand n41163(x41163, x40088, x41162);
  nand n41164(x41164, x40087, x41161);
  nand n41165(x41165, x41164, x41163);
  nand n41167(x41167, x41159, x41163);
  nand n41168(x41168, x40090, x40092);
  nand n41169(x41169, x40089, x40091);
  nand n41170(x41170, x41169, x41168);
  nand n41172(x41172, x40094, x41171);
  nand n41173(x41173, x40093, x41170);
  nand n41174(x41174, x41173, x41172);
  nand n41176(x41176, x41168, x41172);
  nand n41177(x41177, x40096, x40098);
  nand n41178(x41178, x40095, x40097);
  nand n41179(x41179, x41178, x41177);
  nand n41180(x41180, x40100, x40102);
  nand n41181(x41181, x40099, x40101);
  nand n41182(x41182, x41181, x41180);
  nand n41184(x41184, x40104, x41183);
  nand n41185(x41185, x40103, x41182);
  nand n41186(x41186, x41185, x41184);
  nand n41187(x41187, x41180, x41184);
  nand n41188(x41188, x40106, x40108);
  nand n41189(x41189, x40105, x40107);
  nand n41190(x41190, x41189, x41188);
  nand n41192(x41192, x40110, x41191);
  nand n41193(x41193, x40109, x41190);
  nand n41194(x41194, x41193, x41192);
  nand n41196(x41196, x41188, x41192);
  nand n41197(x41197, x40112, x40114);
  nand n41198(x41198, x40111, x40113);
  nand n41199(x41199, x41198, x41197);
  nand n41201(x41201, x40116, x41200);
  nand n41202(x41202, x40115, x41199);
  nand n41203(x41203, x41202, x41201);
  nand n41205(x41205, x41197, x41201);
  nand n41206(x41206, x40118, x40120);
  nand n41207(x41207, x40117, x40119);
  nand n41208(x41208, x41207, x41206);
  nand n41210(x41210, x40122, x41209);
  nand n41211(x41211, x40121, x41208);
  nand n41212(x41212, x41211, x41210);
  nand n41214(x41214, x41206, x41210);
  nand n41215(x41215, x40124, x40126);
  nand n41216(x41216, x40123, x40125);
  nand n41217(x41217, x41216, x41215);
  nand n41219(x41219, x40128, x41218);
  nand n41220(x41220, x40127, x41217);
  nand n41221(x41221, x41220, x41219);
  nand n41222(x41222, x41215, x41219);
  nand n41223(x41223, x40130, x40132);
  nand n41224(x41224, x40129, x40131);
  nand n41225(x41225, x41224, x41223);
  nand n41227(x41227, x40134, x41226);
  nand n41228(x41228, x40133, x41225);
  nand n41229(x41229, x41228, x41227);
  nand n41231(x41231, x41223, x41227);
  nand n41232(x41232, x40136, x40138);
  nand n41233(x41233, x40135, x40137);
  nand n41234(x41234, x41233, x41232);
  nand n41236(x41236, x40140, x41235);
  nand n41237(x41237, x40139, x41234);
  nand n41238(x41238, x41237, x41236);
  nand n41240(x41240, x41232, x41236);
  nand n41241(x41241, x40142, x40144);
  nand n41242(x41242, x40141, x40143);
  nand n41243(x41243, x41242, x41241);
  nand n41245(x41245, x40146, x41244);
  nand n41246(x41246, x40145, x41243);
  nand n41247(x41247, x41246, x41245);
  nand n41249(x41249, x41241, x41245);
  nand n41250(x41250, x40149, x40151);
  nand n41251(x41251, x40148, x40150);
  nand n41252(x41252, x41251, x41250);
  nand n41254(x41254, x40153, x41253);
  nand n41255(x41255, x40152, x41252);
  nand n41256(x41256, x41255, x41254);
  nand n41257(x41257, x41250, x41254);
  nand n41258(x41258, x40155, x40157);
  nand n41259(x41259, x40154, x40156);
  nand n41260(x41260, x41259, x41258);
  nand n41262(x41262, x40159, x41261);
  nand n41263(x41263, x40158, x41260);
  nand n41264(x41264, x41263, x41262);
  nand n41266(x41266, x41258, x41262);
  nand n41267(x41267, x40161, x40163);
  nand n41268(x41268, x40160, x40162);
  nand n41269(x41269, x41268, x41267);
  nand n41271(x41271, x40165, x41270);
  nand n41272(x41272, x40164, x41269);
  nand n41273(x41273, x41272, x41271);
  nand n41275(x41275, x41267, x41271);
  nand n41276(x41276, x40167, x40169);
  nand n41277(x41277, x40166, x40168);
  nand n41278(x41278, x41277, x41276);
  nand n41280(x41280, x40171, x41279);
  nand n41281(x41281, x40170, x41278);
  nand n41282(x41282, x41281, x41280);
  nand n41284(x41284, x41276, x41280);
  nand n41285(x41285, x40173, x40175);
  nand n41286(x41286, x40172, x40174);
  nand n41287(x41287, x41286, x41285);
  nand n41288(x41288, x40177, x40179);
  nand n41289(x41289, x40176, x40178);
  nand n41290(x41290, x41289, x41288);
  nand n41292(x41292, x40181, x41291);
  nand n41293(x41293, x40180, x41290);
  nand n41294(x41294, x41293, x41292);
  nand n41295(x41295, x41288, x41292);
  nand n41296(x41296, x40183, x40185);
  nand n41297(x41297, x40182, x40184);
  nand n41298(x41298, x41297, x41296);
  nand n41300(x41300, x40187, x41299);
  nand n41301(x41301, x40186, x41298);
  nand n41302(x41302, x41301, x41300);
  nand n41304(x41304, x41296, x41300);
  nand n41305(x41305, x40189, x40191);
  nand n41306(x41306, x40188, x40190);
  nand n41307(x41307, x41306, x41305);
  nand n41309(x41309, x40193, x41308);
  nand n41310(x41310, x40192, x41307);
  nand n41311(x41311, x41310, x41309);
  nand n41313(x41313, x41305, x41309);
  nand n41314(x41314, x40195, x40197);
  nand n41315(x41315, x40194, x40196);
  nand n41316(x41316, x41315, x41314);
  nand n41318(x41318, x40199, x41317);
  nand n41319(x41319, x40198, x41316);
  nand n41320(x41320, x41319, x41318);
  nand n41322(x41322, x41314, x41318);
  nand n41323(x41323, x40201, x40203);
  nand n41324(x41324, x40200, x40202);
  nand n41325(x41325, x41324, x41323);
  nand n41327(x41327, x40205, x41326);
  nand n41328(x41328, x40204, x41325);
  nand n41329(x41329, x41328, x41327);
  nand n41330(x41330, x41323, x41327);
  nand n41331(x41331, x40207, x40209);
  nand n41332(x41332, x40206, x40208);
  nand n41333(x41333, x41332, x41331);
  nand n41335(x41335, x40211, x41334);
  nand n41336(x41336, x40210, x41333);
  nand n41337(x41337, x41336, x41335);
  nand n41338(x41338, x41331, x41335);
  nand n41339(x41339, x40213, x40215);
  nand n41340(x41340, x40212, x40214);
  nand n41341(x41341, x41340, x41339);
  nand n41343(x41343, x40217, x41342);
  nand n41344(x41344, x40216, x41341);
  nand n41345(x41345, x41344, x41343);
  nand n41347(x41347, x41339, x41343);
  nand n41348(x41348, x40219, x40221);
  nand n41349(x41349, x40218, x40220);
  nand n41350(x41350, x41349, x41348);
  nand n41352(x41352, x40223, x41351);
  nand n41353(x41353, x40222, x41350);
  nand n41354(x41354, x41353, x41352);
  nand n41356(x41356, x41348, x41352);
  nand n41357(x41357, x40225, x40227);
  nand n41358(x41358, x40224, x40226);
  nand n41359(x41359, x41358, x41357);
  nand n41361(x41361, x40229, x41360);
  nand n41362(x41362, x40228, x41359);
  nand n41363(x41363, x41362, x41361);
  nand n41365(x41365, x41357, x41361);
  nand n41366(x41366, x40231, x40233);
  nand n41367(x41367, x40230, x40232);
  nand n41368(x41368, x41367, x41366);
  nand n41370(x41370, x40235, x41369);
  nand n41371(x41371, x40234, x41368);
  nand n41372(x41372, x41371, x41370);
  nand n41374(x41374, x41366, x41370);
  nand n41375(x41375, x40238, x40240);
  nand n41376(x41376, x40237, x40239);
  nand n41377(x41377, x41376, x41375);
  nand n41379(x41379, x40242, x41378);
  nand n41380(x41380, x40241, x41377);
  nand n41381(x41381, x41380, x41379);
  nand n41382(x41382, x41375, x41379);
  nand n41383(x41383, x40244, x40246);
  nand n41384(x41384, x40243, x40245);
  nand n41385(x41385, x41384, x41383);
  nand n41387(x41387, x40248, x41386);
  nand n41388(x41388, x40247, x41385);
  nand n41389(x41389, x41388, x41387);
  nand n41391(x41391, x41383, x41387);
  nand n41392(x41392, x40250, x40252);
  nand n41393(x41393, x40249, x40251);
  nand n41394(x41394, x41393, x41392);
  nand n41396(x41396, x40254, x41395);
  nand n41397(x41397, x40253, x41394);
  nand n41398(x41398, x41397, x41396);
  nand n41400(x41400, x41392, x41396);
  nand n41401(x41401, x40256, x40258);
  nand n41402(x41402, x40255, x40257);
  nand n41403(x41403, x41402, x41401);
  nand n41405(x41405, x40260, x41404);
  nand n41406(x41406, x40259, x41403);
  nand n41407(x41407, x41406, x41405);
  nand n41409(x41409, x41401, x41405);
  nand n41410(x41410, x40262, x40264);
  nand n41411(x41411, x40261, x40263);
  nand n41412(x41412, x41411, x41410);
  nand n41414(x41414, x40266, x41413);
  nand n41415(x41415, x40265, x41412);
  nand n41416(x41416, x41415, x41414);
  nand n41418(x41418, x41410, x41414);
  nand n41419(x41419, x40268, x40270);
  nand n41420(x41420, x40267, x40269);
  nand n41421(x41421, x41420, x41419);
  nand n41422(x41422, x40272, x40274);
  nand n41423(x41423, x40271, x40273);
  nand n41424(x41424, x41423, x41422);
  nand n41426(x41426, x40276, x41425);
  nand n41427(x41427, x40275, x41424);
  nand n41428(x41428, x41427, x41426);
  nand n41429(x41429, x41422, x41426);
  nand n41430(x41430, x40278, x40280);
  nand n41431(x41431, x40277, x40279);
  nand n41432(x41432, x41431, x41430);
  nand n41434(x41434, x40282, x41433);
  nand n41435(x41435, x40281, x41432);
  nand n41436(x41436, x41435, x41434);
  nand n41438(x41438, x41430, x41434);
  nand n41439(x41439, x40284, x40286);
  nand n41440(x41440, x40283, x40285);
  nand n41441(x41441, x41440, x41439);
  nand n41443(x41443, x40288, x41442);
  nand n41444(x41444, x40287, x41441);
  nand n41445(x41445, x41444, x41443);
  nand n41447(x41447, x41439, x41443);
  nand n41448(x41448, x40290, x40292);
  nand n41449(x41449, x40289, x40291);
  nand n41450(x41450, x41449, x41448);
  nand n41452(x41452, x40294, x41451);
  nand n41453(x41453, x40293, x41450);
  nand n41454(x41454, x41453, x41452);
  nand n41456(x41456, x41448, x41452);
  nand n41457(x41457, x40296, x40298);
  nand n41458(x41458, x40295, x40297);
  nand n41459(x41459, x41458, x41457);
  nand n41461(x41461, x40300, x41460);
  nand n41462(x41462, x40299, x41459);
  nand n41463(x41463, x41462, x41461);
  nand n41465(x41465, x41457, x41461);
  nand n41466(x41466, x40302, x40304);
  nand n41467(x41467, x40301, x40303);
  nand n41468(x41468, x41467, x41466);
  nand n41470(x41470, x40306, x41469);
  nand n41471(x41471, x40305, x41468);
  nand n41472(x41472, x41471, x41470);
  nand n41474(x41474, x41466, x41470);
  nand n41475(x41475, x40308, x40310);
  nand n41476(x41476, x40307, x40309);
  nand n41477(x41477, x41476, x41475);
  nand n41479(x41479, x40312, x41478);
  nand n41480(x41480, x40311, x41477);
  nand n41481(x41481, x41480, x41479);
  nand n41482(x41482, x41475, x41479);
  nand n41483(x41483, x40314, x40316);
  nand n41484(x41484, x40313, x40315);
  nand n41485(x41485, x41484, x41483);
  nand n41487(x41487, x40318, x41486);
  nand n41488(x41488, x40317, x41485);
  nand n41489(x41489, x41488, x41487);
  nand n41491(x41491, x41483, x41487);
  nand n41492(x41492, x40320, x40322);
  nand n41493(x41493, x40319, x40321);
  nand n41494(x41494, x41493, x41492);
  nand n41496(x41496, x40324, x41495);
  nand n41497(x41497, x40323, x41494);
  nand n41498(x41498, x41497, x41496);
  nand n41500(x41500, x41492, x41496);
  nand n41501(x41501, x40326, x40328);
  nand n41502(x41502, x40325, x40327);
  nand n41503(x41503, x41502, x41501);
  nand n41505(x41505, x40330, x41504);
  nand n41506(x41506, x40329, x41503);
  nand n41507(x41507, x41506, x41505);
  nand n41509(x41509, x41501, x41505);
  nand n41510(x41510, x40332, x40334);
  nand n41511(x41511, x40331, x40333);
  nand n41512(x41512, x41511, x41510);
  nand n41514(x41514, x40336, x41513);
  nand n41515(x41515, x40335, x41512);
  nand n41516(x41516, x41515, x41514);
  nand n41518(x41518, x41510, x41514);
  nand n41519(x41519, x40338, x40340);
  nand n41520(x41520, x40337, x40339);
  nand n41521(x41521, x41520, x41519);
  nand n41523(x41523, x40342, x41522);
  nand n41524(x41524, x40341, x41521);
  nand n41525(x41525, x41524, x41523);
  nand n41527(x41527, x41519, x41523);
  nand n41528(x41528, x40345, x40347);
  nand n41529(x41529, x40344, x40346);
  nand n41530(x41530, x41529, x41528);
  nand n41532(x41532, x40349, x41531);
  nand n41533(x41533, x40348, x41530);
  nand n41534(x41534, x41533, x41532);
  nand n41535(x41535, x41528, x41532);
  nand n41536(x41536, x40351, x40353);
  nand n41537(x41537, x40350, x40352);
  nand n41538(x41538, x41537, x41536);
  nand n41540(x41540, x40355, x41539);
  nand n41541(x41541, x40354, x41538);
  nand n41542(x41542, x41541, x41540);
  nand n41544(x41544, x41536, x41540);
  nand n41545(x41545, x40357, x40359);
  nand n41546(x41546, x40356, x40358);
  nand n41547(x41547, x41546, x41545);
  nand n41549(x41549, x40361, x41548);
  nand n41550(x41550, x40360, x41547);
  nand n41551(x41551, x41550, x41549);
  nand n41553(x41553, x41545, x41549);
  nand n41554(x41554, x40363, x40365);
  nand n41555(x41555, x40362, x40364);
  nand n41556(x41556, x41555, x41554);
  nand n41558(x41558, x40367, x41557);
  nand n41559(x41559, x40366, x41556);
  nand n41560(x41560, x41559, x41558);
  nand n41562(x41562, x41554, x41558);
  nand n41563(x41563, x40369, x40371);
  nand n41564(x41564, x40368, x40370);
  nand n41565(x41565, x41564, x41563);
  nand n41567(x41567, x40373, x41566);
  nand n41568(x41568, x40372, x41565);
  nand n41569(x41569, x41568, x41567);
  nand n41571(x41571, x41563, x41567);
  nand n41572(x41572, x40375, x40377);
  nand n41573(x41573, x40374, x40376);
  nand n41574(x41574, x41573, x41572);
  nand n41576(x41576, x40379, x41575);
  nand n41577(x41577, x40378, x41574);
  nand n41578(x41578, x41577, x41576);
  nand n41580(x41580, x41572, x41576);
  nand n41581(x41581, x40381, x40383);
  nand n41582(x41582, x40380, x40382);
  nand n41583(x41583, x41582, x41581);
  nand n41584(x41584, x40385, x40387);
  nand n41585(x41585, x40384, x40386);
  nand n41586(x41586, x41585, x41584);
  nand n41588(x41588, x40389, x41587);
  nand n41589(x41589, x40388, x41586);
  nand n41590(x41590, x41589, x41588);
  nand n41591(x41591, x41584, x41588);
  nand n41592(x41592, x40391, x40393);
  nand n41593(x41593, x40390, x40392);
  nand n41594(x41594, x41593, x41592);
  nand n41596(x41596, x40395, x41595);
  nand n41597(x41597, x40394, x41594);
  nand n41598(x41598, x41597, x41596);
  nand n41600(x41600, x41592, x41596);
  nand n41601(x41601, x40397, x40399);
  nand n41602(x41602, x40396, x40398);
  nand n41603(x41603, x41602, x41601);
  nand n41605(x41605, x40401, x41604);
  nand n41606(x41606, x40400, x41603);
  nand n41607(x41607, x41606, x41605);
  nand n41609(x41609, x41601, x41605);
  nand n41610(x41610, x40403, x40405);
  nand n41611(x41611, x40402, x40404);
  nand n41612(x41612, x41611, x41610);
  nand n41614(x41614, x40407, x41613);
  nand n41615(x41615, x40406, x41612);
  nand n41616(x41616, x41615, x41614);
  nand n41618(x41618, x41610, x41614);
  nand n41619(x41619, x40409, x40411);
  nand n41620(x41620, x40408, x40410);
  nand n41621(x41621, x41620, x41619);
  nand n41623(x41623, x40413, x41622);
  nand n41624(x41624, x40412, x41621);
  nand n41625(x41625, x41624, x41623);
  nand n41627(x41627, x41619, x41623);
  nand n41628(x41628, x40415, x40417);
  nand n41629(x41629, x40414, x40416);
  nand n41630(x41630, x41629, x41628);
  nand n41632(x41632, x40419, x41631);
  nand n41633(x41633, x40418, x41630);
  nand n41634(x41634, x41633, x41632);
  nand n41636(x41636, x41628, x41632);
  nand n41637(x41637, x40421, x40423);
  nand n41638(x41638, x40420, x40422);
  nand n41639(x41639, x41638, x41637);
  nand n41641(x41641, x40425, x41640);
  nand n41642(x41642, x40424, x41639);
  nand n41643(x41643, x41642, x41641);
  nand n41645(x41645, x41637, x41641);
  nand n41646(x41646, x40427, x40429);
  nand n41647(x41647, x40426, x40428);
  nand n41648(x41648, x41647, x41646);
  nand n41650(x41650, x40431, x41649);
  nand n41651(x41651, x40430, x41648);
  nand n41652(x41652, x41651, x41650);
  nand n41653(x41653, x41646, x41650);
  nand n41654(x41654, x40433, x40435);
  nand n41655(x41655, x40432, x40434);
  nand n41656(x41656, x41655, x41654);
  nand n41658(x41658, x40437, x41657);
  nand n41659(x41659, x40436, x41656);
  nand n41660(x41660, x41659, x41658);
  nand n41662(x41662, x41654, x41658);
  nand n41663(x41663, x40439, x40441);
  nand n41664(x41664, x40438, x40440);
  nand n41665(x41665, x41664, x41663);
  nand n41667(x41667, x40443, x41666);
  nand n41668(x41668, x40442, x41665);
  nand n41669(x41669, x41668, x41667);
  nand n41671(x41671, x41663, x41667);
  nand n41672(x41672, x40445, x40447);
  nand n41673(x41673, x40444, x40446);
  nand n41674(x41674, x41673, x41672);
  nand n41676(x41676, x40449, x41675);
  nand n41677(x41677, x40448, x41674);
  nand n41678(x41678, x41677, x41676);
  nand n41680(x41680, x41672, x41676);
  nand n41681(x41681, x40451, x40453);
  nand n41682(x41682, x40450, x40452);
  nand n41683(x41683, x41682, x41681);
  nand n41685(x41685, x40455, x41684);
  nand n41686(x41686, x40454, x41683);
  nand n41687(x41687, x41686, x41685);
  nand n41689(x41689, x41681, x41685);
  nand n41690(x41690, x40457, x40459);
  nand n41691(x41691, x40456, x40458);
  nand n41692(x41692, x41691, x41690);
  nand n41694(x41694, x40461, x41693);
  nand n41695(x41695, x40460, x41692);
  nand n41696(x41696, x41695, x41694);
  nand n41698(x41698, x41690, x41694);
  nand n41699(x41699, x40463, x40465);
  nand n41700(x41700, x40462, x40464);
  nand n41701(x41701, x41700, x41699);
  nand n41703(x41703, x40467, x41702);
  nand n41704(x41704, x40466, x41701);
  nand n41705(x41705, x41704, x41703);
  nand n41707(x41707, x41699, x41703);
  nand n41708(x41708, x40470, x40472);
  nand n41709(x41709, x40469, x40471);
  nand n41710(x41710, x41709, x41708);
  nand n41712(x41712, x40474, x41711);
  nand n41713(x41713, x40473, x41710);
  nand n41714(x41714, x41713, x41712);
  nand n41715(x41715, x41708, x41712);
  nand n41716(x41716, x40476, x40478);
  nand n41717(x41717, x40475, x40477);
  nand n41718(x41718, x41717, x41716);
  nand n41720(x41720, x40480, x41719);
  nand n41721(x41721, x40479, x41718);
  nand n41722(x41722, x41721, x41720);
  nand n41724(x41724, x41716, x41720);
  nand n41725(x41725, x40482, x40484);
  nand n41726(x41726, x40481, x40483);
  nand n41727(x41727, x41726, x41725);
  nand n41729(x41729, x40486, x41728);
  nand n41730(x41730, x40485, x41727);
  nand n41731(x41731, x41730, x41729);
  nand n41733(x41733, x41725, x41729);
  nand n41734(x41734, x40488, x40490);
  nand n41735(x41735, x40487, x40489);
  nand n41736(x41736, x41735, x41734);
  nand n41738(x41738, x40492, x41737);
  nand n41739(x41739, x40491, x41736);
  nand n41740(x41740, x41739, x41738);
  nand n41742(x41742, x41734, x41738);
  nand n41743(x41743, x40494, x40496);
  nand n41744(x41744, x40493, x40495);
  nand n41745(x41745, x41744, x41743);
  nand n41747(x41747, x40498, x41746);
  nand n41748(x41748, x40497, x41745);
  nand n41749(x41749, x41748, x41747);
  nand n41751(x41751, x41743, x41747);
  nand n41752(x41752, x40500, x40502);
  nand n41753(x41753, x40499, x40501);
  nand n41754(x41754, x41753, x41752);
  nand n41756(x41756, x40504, x41755);
  nand n41757(x41757, x40503, x41754);
  nand n41758(x41758, x41757, x41756);
  nand n41760(x41760, x41752, x41756);
  nand n41761(x41761, x40506, x40508);
  nand n41762(x41762, x40505, x40507);
  nand n41763(x41763, x41762, x41761);
  nand n41765(x41765, x40510, x41764);
  nand n41766(x41766, x40509, x41763);
  nand n41767(x41767, x41766, x41765);
  nand n41769(x41769, x41761, x41765);
  nand n41770(x41770, x40512, x40514);
  nand n41771(x41771, x40511, x40513);
  nand n41772(x41772, x41771, x41770);
  nand n41773(x41773, x40516, x40518);
  nand n41774(x41774, x40515, x40517);
  nand n41775(x41775, x41774, x41773);
  nand n41777(x41777, x40520, x41776);
  nand n41778(x41778, x40519, x41775);
  nand n41779(x41779, x41778, x41777);
  nand n41780(x41780, x41773, x41777);
  nand n41781(x41781, x40522, x40524);
  nand n41782(x41782, x40521, x40523);
  nand n41783(x41783, x41782, x41781);
  nand n41785(x41785, x40526, x41784);
  nand n41786(x41786, x40525, x41783);
  nand n41787(x41787, x41786, x41785);
  nand n41789(x41789, x41781, x41785);
  nand n41790(x41790, x40528, x40530);
  nand n41791(x41791, x40527, x40529);
  nand n41792(x41792, x41791, x41790);
  nand n41794(x41794, x40532, x41793);
  nand n41795(x41795, x40531, x41792);
  nand n41796(x41796, x41795, x41794);
  nand n41798(x41798, x41790, x41794);
  nand n41799(x41799, x40534, x40536);
  nand n41800(x41800, x40533, x40535);
  nand n41801(x41801, x41800, x41799);
  nand n41803(x41803, x40538, x41802);
  nand n41804(x41804, x40537, x41801);
  nand n41805(x41805, x41804, x41803);
  nand n41807(x41807, x41799, x41803);
  nand n41808(x41808, x40540, x40542);
  nand n41809(x41809, x40539, x40541);
  nand n41810(x41810, x41809, x41808);
  nand n41812(x41812, x40544, x41811);
  nand n41813(x41813, x40543, x41810);
  nand n41814(x41814, x41813, x41812);
  nand n41816(x41816, x41808, x41812);
  nand n41817(x41817, x40546, x40548);
  nand n41818(x41818, x40545, x40547);
  nand n41819(x41819, x41818, x41817);
  nand n41821(x41821, x40550, x41820);
  nand n41822(x41822, x40549, x41819);
  nand n41823(x41823, x41822, x41821);
  nand n41825(x41825, x41817, x41821);
  nand n41826(x41826, x40552, x40554);
  nand n41827(x41827, x40551, x40553);
  nand n41828(x41828, x41827, x41826);
  nand n41830(x41830, x40556, x41829);
  nand n41831(x41831, x40555, x41828);
  nand n41832(x41832, x41831, x41830);
  nand n41834(x41834, x41826, x41830);
  nand n41835(x41835, x40558, x40560);
  nand n41836(x41836, x40557, x40559);
  nand n41837(x41837, x41836, x41835);
  nand n41839(x41839, x40562, x41838);
  nand n41840(x41840, x40561, x41837);
  nand n41841(x41841, x41840, x41839);
  nand n41842(x41842, x41835, x41839);
  nand n41843(x41843, x40564, x40566);
  nand n41844(x41844, x40563, x40565);
  nand n41845(x41845, x41844, x41843);
  nand n41847(x41847, x40568, x41846);
  nand n41848(x41848, x40567, x41845);
  nand n41849(x41849, x41848, x41847);
  nand n41850(x41850, x41843, x41847);
  nand n41851(x41851, x40570, x40572);
  nand n41852(x41852, x40569, x40571);
  nand n41853(x41853, x41852, x41851);
  nand n41855(x41855, x40574, x41854);
  nand n41856(x41856, x40573, x41853);
  nand n41857(x41857, x41856, x41855);
  nand n41859(x41859, x41851, x41855);
  nand n41860(x41860, x40576, x40578);
  nand n41861(x41861, x40575, x40577);
  nand n41862(x41862, x41861, x41860);
  nand n41864(x41864, x40580, x41863);
  nand n41865(x41865, x40579, x41862);
  nand n41866(x41866, x41865, x41864);
  nand n41868(x41868, x41860, x41864);
  nand n41869(x41869, x40582, x40584);
  nand n41870(x41870, x40581, x40583);
  nand n41871(x41871, x41870, x41869);
  nand n41873(x41873, x40586, x41872);
  nand n41874(x41874, x40585, x41871);
  nand n41875(x41875, x41874, x41873);
  nand n41877(x41877, x41869, x41873);
  nand n41878(x41878, x40588, x40590);
  nand n41879(x41879, x40587, x40589);
  nand n41880(x41880, x41879, x41878);
  nand n41882(x41882, x40592, x41881);
  nand n41883(x41883, x40591, x41880);
  nand n41884(x41884, x41883, x41882);
  nand n41886(x41886, x41878, x41882);
  nand n41887(x41887, x40594, x40596);
  nand n41888(x41888, x40593, x40595);
  nand n41889(x41889, x41888, x41887);
  nand n41891(x41891, x40598, x41890);
  nand n41892(x41892, x40597, x41889);
  nand n41893(x41893, x41892, x41891);
  nand n41895(x41895, x41887, x41891);
  nand n41896(x41896, x40600, x40602);
  nand n41897(x41897, x40599, x40601);
  nand n41898(x41898, x41897, x41896);
  nand n41900(x41900, x40604, x41899);
  nand n41901(x41901, x40603, x41898);
  nand n41902(x41902, x41901, x41900);
  nand n41904(x41904, x41896, x41900);
  nand n41905(x41905, x40606, x40608);
  nand n41906(x41906, x40605, x40607);
  nand n41907(x41907, x41906, x41905);
  nand n41909(x41909, x40610, x41908);
  nand n41910(x41910, x40609, x41907);
  nand n41911(x41911, x41910, x41909);
  nand n41913(x41913, x41905, x41909);
  nand n41914(x41914, x40613, x40615);
  nand n41915(x41915, x40612, x40614);
  nand n41916(x41916, x41915, x41914);
  nand n41918(x41918, x40617, x41917);
  nand n41919(x41919, x40616, x41916);
  nand n41920(x41920, x41919, x41918);
  nand n41921(x41921, x41914, x41918);
  nand n41922(x41922, x40619, x40621);
  nand n41923(x41923, x40618, x40620);
  nand n41924(x41924, x41923, x41922);
  nand n41926(x41926, x40623, x41925);
  nand n41927(x41927, x40622, x41924);
  nand n41928(x41928, x41927, x41926);
  nand n41930(x41930, x41922, x41926);
  nand n41931(x41931, x40625, x40627);
  nand n41932(x41932, x40624, x40626);
  nand n41933(x41933, x41932, x41931);
  nand n41935(x41935, x40629, x41934);
  nand n41936(x41936, x40628, x41933);
  nand n41937(x41937, x41936, x41935);
  nand n41939(x41939, x41931, x41935);
  nand n41940(x41940, x40631, x40633);
  nand n41941(x41941, x40630, x40632);
  nand n41942(x41942, x41941, x41940);
  nand n41944(x41944, x40635, x41943);
  nand n41945(x41945, x40634, x41942);
  nand n41946(x41946, x41945, x41944);
  nand n41948(x41948, x41940, x41944);
  nand n41949(x41949, x40637, x40639);
  nand n41950(x41950, x40636, x40638);
  nand n41951(x41951, x41950, x41949);
  nand n41953(x41953, x40641, x41952);
  nand n41954(x41954, x40640, x41951);
  nand n41955(x41955, x41954, x41953);
  nand n41957(x41957, x41949, x41953);
  nand n41958(x41958, x40643, x40645);
  nand n41959(x41959, x40642, x40644);
  nand n41960(x41960, x41959, x41958);
  nand n41962(x41962, x40647, x41961);
  nand n41963(x41963, x40646, x41960);
  nand n41964(x41964, x41963, x41962);
  nand n41966(x41966, x41958, x41962);
  nand n41967(x41967, x40649, x40651);
  nand n41968(x41968, x40648, x40650);
  nand n41969(x41969, x41968, x41967);
  nand n41971(x41971, x40653, x41970);
  nand n41972(x41972, x40652, x41969);
  nand n41973(x41973, x41972, x41971);
  nand n41975(x41975, x41967, x41971);
  nand n41976(x41976, x40655, x40657);
  nand n41977(x41977, x40654, x40656);
  nand n41978(x41978, x41977, x41976);
  nand n41980(x41980, x40659, x41979);
  nand n41981(x41981, x40658, x41978);
  nand n41982(x41982, x41981, x41980);
  nand n41984(x41984, x41976, x41980);
  nand n41985(x41985, x40661, x40663);
  nand n41986(x41986, x40660, x40662);
  nand n41987(x41987, x41986, x41985);
  nand n41988(x41988, x40665, x40667);
  nand n41989(x41989, x40664, x40666);
  nand n41990(x41990, x41989, x41988);
  nand n41992(x41992, x40669, x41991);
  nand n41993(x41993, x40668, x41990);
  nand n41994(x41994, x41993, x41992);
  nand n41995(x41995, x41988, x41992);
  nand n41996(x41996, x40671, x40673);
  nand n41997(x41997, x40670, x40672);
  nand n41998(x41998, x41997, x41996);
  nand n42000(x42000, x40675, x41999);
  nand n42001(x42001, x40674, x41998);
  nand n42002(x42002, x42001, x42000);
  nand n42004(x42004, x41996, x42000);
  nand n42005(x42005, x40677, x40679);
  nand n42006(x42006, x40676, x40678);
  nand n42007(x42007, x42006, x42005);
  nand n42009(x42009, x40681, x42008);
  nand n42010(x42010, x40680, x42007);
  nand n42011(x42011, x42010, x42009);
  nand n42013(x42013, x42005, x42009);
  nand n42014(x42014, x40683, x40685);
  nand n42015(x42015, x40682, x40684);
  nand n42016(x42016, x42015, x42014);
  nand n42018(x42018, x40687, x42017);
  nand n42019(x42019, x40686, x42016);
  nand n42020(x42020, x42019, x42018);
  nand n42022(x42022, x42014, x42018);
  nand n42023(x42023, x40689, x40691);
  nand n42024(x42024, x40688, x40690);
  nand n42025(x42025, x42024, x42023);
  nand n42027(x42027, x40693, x42026);
  nand n42028(x42028, x40692, x42025);
  nand n42029(x42029, x42028, x42027);
  nand n42031(x42031, x42023, x42027);
  nand n42032(x42032, x40695, x40697);
  nand n42033(x42033, x40694, x40696);
  nand n42034(x42034, x42033, x42032);
  nand n42036(x42036, x40699, x42035);
  nand n42037(x42037, x40698, x42034);
  nand n42038(x42038, x42037, x42036);
  nand n42040(x42040, x42032, x42036);
  nand n42041(x42041, x40701, x40703);
  nand n42042(x42042, x40700, x40702);
  nand n42043(x42043, x42042, x42041);
  nand n42045(x42045, x40705, x42044);
  nand n42046(x42046, x40704, x42043);
  nand n42047(x42047, x42046, x42045);
  nand n42049(x42049, x42041, x42045);
  nand n42050(x42050, x40707, x40709);
  nand n42051(x42051, x40706, x40708);
  nand n42052(x42052, x42051, x42050);
  nand n42054(x42054, x40711, x42053);
  nand n42055(x42055, x40710, x42052);
  nand n42056(x42056, x42055, x42054);
  nand n42058(x42058, x42050, x42054);
  nand n42059(x42059, x40713, x40715);
  nand n42060(x42060, x40712, x40714);
  nand n42061(x42061, x42060, x42059);
  nand n42063(x42063, x40717, x42062);
  nand n42064(x42064, x40716, x42061);
  nand n42065(x42065, x42064, x42063);
  nand n42067(x42067, x42059, x42063);
  nand n42068(x42068, x40719, x40721);
  nand n42069(x42069, x40718, x40720);
  nand n42070(x42070, x42069, x42068);
  nand n42072(x42072, x40723, x42071);
  nand n42073(x42073, x40722, x42070);
  nand n42074(x42074, x42073, x42072);
  nand n42075(x42075, x42068, x42072);
  nand n42076(x42076, x40725, x40727);
  nand n42077(x42077, x40724, x40726);
  nand n42078(x42078, x42077, x42076);
  nand n42080(x42080, x40729, x42079);
  nand n42081(x42081, x40728, x42078);
  nand n42082(x42082, x42081, x42080);
  nand n42084(x42084, x42076, x42080);
  nand n42085(x42085, x40731, x40733);
  nand n42086(x42086, x40730, x40732);
  nand n42087(x42087, x42086, x42085);
  nand n42089(x42089, x40735, x42088);
  nand n42090(x42090, x40734, x42087);
  nand n42091(x42091, x42090, x42089);
  nand n42093(x42093, x42085, x42089);
  nand n42094(x42094, x40737, x40739);
  nand n42095(x42095, x40736, x40738);
  nand n42096(x42096, x42095, x42094);
  nand n42098(x42098, x40741, x42097);
  nand n42099(x42099, x40740, x42096);
  nand n42100(x42100, x42099, x42098);
  nand n42102(x42102, x42094, x42098);
  nand n42103(x42103, x40743, x40745);
  nand n42104(x42104, x40742, x40744);
  nand n42105(x42105, x42104, x42103);
  nand n42107(x42107, x40747, x42106);
  nand n42108(x42108, x40746, x42105);
  nand n42109(x42109, x42108, x42107);
  nand n42111(x42111, x42103, x42107);
  nand n42112(x42112, x40749, x40751);
  nand n42113(x42113, x40748, x40750);
  nand n42114(x42114, x42113, x42112);
  nand n42116(x42116, x40753, x42115);
  nand n42117(x42117, x40752, x42114);
  nand n42118(x42118, x42117, x42116);
  nand n42120(x42120, x42112, x42116);
  nand n42121(x42121, x40755, x40757);
  nand n42122(x42122, x40754, x40756);
  nand n42123(x42123, x42122, x42121);
  nand n42125(x42125, x40759, x42124);
  nand n42126(x42126, x40758, x42123);
  nand n42127(x42127, x42126, x42125);
  nand n42129(x42129, x42121, x42125);
  nand n42130(x42130, x40761, x40763);
  nand n42131(x42131, x40760, x40762);
  nand n42132(x42132, x42131, x42130);
  nand n42134(x42134, x40765, x42133);
  nand n42135(x42135, x40764, x42132);
  nand n42136(x42136, x42135, x42134);
  nand n42138(x42138, x42130, x42134);
  nand n42139(x42139, x40767, x40769);
  nand n42140(x42140, x40766, x40768);
  nand n42141(x42141, x42140, x42139);
  nand n42143(x42143, x40771, x42142);
  nand n42144(x42144, x40770, x42141);
  nand n42145(x42145, x42144, x42143);
  nand n42147(x42147, x42139, x42143);
  nand n42148(x42148, x40774, x40776);
  nand n42149(x42149, x40773, x40775);
  nand n42150(x42150, x42149, x42148);
  nand n42152(x42152, x40778, x42151);
  nand n42153(x42153, x40777, x42150);
  nand n42154(x42154, x42153, x42152);
  nand n42155(x42155, x42148, x42152);
  nand n42156(x42156, x40780, x40782);
  nand n42157(x42157, x40779, x40781);
  nand n42158(x42158, x42157, x42156);
  nand n42160(x42160, x40784, x42159);
  nand n42161(x42161, x40783, x42158);
  nand n42162(x42162, x42161, x42160);
  nand n42164(x42164, x42156, x42160);
  nand n42165(x42165, x40786, x40788);
  nand n42166(x42166, x40785, x40787);
  nand n42167(x42167, x42166, x42165);
  nand n42169(x42169, x40790, x42168);
  nand n42170(x42170, x40789, x42167);
  nand n42171(x42171, x42170, x42169);
  nand n42173(x42173, x42165, x42169);
  nand n42174(x42174, x40792, x40794);
  nand n42175(x42175, x40791, x40793);
  nand n42176(x42176, x42175, x42174);
  nand n42178(x42178, x40796, x42177);
  nand n42179(x42179, x40795, x42176);
  nand n42180(x42180, x42179, x42178);
  nand n42182(x42182, x42174, x42178);
  nand n42183(x42183, x40798, x40800);
  nand n42184(x42184, x40797, x40799);
  nand n42185(x42185, x42184, x42183);
  nand n42187(x42187, x40802, x42186);
  nand n42188(x42188, x40801, x42185);
  nand n42189(x42189, x42188, x42187);
  nand n42191(x42191, x42183, x42187);
  nand n42192(x42192, x40804, x40806);
  nand n42193(x42193, x40803, x40805);
  nand n42194(x42194, x42193, x42192);
  nand n42196(x42196, x40808, x42195);
  nand n42197(x42197, x40807, x42194);
  nand n42198(x42198, x42197, x42196);
  nand n42200(x42200, x42192, x42196);
  nand n42201(x42201, x40810, x40812);
  nand n42202(x42202, x40809, x40811);
  nand n42203(x42203, x42202, x42201);
  nand n42205(x42205, x40814, x42204);
  nand n42206(x42206, x40813, x42203);
  nand n42207(x42207, x42206, x42205);
  nand n42209(x42209, x42201, x42205);
  nand n42210(x42210, x40816, x40818);
  nand n42211(x42211, x40815, x40817);
  nand n42212(x42212, x42211, x42210);
  nand n42214(x42214, x40820, x42213);
  nand n42215(x42215, x40819, x42212);
  nand n42216(x42216, x42215, x42214);
  nand n42218(x42218, x42210, x42214);
  nand n42219(x42219, x40822, x40824);
  nand n42220(x42220, x40821, x40823);
  nand n42221(x42221, x42220, x42219);
  nand n42223(x42223, x40826, x42222);
  nand n42224(x42224, x40825, x42221);
  nand n42225(x42225, x42224, x42223);
  nand n42227(x42227, x42219, x42223);
  nand n42228(x42228, x40828, x40830);
  nand n42229(x42229, x40827, x40829);
  nand n42230(x42230, x42229, x42228);
  nand n42231(x42231, x40832, x40834);
  nand n42232(x42232, x40831, x40833);
  nand n42233(x42233, x42232, x42231);
  nand n42235(x42235, x40836, x42234);
  nand n42236(x42236, x40835, x42233);
  nand n42237(x42237, x42236, x42235);
  nand n42239(x42239, x42231, x42235);
  nand n42240(x42240, x40838, x40840);
  nand n42241(x42241, x40837, x40839);
  nand n42242(x42242, x42241, x42240);
  nand n42244(x42244, x40842, x42243);
  nand n42245(x42245, x40841, x42242);
  nand n42246(x42246, x42245, x42244);
  nand n42248(x42248, x42240, x42244);
  nand n42249(x42249, x40844, x40846);
  nand n42250(x42250, x40843, x40845);
  nand n42251(x42251, x42250, x42249);
  nand n42253(x42253, x40848, x42252);
  nand n42254(x42254, x40847, x42251);
  nand n42255(x42255, x42254, x42253);
  nand n42257(x42257, x42249, x42253);
  nand n42258(x42258, x40850, x40852);
  nand n42259(x42259, x40849, x40851);
  nand n42260(x42260, x42259, x42258);
  nand n42262(x42262, x40854, x42261);
  nand n42263(x42263, x40853, x42260);
  nand n42264(x42264, x42263, x42262);
  nand n42266(x42266, x42258, x42262);
  nand n42267(x42267, x40856, x40858);
  nand n42268(x42268, x40855, x40857);
  nand n42269(x42269, x42268, x42267);
  nand n42271(x42271, x40860, x42270);
  nand n42272(x42272, x40859, x42269);
  nand n42273(x42273, x42272, x42271);
  nand n42275(x42275, x42267, x42271);
  nand n42276(x42276, x40862, x40864);
  nand n42277(x42277, x40861, x40863);
  nand n42278(x42278, x42277, x42276);
  nand n42280(x42280, x40866, x42279);
  nand n42281(x42281, x40865, x42278);
  nand n42282(x42282, x42281, x42280);
  nand n42284(x42284, x42276, x42280);
  nand n42285(x42285, x40868, x40870);
  nand n42286(x42286, x40867, x40869);
  nand n42287(x42287, x42286, x42285);
  nand n42289(x42289, x40872, x42288);
  nand n42290(x42290, x40871, x42287);
  nand n42291(x42291, x42290, x42289);
  nand n42293(x42293, x42285, x42289);
  nand n42294(x42294, x40874, x40876);
  nand n42295(x42295, x40873, x40875);
  nand n42296(x42296, x42295, x42294);
  nand n42298(x42298, x40878, x42297);
  nand n42299(x42299, x40877, x42296);
  nand n42300(x42300, x42299, x42298);
  nand n42302(x42302, x42294, x42298);
  nand n42303(x42303, x40880, x40882);
  nand n42304(x42304, x40879, x40881);
  nand n42305(x42305, x42304, x42303);
  nand n42307(x42307, x40884, x42306);
  nand n42308(x42308, x40883, x42305);
  nand n42309(x42309, x42308, x42307);
  nand n42311(x42311, x42303, x42307);
  nand n42312(x42312, x40886, x40888);
  nand n42313(x42313, x40885, x40887);
  nand n42314(x42314, x42313, x42312);
  nand n42316(x42316, x40890, x42315);
  nand n42317(x42317, x40889, x42314);
  nand n42318(x42318, x42317, x42316);
  nand n42320(x42320, x42312, x42316);
  nand n42321(x42321, x40892, x40894);
  nand n42322(x42322, x40891, x40893);
  nand n42323(x42323, x42322, x42321);
  nand n42325(x42325, x40896, x42324);
  nand n42326(x42326, x40895, x42323);
  nand n42327(x42327, x42326, x42325);
  nand n42329(x42329, x42321, x42325);
  nand n42330(x42330, x40898, x40900);
  nand n42331(x42331, x40897, x40899);
  nand n42332(x42332, x42331, x42330);
  nand n42334(x42334, x40902, x42333);
  nand n42335(x42335, x40901, x42332);
  nand n42336(x42336, x42335, x42334);
  nand n42338(x42338, x42330, x42334);
  nand n42339(x42339, x40904, x40906);
  nand n42340(x42340, x40903, x40905);
  nand n42341(x42341, x42340, x42339);
  nand n42343(x42343, x40908, x42342);
  nand n42344(x42344, x40907, x42341);
  nand n42345(x42345, x42344, x42343);
  nand n42347(x42347, x42339, x42343);
  nand n42348(x42348, x40910, x40912);
  nand n42349(x42349, x40909, x40911);
  nand n42350(x42350, x42349, x42348);
  nand n42352(x42352, x40914, x42351);
  nand n42353(x42353, x40913, x42350);
  nand n42354(x42354, x42353, x42352);
  nand n42356(x42356, x42348, x42352);
  nand n42357(x42357, x40916, x40918);
  nand n42358(x42358, x40915, x40917);
  nand n42359(x42359, x42358, x42357);
  nand n42361(x42361, x40920, x42360);
  nand n42362(x42362, x40919, x42359);
  nand n42363(x42363, x42362, x42361);
  nand n42365(x42365, x42357, x42361);
  nand n42366(x42366, x40922, x40924);
  nand n42367(x42367, x40921, x40923);
  nand n42368(x42368, x42367, x42366);
  nand n42370(x42370, x40926, x42369);
  nand n42371(x42371, x40925, x42368);
  nand n42372(x42372, x42371, x42370);
  nand n42374(x42374, x42366, x42370);
  nand n42375(x42375, x40928, x40930);
  nand n42376(x42376, x40927, x40929);
  nand n42377(x42377, x42376, x42375);
  nand n42379(x42379, x40932, x42378);
  nand n42380(x42380, x40931, x42377);
  nand n42381(x42381, x42380, x42379);
  nand n42383(x42383, x42375, x42379);
  nand n42384(x42384, x40934, x40936);
  nand n42385(x42385, x40933, x40935);
  nand n42386(x42386, x42385, x42384);
  nand n42388(x42388, x40938, x42387);
  nand n42389(x42389, x40937, x42386);
  nand n42390(x42390, x42389, x42388);
  nand n42392(x42392, x42384, x42388);
  nand n42393(x42393, x40940, x40942);
  nand n42394(x42394, x40939, x40941);
  nand n42395(x42395, x42394, x42393);
  nand n42397(x42397, x40944, x42396);
  nand n42398(x42398, x40943, x42395);
  nand n42399(x42399, x42398, x42397);
  nand n42401(x42401, x42393, x42397);
  nand n42402(x42402, x40946, x40948);
  nand n42403(x42403, x40945, x40947);
  nand n42404(x42404, x42403, x42402);
  nand n42406(x42406, x40950, x42405);
  nand n42407(x42407, x40949, x42404);
  nand n42408(x42408, x42407, x42406);
  nand n42410(x42410, x42402, x42406);
  nand n42411(x42411, x40953, x40955);
  nand n42412(x42412, x40952, x40954);
  nand n42413(x42413, x42412, x42411);
  nand n42415(x42415, x40957, x42414);
  nand n42416(x42416, x40956, x42413);
  nand n42417(x42417, x42416, x42415);
  nand n42419(x42419, x40959, x40961);
  nand n42420(x42420, x40958, x40960);
  nand n42421(x42421, x42420, x42419);
  nand n42423(x42423, x40963, x42422);
  nand n42424(x42424, x40962, x42421);
  nand n42425(x42425, x42424, x42423);
  nand n42427(x42427, x40965, x40967);
  nand n42428(x42428, x40964, x40966);
  nand n42429(x42429, x42428, x42427);
  nand n42431(x42431, x40969, x42430);
  nand n42432(x42432, x40968, x42429);
  nand n42433(x42433, x42432, x42431);
  nand n42435(x42435, x40971, x40973);
  nand n42436(x42436, x40970, x40972);
  nand n42437(x42437, x42436, x42435);
  nand n42439(x42439, x40975, x42438);
  nand n42440(x42440, x40974, x42437);
  nand n42441(x42441, x42440, x42439);
  nand n42443(x42443, x40977, x40979);
  nand n42444(x42444, x40976, x40978);
  nand n42445(x42445, x42444, x42443);
  nand n42447(x42447, x40981, x42446);
  nand n42448(x42448, x40980, x42445);
  nand n42449(x42449, x42448, x42447);
  nand n42451(x42451, x40983, x40985);
  nand n42452(x42452, x40982, x40984);
  nand n42453(x42453, x42452, x42451);
  nand n42455(x42455, x40987, x42454);
  nand n42456(x42456, x40986, x42453);
  nand n42457(x42457, x42456, x42455);
  nand n42459(x42459, x40989, x40991);
  nand n42460(x42460, x40988, x40990);
  nand n42461(x42461, x42460, x42459);
  nand n42463(x42463, x40993, x42462);
  nand n42464(x42464, x40992, x42461);
  nand n42465(x42465, x42464, x42463);
  nand n42467(x42467, x40995, x40997);
  nand n42468(x42468, x40994, x40996);
  nand n42469(x42469, x42468, x42467);
  nand n42471(x42471, x40999, x42470);
  nand n42472(x42472, x40998, x42469);
  nand n42473(x42473, x42472, x42471);
  nand n42475(x42475, x41001, x41003);
  nand n42476(x42476, x41000, x41002);
  nand n42477(x42477, x42476, x42475);
  nand n42479(x42479, x41005, x42478);
  nand n42480(x42480, x41004, x42477);
  nand n42481(x42481, x42480, x42479);
  nand n42483(x42483, x41007, x41009);
  nand n42484(x42484, x41006, x41008);
  nand n42485(x42485, x42484, x42483);
  nand n42487(x42487, x41011, x42486);
  nand n42488(x42488, x41010, x42485);
  nand n42489(x42489, x42488, x42487);
  nand n42491(x42491, x41013, x41015);
  nand n42492(x42492, x41012, x41014);
  nand n42493(x42493, x42492, x42491);
  nand n42497(x42497, x41042, x84939);
  nand n42499(x42499, x42498, x41043);
  nand n42500(x42500, x42499, x42497);
  nand n42501(x42501, x41053, x41061);
  nand n42504(x42504, x42503, x42502);
  nand n42505(x42505, x42504, x42501);
  nand n42506(x42506, x41077, x84940);
  nand n42507(x42507, x41076, x40023);
  nand n42508(x42508, x42507, x42506);
  nand n42509(x42509, x41069, x41078);
  nand n42512(x42512, x42511, x42510);
  nand n42513(x42513, x42512, x42509);
  nand n42514(x42514, x41094, x84941);
  nand n42515(x42515, x41093, x41098);
  nand n42516(x42516, x42515, x42514);
  nand n42517(x42517, x41086, x41095);
  nand n42520(x42520, x42519, x42518);
  nand n42521(x42521, x42520, x42517);
  nand n42523(x42523, x84942, x42522);
  nand n42524(x42524, x41096, x42521);
  nand n42525(x42525, x42524, x42523);
  nand n42526(x42526, x42517, x42523);
  nand n42527(x42527, x41114, x41123);
  nand n42528(x42528, x41113, x41122);
  nand n42529(x42529, x42528, x42527);
  nand n42530(x42530, x41106, x41115);
  nand n42533(x42533, x42532, x42531);
  nand n42534(x42534, x42533, x42530);
  nand n42536(x42536, x41124, x42535);
  nand n42538(x42538, x42537, x42534);
  nand n42539(x42539, x42538, x42536);
  nand n42540(x42540, x42530, x42536);
  nand n42541(x42541, x41140, x41149);
  nand n42542(x42542, x41139, x41148);
  nand n42543(x42543, x42542, x42541);
  nand n42545(x42545, x84943, x42544);
  nand n42546(x42546, x40076, x42543);
  nand n42547(x42547, x42546, x42545);
  nand n42549(x42549, x42541, x42545);
  nand n42550(x42550, x41132, x41141);
  nand n42553(x42553, x42552, x42551);
  nand n42554(x42554, x42553, x42550);
  nand n42556(x42556, x41150, x42555);
  nand n42558(x42558, x42557, x42554);
  nand n42559(x42559, x42558, x42556);
  nand n42560(x42560, x42550, x42556);
  nand n42561(x42561, x41166, x41175);
  nand n42562(x42562, x41165, x41174);
  nand n42563(x42563, x42562, x42561);
  nand n42565(x42565, x84944, x42564);
  nand n42566(x42566, x41179, x42563);
  nand n42567(x42567, x42566, x42565);
  nand n42569(x42569, x42561, x42565);
  nand n42570(x42570, x41158, x41167);
  nand n42573(x42573, x42572, x42571);
  nand n42574(x42574, x42573, x42570);
  nand n42576(x42576, x41176, x42575);
  nand n42578(x42578, x42577, x42574);
  nand n42579(x42579, x42578, x42576);
  nand n42580(x42580, x42570, x42576);
  nand n42581(x42581, x41195, x41204);
  nand n42582(x42582, x41194, x41203);
  nand n42583(x42583, x42582, x42581);
  nand n42585(x42585, x41213, x42584);
  nand n42586(x42586, x41212, x42583);
  nand n42587(x42587, x42586, x42585);
  nand n42589(x42589, x42581, x42585);
  nand n42590(x42590, x41187, x41196);
  nand n42593(x42593, x42592, x42591);
  nand n42594(x42594, x42593, x42590);
  nand n42596(x42596, x41205, x42595);
  nand n42598(x42598, x42597, x42594);
  nand n42599(x42599, x42598, x42596);
  nand n42600(x42600, x42590, x42596);
  nand n42602(x42602, x41230, x41239);
  nand n42603(x42603, x41229, x41238);
  nand n42604(x42604, x42603, x42602);
  nand n42606(x42606, x41248, x42605);
  nand n42607(x42607, x41247, x42604);
  nand n42608(x42608, x42607, x42606);
  nand n42610(x42610, x42602, x42606);
  nand n42611(x42611, x41222, x41231);
  nand n42614(x42614, x42613, x42612);
  nand n42615(x42615, x42614, x42611);
  nand n42617(x42617, x41240, x42616);
  nand n42619(x42619, x42618, x42615);
  nand n42620(x42620, x42619, x42617);
  nand n42621(x42621, x42611, x42617);
  nand n42623(x42623, x41265, x41274);
  nand n42624(x42624, x41264, x41273);
  nand n42625(x42625, x42624, x42623);
  nand n42627(x42627, x41283, x42626);
  nand n42628(x42628, x41282, x42625);
  nand n42629(x42629, x42628, x42627);
  nand n42631(x42631, x42623, x42627);
  nand n42632(x42632, x41257, x41266);
  nand n42635(x42635, x42634, x42633);
  nand n42636(x42636, x42635, x42632);
  nand n42638(x42638, x41275, x42637);
  nand n42640(x42640, x42639, x42636);
  nand n42641(x42641, x42640, x42638);
  nand n42642(x42642, x42632, x42638);
  nand n42643(x42643, x41284, x84945);
  nand n42645(x42645, x42644, x41285);
  nand n42646(x42646, x42645, x42643);
  nand n42647(x42647, x41303, x41312);
  nand n42648(x42648, x41302, x41311);
  nand n42649(x42649, x42648, x42647);
  nand n42651(x42651, x41321, x42650);
  nand n42652(x42652, x41320, x42649);
  nand n42653(x42653, x42652, x42651);
  nand n42655(x42655, x42647, x42651);
  nand n42656(x42656, x41295, x41304);
  nand n42659(x42659, x42658, x42657);
  nand n42660(x42660, x42659, x42656);
  nand n42662(x42662, x41313, x42661);
  nand n42664(x42664, x42663, x42660);
  nand n42665(x42665, x42664, x42662);
  nand n42666(x42666, x42656, x42662);
  nand n42667(x42667, x41322, x41330);
  nand n42670(x42670, x42669, x42668);
  nand n42671(x42671, x42670, x42667);
  nand n42672(x42672, x41346, x41355);
  nand n42673(x42673, x41345, x41354);
  nand n42674(x42674, x42673, x42672);
  nand n42676(x42676, x41364, x42675);
  nand n42677(x42677, x41363, x42674);
  nand n42678(x42678, x42677, x42676);
  nand n42680(x42680, x42672, x42676);
  nand n42681(x42681, x41373, x84946);
  nand n42682(x42682, x41372, x40236);
  nand n42683(x42683, x42682, x42681);
  nand n42684(x42684, x41338, x41347);
  nand n42687(x42687, x42686, x42685);
  nand n42688(x42688, x42687, x42684);
  nand n42690(x42690, x41356, x42689);
  nand n42692(x42692, x42691, x42688);
  nand n42693(x42693, x42692, x42690);
  nand n42694(x42694, x42684, x42690);
  nand n42695(x42695, x41365, x41374);
  nand n42698(x42698, x42697, x42696);
  nand n42699(x42699, x42698, x42695);
  nand n42700(x42700, x41390, x41399);
  nand n42701(x42701, x41389, x41398);
  nand n42702(x42702, x42701, x42700);
  nand n42704(x42704, x41408, x42703);
  nand n42705(x42705, x41407, x42702);
  nand n42706(x42706, x42705, x42704);
  nand n42708(x42708, x42700, x42704);
  nand n42709(x42709, x41417, x84947);
  nand n42710(x42710, x41416, x41421);
  nand n42711(x42711, x42710, x42709);
  nand n42712(x42712, x41382, x41391);
  nand n42715(x42715, x42714, x42713);
  nand n42716(x42716, x42715, x42712);
  nand n42718(x42718, x41400, x42717);
  nand n42720(x42720, x42719, x42716);
  nand n42721(x42721, x42720, x42718);
  nand n42722(x42722, x42712, x42718);
  nand n42723(x42723, x41409, x41418);
  nand n42726(x42726, x42725, x42724);
  nand n42727(x42727, x42726, x42723);
  nand n42729(x42729, x84948, x42728);
  nand n42730(x42730, x41419, x42727);
  nand n42731(x42731, x42730, x42729);
  nand n42733(x42733, x42723, x42729);
  nand n42734(x42734, x41437, x41446);
  nand n42735(x42735, x41436, x41445);
  nand n42736(x42736, x42735, x42734);
  nand n42738(x42738, x41455, x42737);
  nand n42739(x42739, x41454, x42736);
  nand n42740(x42740, x42739, x42738);
  nand n42742(x42742, x42734, x42738);
  nand n42743(x42743, x41464, x41473);
  nand n42744(x42744, x41463, x41472);
  nand n42745(x42745, x42744, x42743);
  nand n42746(x42746, x41429, x41438);
  nand n42749(x42749, x42748, x42747);
  nand n42750(x42750, x42749, x42746);
  nand n42752(x42752, x41447, x42751);
  nand n42754(x42754, x42753, x42750);
  nand n42755(x42755, x42754, x42752);
  nand n42756(x42756, x42746, x42752);
  nand n42757(x42757, x41456, x41465);
  nand n42760(x42760, x42759, x42758);
  nand n42761(x42761, x42760, x42757);
  nand n42763(x42763, x41474, x42762);
  nand n42765(x42765, x42764, x42761);
  nand n42766(x42766, x42765, x42763);
  nand n42768(x42768, x42757, x42763);
  nand n42769(x42769, x41490, x41499);
  nand n42770(x42770, x41489, x41498);
  nand n42771(x42771, x42770, x42769);
  nand n42773(x42773, x41508, x42772);
  nand n42774(x42774, x41507, x42771);
  nand n42775(x42775, x42774, x42773);
  nand n42777(x42777, x42769, x42773);
  nand n42778(x42778, x41517, x41526);
  nand n42779(x42779, x41516, x41525);
  nand n42780(x42780, x42779, x42778);
  nand n42782(x42782, x84949, x42781);
  nand n42783(x42783, x40343, x42780);
  nand n42784(x42784, x42783, x42782);
  nand n42785(x42785, x42778, x42782);
  nand n42786(x42786, x41482, x41491);
  nand n42789(x42789, x42788, x42787);
  nand n42790(x42790, x42789, x42786);
  nand n42792(x42792, x41500, x42791);
  nand n42794(x42794, x42793, x42790);
  nand n42795(x42795, x42794, x42792);
  nand n42796(x42796, x42786, x42792);
  nand n42797(x42797, x41509, x41518);
  nand n42800(x42800, x42799, x42798);
  nand n42801(x42801, x42800, x42797);
  nand n42803(x42803, x41527, x42802);
  nand n42805(x42805, x42804, x42801);
  nand n42806(x42806, x42805, x42803);
  nand n42808(x42808, x42797, x42803);
  nand n42809(x42809, x41543, x41552);
  nand n42810(x42810, x41542, x41551);
  nand n42811(x42811, x42810, x42809);
  nand n42813(x42813, x41561, x42812);
  nand n42814(x42814, x41560, x42811);
  nand n42815(x42815, x42814, x42813);
  nand n42817(x42817, x42809, x42813);
  nand n42818(x42818, x41570, x41579);
  nand n42819(x42819, x41569, x41578);
  nand n42820(x42820, x42819, x42818);
  nand n42822(x42822, x84950, x42821);
  nand n42823(x42823, x41583, x42820);
  nand n42824(x42824, x42823, x42822);
  nand n42825(x42825, x42818, x42822);
  nand n42826(x42826, x41535, x41544);
  nand n42829(x42829, x42828, x42827);
  nand n42830(x42830, x42829, x42826);
  nand n42832(x42832, x41553, x42831);
  nand n42834(x42834, x42833, x42830);
  nand n42835(x42835, x42834, x42832);
  nand n42836(x42836, x42826, x42832);
  nand n42837(x42837, x41562, x41571);
  nand n42840(x42840, x42839, x42838);
  nand n42841(x42841, x42840, x42837);
  nand n42843(x42843, x41580, x42842);
  nand n42845(x42845, x42844, x42841);
  nand n42846(x42846, x42845, x42843);
  nand n42848(x42848, x42837, x42843);
  nand n42849(x42849, x41599, x41608);
  nand n42850(x42850, x41598, x41607);
  nand n42851(x42851, x42850, x42849);
  nand n42853(x42853, x41617, x42852);
  nand n42854(x42854, x41616, x42851);
  nand n42855(x42855, x42854, x42853);
  nand n42857(x42857, x42849, x42853);
  nand n42858(x42858, x41626, x41635);
  nand n42859(x42859, x41625, x41634);
  nand n42860(x42860, x42859, x42858);
  nand n42862(x42862, x41644, x42861);
  nand n42863(x42863, x41643, x42860);
  nand n42864(x42864, x42863, x42862);
  nand n42865(x42865, x42858, x42862);
  nand n42866(x42866, x41591, x41600);
  nand n42869(x42869, x42868, x42867);
  nand n42870(x42870, x42869, x42866);
  nand n42872(x42872, x41609, x42871);
  nand n42874(x42874, x42873, x42870);
  nand n42875(x42875, x42874, x42872);
  nand n42876(x42876, x42866, x42872);
  nand n42877(x42877, x41618, x41627);
  nand n42880(x42880, x42879, x42878);
  nand n42881(x42881, x42880, x42877);
  nand n42883(x42883, x41636, x42882);
  nand n42885(x42885, x42884, x42881);
  nand n42886(x42886, x42885, x42883);
  nand n42888(x42888, x42877, x42883);
  nand n42890(x42890, x41661, x41670);
  nand n42891(x42891, x41660, x41669);
  nand n42892(x42892, x42891, x42890);
  nand n42894(x42894, x41679, x42893);
  nand n42895(x42895, x41678, x42892);
  nand n42896(x42896, x42895, x42894);
  nand n42898(x42898, x42890, x42894);
  nand n42899(x42899, x41688, x41697);
  nand n42900(x42900, x41687, x41696);
  nand n42901(x42901, x42900, x42899);
  nand n42903(x42903, x41706, x42902);
  nand n42904(x42904, x41705, x42901);
  nand n42905(x42905, x42904, x42903);
  nand n42907(x42907, x42899, x42903);
  nand n42908(x42908, x41653, x41662);
  nand n42911(x42911, x42910, x42909);
  nand n42912(x42912, x42911, x42908);
  nand n42914(x42914, x41671, x42913);
  nand n42916(x42916, x42915, x42912);
  nand n42917(x42917, x42916, x42914);
  nand n42918(x42918, x42908, x42914);
  nand n42919(x42919, x41680, x41689);
  nand n42922(x42922, x42921, x42920);
  nand n42923(x42923, x42922, x42919);
  nand n42925(x42925, x41698, x42924);
  nand n42927(x42927, x42926, x42923);
  nand n42928(x42928, x42927, x42925);
  nand n42930(x42930, x42919, x42925);
  nand n42932(x42932, x41723, x41732);
  nand n42933(x42933, x41722, x41731);
  nand n42934(x42934, x42933, x42932);
  nand n42936(x42936, x41741, x42935);
  nand n42937(x42937, x41740, x42934);
  nand n42938(x42938, x42937, x42936);
  nand n42940(x42940, x42932, x42936);
  nand n42941(x42941, x41750, x41759);
  nand n42942(x42942, x41749, x41758);
  nand n42943(x42943, x42942, x42941);
  nand n42945(x42945, x41768, x42944);
  nand n42946(x42946, x41767, x42943);
  nand n42947(x42947, x42946, x42945);
  nand n42949(x42949, x42941, x42945);
  nand n42950(x42950, x41715, x41724);
  nand n42953(x42953, x42952, x42951);
  nand n42954(x42954, x42953, x42950);
  nand n42956(x42956, x41733, x42955);
  nand n42958(x42958, x42957, x42954);
  nand n42959(x42959, x42958, x42956);
  nand n42960(x42960, x42950, x42956);
  nand n42961(x42961, x41742, x41751);
  nand n42964(x42964, x42963, x42962);
  nand n42965(x42965, x42964, x42961);
  nand n42967(x42967, x41760, x42966);
  nand n42969(x42969, x42968, x42965);
  nand n42970(x42970, x42969, x42967);
  nand n42972(x42972, x42961, x42967);
  nand n42973(x42973, x41769, x84951);
  nand n42975(x42975, x42974, x41770);
  nand n42976(x42976, x42975, x42973);
  nand n42977(x42977, x41788, x41797);
  nand n42978(x42978, x41787, x41796);
  nand n42979(x42979, x42978, x42977);
  nand n42981(x42981, x41806, x42980);
  nand n42982(x42982, x41805, x42979);
  nand n42983(x42983, x42982, x42981);
  nand n42985(x42985, x42977, x42981);
  nand n42986(x42986, x41815, x41824);
  nand n42987(x42987, x41814, x41823);
  nand n42988(x42988, x42987, x42986);
  nand n42990(x42990, x41833, x42989);
  nand n42991(x42991, x41832, x42988);
  nand n42992(x42992, x42991, x42990);
  nand n42994(x42994, x42986, x42990);
  nand n42995(x42995, x41780, x41789);
  nand n42998(x42998, x42997, x42996);
  nand n42999(x42999, x42998, x42995);
  nand n43001(x43001, x41798, x43000);
  nand n43003(x43003, x43002, x42999);
  nand n43004(x43004, x43003, x43001);
  nand n43005(x43005, x42995, x43001);
  nand n43006(x43006, x41807, x41816);
  nand n43009(x43009, x43008, x43007);
  nand n43010(x43010, x43009, x43006);
  nand n43012(x43012, x41825, x43011);
  nand n43014(x43014, x43013, x43010);
  nand n43015(x43015, x43014, x43012);
  nand n43017(x43017, x43006, x43012);
  nand n43018(x43018, x41834, x41842);
  nand n43021(x43021, x43020, x43019);
  nand n43022(x43022, x43021, x43018);
  nand n43023(x43023, x41858, x41867);
  nand n43024(x43024, x41857, x41866);
  nand n43025(x43025, x43024, x43023);
  nand n43027(x43027, x41876, x43026);
  nand n43028(x43028, x41875, x43025);
  nand n43029(x43029, x43028, x43027);
  nand n43031(x43031, x43023, x43027);
  nand n43032(x43032, x41885, x41894);
  nand n43033(x43033, x41884, x41893);
  nand n43034(x43034, x43033, x43032);
  nand n43036(x43036, x41903, x43035);
  nand n43037(x43037, x41902, x43034);
  nand n43038(x43038, x43037, x43036);
  nand n43040(x43040, x43032, x43036);
  nand n43041(x43041, x41912, x84952);
  nand n43042(x43042, x41911, x40611);
  nand n43043(x43043, x43042, x43041);
  nand n43044(x43044, x41850, x41859);
  nand n43047(x43047, x43046, x43045);
  nand n43048(x43048, x43047, x43044);
  nand n43050(x43050, x41868, x43049);
  nand n43052(x43052, x43051, x43048);
  nand n43053(x43053, x43052, x43050);
  nand n43055(x43055, x43044, x43050);
  nand n43056(x43056, x41877, x41886);
  nand n43059(x43059, x43058, x43057);
  nand n43060(x43060, x43059, x43056);
  nand n43062(x43062, x41895, x43061);
  nand n43064(x43064, x43063, x43060);
  nand n43065(x43065, x43064, x43062);
  nand n43067(x43067, x43056, x43062);
  nand n43068(x43068, x41904, x41913);
  nand n43071(x43071, x43070, x43069);
  nand n43072(x43072, x43071, x43068);
  nand n43073(x43073, x41929, x41938);
  nand n43074(x43074, x41928, x41937);
  nand n43075(x43075, x43074, x43073);
  nand n43077(x43077, x41947, x43076);
  nand n43078(x43078, x41946, x43075);
  nand n43079(x43079, x43078, x43077);
  nand n43081(x43081, x43073, x43077);
  nand n43082(x43082, x41956, x41965);
  nand n43083(x43083, x41955, x41964);
  nand n43084(x43084, x43083, x43082);
  nand n43086(x43086, x41974, x43085);
  nand n43087(x43087, x41973, x43084);
  nand n43088(x43088, x43087, x43086);
  nand n43090(x43090, x43082, x43086);
  nand n43091(x43091, x41983, x84953);
  nand n43092(x43092, x41982, x41987);
  nand n43093(x43093, x43092, x43091);
  nand n43094(x43094, x41921, x41930);
  nand n43097(x43097, x43096, x43095);
  nand n43098(x43098, x43097, x43094);
  nand n43100(x43100, x41939, x43099);
  nand n43102(x43102, x43101, x43098);
  nand n43103(x43103, x43102, x43100);
  nand n43105(x43105, x43094, x43100);
  nand n43106(x43106, x41948, x41957);
  nand n43109(x43109, x43108, x43107);
  nand n43110(x43110, x43109, x43106);
  nand n43112(x43112, x41966, x43111);
  nand n43114(x43114, x43113, x43110);
  nand n43115(x43115, x43114, x43112);
  nand n43117(x43117, x43106, x43112);
  nand n43118(x43118, x41975, x41984);
  nand n43121(x43121, x43120, x43119);
  nand n43122(x43122, x43121, x43118);
  nand n43124(x43124, x84954, x43123);
  nand n43125(x43125, x41985, x43122);
  nand n43126(x43126, x43125, x43124);
  nand n43128(x43128, x43118, x43124);
  nand n43129(x43129, x42003, x42012);
  nand n43130(x43130, x42002, x42011);
  nand n43131(x43131, x43130, x43129);
  nand n43133(x43133, x42021, x43132);
  nand n43134(x43134, x42020, x43131);
  nand n43135(x43135, x43134, x43133);
  nand n43137(x43137, x43129, x43133);
  nand n43138(x43138, x42030, x42039);
  nand n43139(x43139, x42029, x42038);
  nand n43140(x43140, x43139, x43138);
  nand n43142(x43142, x42048, x43141);
  nand n43143(x43143, x42047, x43140);
  nand n43144(x43144, x43143, x43142);
  nand n43146(x43146, x43138, x43142);
  nand n43147(x43147, x42057, x42066);
  nand n43148(x43148, x42056, x42065);
  nand n43149(x43149, x43148, x43147);
  nand n43150(x43150, x41995, x42004);
  nand n43153(x43153, x43152, x43151);
  nand n43154(x43154, x43153, x43150);
  nand n43156(x43156, x42013, x43155);
  nand n43158(x43158, x43157, x43154);
  nand n43159(x43159, x43158, x43156);
  nand n43161(x43161, x43150, x43156);
  nand n43162(x43162, x42022, x42031);
  nand n43165(x43165, x43164, x43163);
  nand n43166(x43166, x43165, x43162);
  nand n43168(x43168, x42040, x43167);
  nand n43170(x43170, x43169, x43166);
  nand n43171(x43171, x43170, x43168);
  nand n43173(x43173, x43162, x43168);
  nand n43174(x43174, x42049, x42058);
  nand n43177(x43177, x43176, x43175);
  nand n43178(x43178, x43177, x43174);
  nand n43180(x43180, x42067, x43179);
  nand n43182(x43182, x43181, x43178);
  nand n43183(x43183, x43182, x43180);
  nand n43185(x43185, x43174, x43180);
  nand n43186(x43186, x42083, x42092);
  nand n43187(x43187, x42082, x42091);
  nand n43188(x43188, x43187, x43186);
  nand n43190(x43190, x42101, x43189);
  nand n43191(x43191, x42100, x43188);
  nand n43192(x43192, x43191, x43190);
  nand n43194(x43194, x43186, x43190);
  nand n43195(x43195, x42110, x42119);
  nand n43196(x43196, x42109, x42118);
  nand n43197(x43197, x43196, x43195);
  nand n43199(x43199, x42128, x43198);
  nand n43200(x43200, x42127, x43197);
  nand n43201(x43201, x43200, x43199);
  nand n43203(x43203, x43195, x43199);
  nand n43204(x43204, x42137, x42146);
  nand n43205(x43205, x42136, x42145);
  nand n43206(x43206, x43205, x43204);
  nand n43208(x43208, x84955, x43207);
  nand n43209(x43209, x40772, x43206);
  nand n43210(x43210, x43209, x43208);
  nand n43212(x43212, x43204, x43208);
  nand n43213(x43213, x42075, x42084);
  nand n43216(x43216, x43215, x43214);
  nand n43217(x43217, x43216, x43213);
  nand n43219(x43219, x42093, x43218);
  nand n43221(x43221, x43220, x43217);
  nand n43222(x43222, x43221, x43219);
  nand n43224(x43224, x43213, x43219);
  nand n43225(x43225, x42102, x42111);
  nand n43228(x43228, x43227, x43226);
  nand n43229(x43229, x43228, x43225);
  nand n43231(x43231, x42120, x43230);
  nand n43233(x43233, x43232, x43229);
  nand n43234(x43234, x43233, x43231);
  nand n43236(x43236, x43225, x43231);
  nand n43237(x43237, x42129, x42138);
  nand n43240(x43240, x43239, x43238);
  nand n43241(x43241, x43240, x43237);
  nand n43243(x43243, x42147, x43242);
  nand n43245(x43245, x43244, x43241);
  nand n43246(x43246, x43245, x43243);
  nand n43248(x43248, x43237, x43243);
  nand n43249(x43249, x42163, x42172);
  nand n43250(x43250, x42162, x42171);
  nand n43251(x43251, x43250, x43249);
  nand n43253(x43253, x42181, x43252);
  nand n43254(x43254, x42180, x43251);
  nand n43255(x43255, x43254, x43253);
  nand n43257(x43257, x43249, x43253);
  nand n43258(x43258, x42190, x42199);
  nand n43259(x43259, x42189, x42198);
  nand n43260(x43260, x43259, x43258);
  nand n43262(x43262, x42208, x43261);
  nand n43263(x43263, x42207, x43260);
  nand n43264(x43264, x43263, x43262);
  nand n43266(x43266, x43258, x43262);
  nand n43267(x43267, x42217, x42226);
  nand n43268(x43268, x42216, x42225);
  nand n43269(x43269, x43268, x43267);
  nand n43271(x43271, x84956, x43270);
  nand n43272(x43272, x42230, x43269);
  nand n43273(x43273, x43272, x43271);
  nand n43275(x43275, x43267, x43271);
  nand n43276(x43276, x42155, x42164);
  nand n43279(x43279, x43278, x43277);
  nand n43280(x43280, x43279, x43276);
  nand n43282(x43282, x42173, x43281);
  nand n43284(x43284, x43283, x43280);
  nand n43285(x43285, x43284, x43282);
  nand n43287(x43287, x43276, x43282);
  nand n43288(x43288, x42182, x42191);
  nand n43291(x43291, x43290, x43289);
  nand n43292(x43292, x43291, x43288);
  nand n43294(x43294, x42200, x43293);
  nand n43296(x43296, x43295, x43292);
  nand n43297(x43297, x43296, x43294);
  nand n43299(x43299, x43288, x43294);
  nand n43300(x43300, x42209, x42218);
  nand n43303(x43303, x43302, x43301);
  nand n43304(x43304, x43303, x43300);
  nand n43306(x43306, x42227, x43305);
  nand n43308(x43308, x43307, x43304);
  nand n43309(x43309, x43308, x43306);
  nand n43311(x43311, x43300, x43306);
  nand n43312(x43312, x42238, x84999);
  nand n43313(x43313, x42237, x42228);
  nand n43314(x43314, x43313, x43312);
  nand n43316(x43316, x42247, x42256);
  nand n43317(x43317, x42246, x42255);
  nand n43318(x43318, x43317, x43316);
  nand n43320(x43320, x42265, x43319);
  nand n43321(x43321, x42264, x43318);
  nand n43322(x43322, x43321, x43320);
  nand n43324(x43324, x43316, x43320);
  nand n43325(x43325, x42274, x42283);
  nand n43326(x43326, x42273, x42282);
  nand n43327(x43327, x43326, x43325);
  nand n43329(x43329, x42292, x43328);
  nand n43330(x43330, x42291, x43327);
  nand n43331(x43331, x43330, x43329);
  nand n43333(x43333, x43325, x43329);
  nand n43334(x43334, x42301, x42310);
  nand n43335(x43335, x42300, x42309);
  nand n43336(x43336, x43335, x43334);
  nand n43338(x43338, x42319, x43337);
  nand n43339(x43339, x42318, x43336);
  nand n43340(x43340, x43339, x43338);
  nand n43342(x43342, x43334, x43338);
  nand n43343(x43343, x42239, x42248);
  nand n43346(x43346, x43345, x43344);
  nand n43347(x43347, x43346, x43343);
  nand n43349(x43349, x42257, x43348);
  nand n43351(x43351, x43350, x43347);
  nand n43352(x43352, x43351, x43349);
  nand n43354(x43354, x43343, x43349);
  nand n43355(x43355, x42266, x42275);
  nand n43358(x43358, x43357, x43356);
  nand n43359(x43359, x43358, x43355);
  nand n43361(x43361, x42284, x43360);
  nand n43363(x43363, x43362, x43359);
  nand n43364(x43364, x43363, x43361);
  nand n43366(x43366, x43355, x43361);
  nand n43367(x43367, x42293, x42302);
  nand n43370(x43370, x43369, x43368);
  nand n43371(x43371, x43370, x43367);
  nand n43373(x43373, x42311, x43372);
  nand n43375(x43375, x43374, x43371);
  nand n43376(x43376, x43375, x43373);
  nand n43378(x43378, x43367, x43373);
  nand n43380(x43380, x42328, x42320);
  nand n43381(x43381, x42327, x43379);
  nand n43382(x43382, x43381, x43380);
  nand n43384(x43384, x42337, x42346);
  nand n43385(x43385, x42336, x42345);
  nand n43386(x43386, x43385, x43384);
  nand n43388(x43388, x42355, x43387);
  nand n43389(x43389, x42354, x43386);
  nand n43390(x43390, x43389, x43388);
  nand n43392(x43392, x43384, x43388);
  nand n43393(x43393, x42364, x42373);
  nand n43394(x43394, x42363, x42372);
  nand n43395(x43395, x43394, x43393);
  nand n43397(x43397, x42382, x43396);
  nand n43398(x43398, x42381, x43395);
  nand n43399(x43399, x43398, x43397);
  nand n43401(x43401, x43393, x43397);
  nand n43402(x43402, x42391, x42400);
  nand n43403(x43403, x42390, x42399);
  nand n43404(x43404, x43403, x43402);
  nand n43406(x43406, x42409, x43405);
  nand n43407(x43407, x42408, x43404);
  nand n43408(x43408, x43407, x43406);
  nand n43410(x43410, x43402, x43406);
  nand n43411(x43411, x42329, x42338);
  nand n43414(x43414, x43413, x43412);
  nand n43415(x43415, x43414, x43411);
  nand n43417(x43417, x42347, x43416);
  nand n43419(x43419, x43418, x43415);
  nand n43420(x43420, x43419, x43417);
  nand n43422(x43422, x42356, x42365);
  nand n43425(x43425, x43424, x43423);
  nand n43426(x43426, x43425, x43422);
  nand n43428(x43428, x42374, x43427);
  nand n43430(x43430, x43429, x43426);
  nand n43431(x43431, x43430, x43428);
  nand n43433(x43433, x42383, x42392);
  nand n43436(x43436, x43435, x43434);
  nand n43437(x43437, x43436, x43433);
  nand n43439(x43439, x42401, x43438);
  nand n43441(x43441, x43440, x43437);
  nand n43442(x43442, x43441, x43439);
  nand n43445(x43445, x42418, x42410);
  nand n43446(x43446, x42417, x43444);
  nand n43447(x43447, x43446, x43445);
  nand n43449(x43449, x42426, x42434);
  nand n43450(x43450, x42425, x42433);
  nand n43451(x43451, x43450, x43449);
  nand n43453(x43453, x42442, x43452);
  nand n43454(x43454, x42441, x43451);
  nand n43455(x43455, x43454, x43453);
  nand n43457(x43457, x42450, x42458);
  nand n43458(x43458, x42449, x42457);
  nand n43459(x43459, x43458, x43457);
  nand n43461(x43461, x42466, x43460);
  nand n43462(x43462, x42465, x43459);
  nand n43463(x43463, x43462, x43461);
  nand n43465(x43465, x42474, x42482);
  nand n43466(x43466, x42473, x42481);
  nand n43467(x43467, x43466, x43465);
  nand n43469(x43469, x42490, x43468);
  nand n43470(x43470, x42489, x43467);
  nand n43471(x43471, x43470, x43469);
  nand n43473(x43473, x84958, x85004);
  nand n43474(x43474, x39988, x41033);
  nand n43475(x43475, x43474, x43473);
  nand n43477(x43477, x84959, x85005);
  nand n43478(x43478, x41045, x41041);
  nand n43479(x43479, x43478, x43477);
  nand n43481(x43481, x84960, x85006);
  nand n43482(x43482, x41060, x41052);
  nand n43483(x43483, x43482, x43481);
  nand n43485(x43485, x84961, x85008);
  nand n43486(x43486, x42508, x41068);
  nand n43487(x43487, x43486, x43485);
  nand n43489(x43489, x84962, x85012);
  nand n43490(x43490, x42516, x41085);
  nand n43491(x43491, x43490, x43489);
  nand n43493(x43493, x84963, x85016);
  nand n43494(x43494, x42529, x41105);
  nand n43495(x43495, x43494, x43493);
  nand n43498(x43498, x42548, x85019);
  nand n43499(x43499, x42547, x41131);
  nand n43500(x43500, x43499, x43498);
  nand n43504(x43504, x42568, x85021);
  nand n43505(x43505, x42567, x41157);
  nand n43506(x43506, x43505, x43504);
  nand n43510(x43510, x84964, x85022);
  nand n43511(x43511, x41177, x42579);
  nand n43512(x43512, x43511, x43510);
  nand n43514(x43514, x42588, x85023);
  nand n43515(x43515, x42587, x41186);
  nand n43516(x43516, x43515, x43514);
  nand n43520(x43520, x41214, x85024);
  nand n43521(x43521, x42601, x42599);
  nand n43522(x43522, x43521, x43520);
  nand n43524(x43524, x42609, x85025);
  nand n43525(x43525, x42608, x41221);
  nand n43526(x43526, x43525, x43524);
  nand n43530(x43530, x41249, x85027);
  nand n43531(x43531, x42622, x42620);
  nand n43532(x43532, x43531, x43530);
  nand n43534(x43534, x42630, x85028);
  nand n43535(x43535, x42629, x41256);
  nand n43536(x43536, x43535, x43534);
  nand n43540(x43540, x84965, x85030);
  nand n43541(x43541, x42646, x42641);
  nand n43542(x43542, x43541, x43540);
  nand n43544(x43544, x42654, x85031);
  nand n43545(x43545, x42653, x41294);
  nand n43546(x43546, x43545, x43544);
  nand n43548(x43548, x42642, x84966);
  nand n43550(x43550, x43549, x42643);
  nand n43551(x43551, x43550, x43548);
  nand n43553(x43553, x84967, x85034);
  nand n43554(x43554, x42671, x42665);
  nand n43555(x43555, x43554, x43553);
  nand n43557(x43557, x42679, x85036);
  nand n43558(x43558, x42678, x41337);
  nand n43559(x43559, x43558, x43557);
  nand n43561(x43561, x42666, x84968);
  nand n43563(x43563, x43562, x42667);
  nand n43564(x43564, x43563, x43561);
  nand n43566(x43566, x84969, x42680);
  nand n43567(x43567, x42681, x43565);
  nand n43568(x43568, x43567, x43566);
  nand n43570(x43570, x84970, x85041);
  nand n43571(x43571, x42699, x42693);
  nand n43572(x43572, x43571, x43570);
  nand n43574(x43574, x42707, x85043);
  nand n43575(x43575, x42706, x41381);
  nand n43576(x43576, x43575, x43574);
  nand n43578(x43578, x42694, x84971);
  nand n43580(x43580, x43579, x42695);
  nand n43581(x43581, x43580, x43578);
  nand n43583(x43583, x84972, x42708);
  nand n43584(x43584, x42709, x43582);
  nand n43585(x43585, x43584, x43583);
  nand n43587(x43587, x42732, x85048);
  nand n43588(x43588, x42731, x42721);
  nand n43589(x43589, x43588, x43587);
  nand n43591(x43591, x42741, x85050);
  nand n43592(x43592, x42740, x41428);
  nand n43593(x43593, x43592, x43591);
  nand n43595(x43595, x42722, x42733);
  nand n43598(x43598, x43597, x43596);
  nand n43599(x43599, x43598, x43595);
  nand n43601(x43601, x84973, x42742);
  nand n43602(x43602, x42743, x43600);
  nand n43603(x43603, x43602, x43601);
  nand n43605(x43605, x42767, x85055);
  nand n43606(x43606, x42766, x42755);
  nand n43607(x43607, x43606, x43605);
  nand n43609(x43609, x42776, x85057);
  nand n43610(x43610, x42775, x41481);
  nand n43611(x43611, x43610, x43609);
  nand n43613(x43613, x42756, x42768);
  nand n43616(x43616, x43615, x43614);
  nand n43617(x43617, x43616, x43613);
  nand n43619(x43619, x42785, x42777);
  nand n43621(x43621, x43620, x43618);
  nand n43622(x43622, x43621, x43619);
  nand n43624(x43624, x42807, x85062);
  nand n43625(x43625, x42806, x42795);
  nand n43626(x43626, x43625, x43624);
  nand n43628(x43628, x42816, x85064);
  nand n43629(x43629, x42815, x41534);
  nand n43630(x43630, x43629, x43628);
  nand n43632(x43632, x42796, x42808);
  nand n43635(x43635, x43634, x43633);
  nand n43636(x43636, x43635, x43632);
  nand n43638(x43638, x42825, x42817);
  nand n43640(x43640, x43639, x43637);
  nand n43641(x43641, x43640, x43638);
  nand n43643(x43643, x42847, x85069);
  nand n43644(x43644, x42846, x42835);
  nand n43645(x43645, x43644, x43643);
  nand n43647(x43647, x84974, x84975);
  nand n43648(x43648, x41581, x41590);
  nand n43649(x43649, x43648, x43647);
  nand n43651(x43651, x42856, x43650);
  nand n43652(x43652, x42855, x43649);
  nand n43653(x43653, x43652, x43651);
  nand n43655(x43655, x43647, x43651);
  nand n43656(x43656, x42836, x42848);
  nand n43659(x43659, x43658, x43657);
  nand n43660(x43660, x43659, x43656);
  nand n43662(x43662, x42865, x42857);
  nand n43664(x43664, x43663, x43661);
  nand n43665(x43665, x43664, x43662);
  nand n43667(x43667, x42887, x85075);
  nand n43668(x43668, x42886, x42875);
  nand n43669(x43669, x43668, x43667);
  nand n43671(x43671, x41645, x84976);
  nand n43672(x43672, x42889, x41652);
  nand n43673(x43673, x43672, x43671);
  nand n43675(x43675, x42897, x43674);
  nand n43676(x43676, x42896, x43673);
  nand n43677(x43677, x43676, x43675);
  nand n43679(x43679, x43671, x43675);
  nand n43680(x43680, x42906, x84977);
  nand n43681(x43681, x42905, x40468);
  nand n43682(x43682, x43681, x43680);
  nand n43683(x43683, x42876, x42888);
  nand n43686(x43686, x43685, x43684);
  nand n43687(x43687, x43686, x43683);
  nand n43689(x43689, x42907, x42898);
  nand n43691(x43691, x43690, x43688);
  nand n43692(x43692, x43691, x43689);
  nand n43694(x43694, x42929, x85082);
  nand n43695(x43695, x42928, x42917);
  nand n43696(x43696, x43695, x43694);
  nand n43698(x43698, x41707, x84978);
  nand n43699(x43699, x42931, x41714);
  nand n43700(x43700, x43699, x43698);
  nand n43702(x43702, x42939, x43701);
  nand n43703(x43703, x42938, x43700);
  nand n43704(x43704, x43703, x43702);
  nand n43706(x43706, x43698, x43702);
  nand n43707(x43707, x42948, x84979);
  nand n43708(x43708, x42947, x41772);
  nand n43709(x43709, x43708, x43707);
  nand n43710(x43710, x42918, x42930);
  nand n43713(x43713, x43712, x43711);
  nand n43714(x43714, x43713, x43710);
  nand n43716(x43716, x42949, x42940);
  nand n43718(x43718, x43717, x43715);
  nand n43719(x43719, x43718, x43716);
  nand n43721(x43721, x42971, x85089);
  nand n43722(x43722, x42970, x42959);
  nand n43723(x43723, x43722, x43721);
  nand n43725(x43725, x84980, x84982);
  nand n43726(x43726, x42976, x41779);
  nand n43727(x43727, x43726, x43725);
  nand n43729(x43729, x42984, x43728);
  nand n43730(x43730, x42983, x43727);
  nand n43731(x43731, x43730, x43729);
  nand n43733(x43733, x43725, x43729);
  nand n43734(x43734, x42993, x84983);
  nand n43735(x43735, x42992, x41841);
  nand n43736(x43736, x43735, x43734);
  nand n43737(x43737, x42960, x42972);
  nand n43740(x43740, x43739, x43738);
  nand n43741(x43741, x43740, x43737);
  nand n43743(x43743, x84981, x43742);
  nand n43744(x43744, x42973, x43741);
  nand n43745(x43745, x43744, x43743);
  nand n43747(x43747, x43737, x43743);
  nand n43749(x43749, x42994, x42985);
  nand n43751(x43751, x43750, x43748);
  nand n43752(x43752, x43751, x43749);
  nand n43754(x43754, x43016, x85094);
  nand n43755(x43755, x43015, x43004);
  nand n43756(x43756, x43755, x43754);
  nand n43758(x43758, x84984, x84986);
  nand n43759(x43759, x43022, x41849);
  nand n43760(x43760, x43759, x43758);
  nand n43762(x43762, x43030, x43761);
  nand n43763(x43763, x43029, x43760);
  nand n43764(x43764, x43763, x43762);
  nand n43766(x43766, x43758, x43762);
  nand n43767(x43767, x43039, x84987);
  nand n43768(x43768, x43038, x43043);
  nand n43769(x43769, x43768, x43767);
  nand n43770(x43770, x43005, x43017);
  nand n43773(x43773, x43772, x43771);
  nand n43774(x43774, x43773, x43770);
  nand n43776(x43776, x84985, x43775);
  nand n43777(x43777, x43018, x43774);
  nand n43778(x43778, x43777, x43776);
  nand n43780(x43780, x43770, x43776);
  nand n43782(x43782, x43040, x43031);
  nand n43784(x43784, x43783, x43781);
  nand n43785(x43785, x43784, x43782);
  nand n43787(x43787, x84988, x43054);
  nand n43788(x43788, x43041, x43053);
  nand n43789(x43789, x43788, x43787);
  nand n43791(x43791, x43066, x43790);
  nand n43792(x43792, x43065, x43789);
  nand n43793(x43793, x43792, x43791);
  nand n43795(x43795, x43787, x43791);
  nand n43796(x43796, x84989, x84991);
  nand n43797(x43797, x43072, x41920);
  nand n43798(x43798, x43797, x43796);
  nand n43800(x43800, x43080, x43799);
  nand n43801(x43801, x43079, x43798);
  nand n43802(x43802, x43801, x43800);
  nand n43804(x43804, x43796, x43800);
  nand n43805(x43805, x43089, x84992);
  nand n43806(x43806, x43088, x43093);
  nand n43807(x43807, x43806, x43805);
  nand n43808(x43808, x43055, x43067);
  nand n43811(x43811, x43810, x43809);
  nand n43812(x43812, x43811, x43808);
  nand n43814(x43814, x84990, x43813);
  nand n43815(x43815, x43068, x43812);
  nand n43816(x43816, x43815, x43814);
  nand n43818(x43818, x43808, x43814);
  nand n43820(x43820, x43090, x43081);
  nand n43822(x43822, x43821, x43819);
  nand n43823(x43823, x43822, x43820);
  nand n43825(x43825, x84993, x43104);
  nand n43826(x43826, x43091, x43103);
  nand n43827(x43827, x43826, x43825);
  nand n43829(x43829, x43116, x43828);
  nand n43830(x43830, x43115, x43827);
  nand n43831(x43831, x43830, x43829);
  nand n43833(x43833, x43825, x43829);
  nand n43834(x43834, x43127, x84994);
  nand n43835(x43835, x43126, x41994);
  nand n43836(x43836, x43835, x43834);
  nand n43838(x43838, x43136, x43837);
  nand n43839(x43839, x43135, x43836);
  nand n43840(x43840, x43839, x43838);
  nand n43842(x43842, x43834, x43838);
  nand n43843(x43843, x43145, x84995);
  nand n43844(x43844, x43144, x43149);
  nand n43845(x43845, x43844, x43843);
  nand n43846(x43846, x43105, x43117);
  nand n43849(x43849, x43848, x43847);
  nand n43850(x43850, x43849, x43846);
  nand n43852(x43852, x43128, x43851);
  nand n43854(x43854, x43853, x43850);
  nand n43855(x43855, x43854, x43852);
  nand n43857(x43857, x43846, x43852);
  nand n43859(x43859, x43146, x43137);
  nand n43861(x43861, x43860, x43858);
  nand n43862(x43862, x43861, x43859);
  nand n43864(x43864, x84996, x43160);
  nand n43865(x43865, x43147, x43159);
  nand n43866(x43866, x43865, x43864);
  nand n43868(x43868, x43172, x43867);
  nand n43869(x43869, x43171, x43866);
  nand n43870(x43870, x43869, x43868);
  nand n43872(x43872, x43864, x43868);
  nand n43873(x43873, x43184, x84997);
  nand n43874(x43874, x43183, x42074);
  nand n43875(x43875, x43874, x43873);
  nand n43877(x43877, x43193, x43876);
  nand n43878(x43878, x43192, x43875);
  nand n43879(x43879, x43878, x43877);
  nand n43881(x43881, x43873, x43877);
  nand n43882(x43882, x43202, x43211);
  nand n43883(x43883, x43201, x43210);
  nand n43884(x43884, x43883, x43882);
  nand n43885(x43885, x43161, x43173);
  nand n43888(x43888, x43887, x43886);
  nand n43889(x43889, x43888, x43885);
  nand n43891(x43891, x43185, x43890);
  nand n43893(x43893, x43892, x43889);
  nand n43894(x43894, x43893, x43891);
  nand n43896(x43896, x43885, x43891);
  nand n43898(x43898, x43203, x43194);
  nand n43900(x43900, x43899, x43897);
  nand n43901(x43901, x43900, x43898);
  nand n43903(x43903, x43212, x43223);
  nand n43905(x43905, x43904, x43222);
  nand n43906(x43906, x43905, x43903);
  nand n43908(x43908, x43235, x43907);
  nand n43909(x43909, x43234, x43906);
  nand n43910(x43910, x43909, x43908);
  nand n43912(x43912, x43903, x43908);
  nand n43913(x43913, x43247, x84998);
  nand n43914(x43914, x43246, x42154);
  nand n43915(x43915, x43914, x43913);
  nand n43917(x43917, x43256, x43916);
  nand n43918(x43918, x43255, x43915);
  nand n43919(x43919, x43918, x43917);
  nand n43921(x43921, x43913, x43917);
  nand n43922(x43922, x43265, x43274);
  nand n43923(x43923, x43264, x43273);
  nand n43924(x43924, x43923, x43922);
  nand n43925(x43925, x43224, x43236);
  nand n43928(x43928, x43927, x43926);
  nand n43929(x43929, x43928, x43925);
  nand n43931(x43931, x43248, x43930);
  nand n43933(x43933, x43932, x43929);
  nand n43934(x43934, x43933, x43931);
  nand n43936(x43936, x43925, x43931);
  nand n43938(x43938, x43266, x43257);
  nand n43940(x43940, x43939, x43937);
  nand n43941(x43941, x43940, x43938);
  nand n43943(x43943, x43275, x43286);
  nand n43945(x43945, x43944, x43285);
  nand n43946(x43946, x43945, x43943);
  nand n43948(x43948, x43298, x43947);
  nand n43949(x43949, x43297, x43946);
  nand n43950(x43950, x43949, x43948);
  nand n43952(x43952, x43943, x43948);
  nand n43953(x43953, x43310, x43315);
  nand n43954(x43954, x43309, x43314);
  nand n43955(x43955, x43954, x43953);
  nand n43957(x43957, x43323, x43956);
  nand n43958(x43958, x43322, x43955);
  nand n43959(x43959, x43958, x43957);
  nand n43961(x43961, x43953, x43957);
  nand n43962(x43962, x43332, x43341);
  nand n43963(x43963, x43331, x43340);
  nand n43964(x43964, x43963, x43962);
  nand n43965(x43965, x43287, x43299);
  nand n43968(x43968, x43967, x43966);
  nand n43969(x43969, x43968, x43965);
  nand n43971(x43971, x43311, x43970);
  nand n43973(x43973, x43972, x43969);
  nand n43974(x43974, x43973, x43971);
  nand n43976(x43976, x43965, x43971);
  nand n43977(x43977, x85000, x43324);
  nand n43979(x43979, x43312, x43978);
  nand n43980(x43980, x43979, x43977);
  nand n43982(x43982, x43333, x43981);
  nand n43984(x43984, x43983, x43980);
  nand n43985(x43985, x43984, x43982);
  nand n43987(x43987, x43977, x43982);
  nand n43988(x43988, x43342, x43353);
  nand n43990(x43990, x43989, x43352);
  nand n43991(x43991, x43990, x43988);
  nand n43993(x43993, x43365, x43992);
  nand n43994(x43994, x43364, x43991);
  nand n43995(x43995, x43994, x43993);
  nand n43997(x43997, x43988, x43993);
  nand n43998(x43998, x43377, x43383);
  nand n43999(x43999, x43376, x43382);
  nand n44000(x44000, x43999, x43998);
  nand n44002(x44002, x43391, x44001);
  nand n44003(x44003, x43390, x44000);
  nand n44004(x44004, x44003, x44002);
  nand n44006(x44006, x43998, x44002);
  nand n44007(x44007, x43400, x43409);
  nand n44008(x44008, x43399, x43408);
  nand n44009(x44009, x44008, x44007);
  nand n44011(x44011, x84957, x44010);
  nand n44012(x44012, x40951, x44009);
  nand n44013(x44013, x44012, x44011);
  nand n44015(x44015, x44007, x44011);
  nand n44016(x44016, x43354, x43366);
  nand n44019(x44019, x44018, x44017);
  nand n44020(x44020, x44019, x44016);
  nand n44022(x44022, x43378, x44021);
  nand n44024(x44024, x44023, x44020);
  nand n44025(x44025, x44024, x44022);
  nand n44027(x44027, x85001, x43392);
  nand n44029(x44029, x43380, x44028);
  nand n44030(x44030, x44029, x44027);
  nand n44032(x44032, x43401, x44031);
  nand n44034(x44034, x44033, x44030);
  nand n44035(x44035, x44034, x44032);
  nand n44037(x44037, x43410, x43421);
  nand n44039(x44039, x44038, x43420);
  nand n44040(x44040, x44039, x44037);
  nand n44042(x44042, x43432, x44041);
  nand n44043(x44043, x43431, x44040);
  nand n44044(x44044, x44043, x44042);
  nand n44046(x44046, x43443, x43448);
  nand n44047(x44047, x43442, x43447);
  nand n44048(x44048, x44047, x44046);
  nand n44050(x44050, x43456, x44049);
  nand n44051(x44051, x43455, x44048);
  nand n44052(x44052, x44051, x44050);
  nand n44054(x44054, x43464, x43472);
  nand n44055(x44055, x43463, x43471);
  nand n44056(x44056, x44055, x44054);
  nand n44058(x44058, x42494, x44057);
  nand n44059(x44059, x42493, x44056);
  nand n44060(x44060, x44059, x44058);
  nand n44062(x44062, x85002, x85003);
  nand n44063(x44063, x41016, x41025);
  nand n44064(x44064, x44063, x44062);
  nand n44065(x44065, x43476, x41026);
  nand n44066(x44066, x43475, x42495);
  nand n44067(x44067, x44066, x44065);
  nand n44068(x44068, x43480, x41034);
  nand n44069(x44069, x43479, x42496);
  nand n44070(x44070, x44069, x44068);
  nand n44072(x44072, x43484, x85113);
  nand n44073(x44073, x43483, x42500);
  nand n44074(x44074, x44073, x44072);
  nand n44076(x44076, x85007, x85114);
  nand n44077(x44077, x42497, x43481);
  nand n44078(x44078, x44077, x44076);
  nand n44079(x44079, x43488, x85115);
  nand n44080(x44080, x43487, x42505);
  nand n44081(x44081, x44080, x44079);
  nand n44083(x44083, x85009, x85117);
  nand n44084(x44084, x42501, x43485);
  nand n44085(x44085, x44084, x44083);
  nand n44086(x44086, x85010, x85011);
  nand n44087(x44087, x42506, x42513);
  nand n44088(x44088, x44087, x44086);
  nand n44090(x44090, x43492, x44089);
  nand n44091(x44091, x43491, x44088);
  nand n44092(x44092, x44091, x44090);
  nand n44094(x44094, x44086, x44090);
  nand n44095(x44095, x85013, x85118);
  nand n44096(x44096, x42509, x43489);
  nand n44097(x44097, x44096, x44095);
  nand n44098(x44098, x85014, x85015);
  nand n44099(x44099, x42514, x42525);
  nand n44100(x44100, x44099, x44098);
  nand n44102(x44102, x43496, x44101);
  nand n44103(x44103, x43495, x44100);
  nand n44104(x44104, x44103, x44102);
  nand n44106(x44106, x44098, x44102);
  nand n44107(x44107, x42526, x85119);
  nand n44108(x44108, x43497, x43493);
  nand n44109(x44109, x44108, x44107);
  nand n44110(x44110, x85017, x85018);
  nand n44111(x44111, x42527, x42539);
  nand n44112(x44112, x44111, x44110);
  nand n44114(x44114, x43501, x44113);
  nand n44115(x44115, x43500, x44112);
  nand n44116(x44116, x44115, x44114);
  nand n44118(x44118, x44110, x44114);
  nand n44119(x44119, x42540, x85120);
  nand n44120(x44120, x43502, x43498);
  nand n44121(x44121, x44120, x44119);
  nand n44122(x44122, x42549, x85020);
  nand n44123(x44123, x43503, x42559);
  nand n44124(x44124, x44123, x44122);
  nand n44126(x44126, x43507, x44125);
  nand n44127(x44127, x43506, x44124);
  nand n44128(x44128, x44127, x44126);
  nand n44130(x44130, x44122, x44126);
  nand n44131(x44131, x42560, x85121);
  nand n44132(x44132, x43508, x43504);
  nand n44133(x44133, x44132, x44131);
  nand n44134(x44134, x42569, x43513);
  nand n44135(x44135, x43509, x43512);
  nand n44136(x44136, x44135, x44134);
  nand n44138(x44138, x43517, x44137);
  nand n44139(x44139, x43516, x44136);
  nand n44140(x44140, x44139, x44138);
  nand n44142(x44142, x44134, x44138);
  nand n44143(x44143, x42580, x85123);
  nand n44144(x44144, x43518, x43514);
  nand n44145(x44145, x44144, x44143);
  nand n44147(x44147, x42589, x43523);
  nand n44148(x44148, x43519, x43522);
  nand n44149(x44149, x44148, x44147);
  nand n44151(x44151, x43527, x44150);
  nand n44152(x44152, x43526, x44149);
  nand n44153(x44153, x44152, x44151);
  nand n44155(x44155, x44147, x44151);
  nand n44156(x44156, x42600, x85125);
  nand n44157(x44157, x43528, x43524);
  nand n44158(x44158, x44157, x44156);
  nand n44160(x44160, x42610, x43533);
  nand n44161(x44161, x43529, x43532);
  nand n44162(x44162, x44161, x44160);
  nand n44164(x44164, x43537, x44163);
  nand n44165(x44165, x43536, x44162);
  nand n44166(x44166, x44165, x44164);
  nand n44168(x44168, x44160, x44164);
  nand n44169(x44169, x42621, x85127);
  nand n44170(x44170, x43538, x43534);
  nand n44171(x44171, x44170, x44169);
  nand n44173(x44173, x42631, x43543);
  nand n44174(x44174, x43539, x43542);
  nand n44175(x44175, x44174, x44173);
  nand n44177(x44177, x43547, x44176);
  nand n44178(x44178, x43546, x44175);
  nand n44179(x44179, x44178, x44177);
  nand n44181(x44181, x44173, x44177);
  nand n44182(x44182, x85033, x85129);
  nand n44183(x44183, x43551, x43544);
  nand n44184(x44184, x44183, x44182);
  nand n44186(x44186, x42655, x43556);
  nand n44187(x44187, x43552, x43555);
  nand n44188(x44188, x44187, x44186);
  nand n44190(x44190, x43560, x44189);
  nand n44191(x44191, x43559, x44188);
  nand n44192(x44192, x44191, x44190);
  nand n44194(x44194, x44186, x44190);
  nand n44195(x44195, x85035, x85130);
  nand n44196(x44196, x43553, x43548);
  nand n44197(x44197, x44196, x44195);
  nand n44199(x44199, x85038, x85132);
  nand n44200(x44200, x43564, x43557);
  nand n44201(x44201, x44200, x44199);
  nand n44203(x44203, x43569, x43573);
  nand n44204(x44204, x43568, x43572);
  nand n44205(x44205, x44204, x44203);
  nand n44207(x44207, x43577, x44206);
  nand n44208(x44208, x43576, x44205);
  nand n44209(x44209, x44208, x44207);
  nand n44211(x44211, x44203, x44207);
  nand n44212(x44212, x85039, x85040);
  nand n44213(x44213, x43561, x43566);
  nand n44214(x44214, x44213, x44212);
  nand n44216(x44216, x85042, x44215);
  nand n44217(x44217, x43570, x44214);
  nand n44218(x44218, x44217, x44216);
  nand n44220(x44220, x44212, x44216);
  nand n44221(x44221, x85045, x85134);
  nand n44222(x44222, x43581, x43574);
  nand n44223(x44223, x44222, x44221);
  nand n44225(x44225, x43586, x43590);
  nand n44226(x44226, x43585, x43589);
  nand n44227(x44227, x44226, x44225);
  nand n44229(x44229, x43594, x44228);
  nand n44230(x44230, x43593, x44227);
  nand n44231(x44231, x44230, x44229);
  nand n44233(x44233, x44225, x44229);
  nand n44234(x44234, x85046, x85047);
  nand n44235(x44235, x43578, x43583);
  nand n44236(x44236, x44235, x44234);
  nand n44238(x44238, x85049, x44237);
  nand n44239(x44239, x43587, x44236);
  nand n44240(x44240, x44239, x44238);
  nand n44242(x44242, x44234, x44238);
  nand n44243(x44243, x85052, x85136);
  nand n44244(x44244, x43599, x43591);
  nand n44245(x44245, x44244, x44243);
  nand n44247(x44247, x43604, x43608);
  nand n44248(x44248, x43603, x43607);
  nand n44249(x44249, x44248, x44247);
  nand n44251(x44251, x43612, x44250);
  nand n44252(x44252, x43611, x44249);
  nand n44253(x44253, x44252, x44251);
  nand n44255(x44255, x44247, x44251);
  nand n44256(x44256, x85053, x85054);
  nand n44257(x44257, x43595, x43601);
  nand n44258(x44258, x44257, x44256);
  nand n44260(x44260, x85056, x44259);
  nand n44261(x44261, x43605, x44258);
  nand n44262(x44262, x44261, x44260);
  nand n44264(x44264, x44256, x44260);
  nand n44265(x44265, x85059, x85138);
  nand n44266(x44266, x43617, x43609);
  nand n44267(x44267, x44266, x44265);
  nand n44269(x44269, x43623, x43627);
  nand n44270(x44270, x43622, x43626);
  nand n44271(x44271, x44270, x44269);
  nand n44273(x44273, x43631, x44272);
  nand n44274(x44274, x43630, x44271);
  nand n44275(x44275, x44274, x44273);
  nand n44277(x44277, x44269, x44273);
  nand n44278(x44278, x85060, x85061);
  nand n44279(x44279, x43613, x43619);
  nand n44280(x44280, x44279, x44278);
  nand n44282(x44282, x85063, x44281);
  nand n44283(x44283, x43624, x44280);
  nand n44284(x44284, x44283, x44282);
  nand n44286(x44286, x44278, x44282);
  nand n44287(x44287, x85066, x85140);
  nand n44288(x44288, x43636, x43628);
  nand n44289(x44289, x44288, x44287);
  nand n44291(x44291, x43642, x43646);
  nand n44292(x44292, x43641, x43645);
  nand n44293(x44293, x44292, x44291);
  nand n44295(x44295, x43654, x44294);
  nand n44296(x44296, x43653, x44293);
  nand n44297(x44297, x44296, x44295);
  nand n44299(x44299, x44291, x44295);
  nand n44300(x44300, x85067, x85068);
  nand n44301(x44301, x43632, x43638);
  nand n44302(x44302, x44301, x44300);
  nand n44304(x44304, x85070, x44303);
  nand n44305(x44305, x43643, x44302);
  nand n44306(x44306, x44305, x44304);
  nand n44308(x44308, x44300, x44304);
  nand n44310(x44310, x85072, x43655);
  nand n44311(x44311, x43660, x44309);
  nand n44312(x44312, x44311, x44310);
  nand n44314(x44314, x43666, x43670);
  nand n44315(x44315, x43665, x43669);
  nand n44316(x44316, x44315, x44314);
  nand n44318(x44318, x43678, x44317);
  nand n44319(x44319, x43677, x44316);
  nand n44320(x44320, x44319, x44318);
  nand n44322(x44322, x44314, x44318);
  nand n44323(x44323, x85073, x85074);
  nand n44324(x44324, x43656, x43662);
  nand n44325(x44325, x44324, x44323);
  nand n44327(x44327, x85076, x44326);
  nand n44328(x44328, x43667, x44325);
  nand n44329(x44329, x44328, x44327);
  nand n44331(x44331, x44323, x44327);
  nand n44332(x44332, x43679, x85078);
  nand n44334(x44334, x44333, x43680);
  nand n44335(x44335, x44334, x44332);
  nand n44337(x44337, x85079, x44336);
  nand n44338(x44338, x43687, x44335);
  nand n44339(x44339, x44338, x44337);
  nand n44341(x44341, x44332, x44337);
  nand n44342(x44342, x43693, x43697);
  nand n44343(x44343, x43692, x43696);
  nand n44344(x44344, x44343, x44342);
  nand n44346(x44346, x43705, x44345);
  nand n44347(x44347, x43704, x44344);
  nand n44348(x44348, x44347, x44346);
  nand n44350(x44350, x44342, x44346);
  nand n44351(x44351, x85080, x85081);
  nand n44352(x44352, x43683, x43689);
  nand n44353(x44353, x44352, x44351);
  nand n44355(x44355, x85083, x44354);
  nand n44356(x44356, x43694, x44353);
  nand n44357(x44357, x44356, x44355);
  nand n44359(x44359, x44351, x44355);
  nand n44360(x44360, x43706, x85085);
  nand n44362(x44362, x44361, x43707);
  nand n44363(x44363, x44362, x44360);
  nand n44365(x44365, x85086, x44364);
  nand n44366(x44366, x43714, x44363);
  nand n44367(x44367, x44366, x44365);
  nand n44369(x44369, x44360, x44365);
  nand n44370(x44370, x43720, x43724);
  nand n44371(x44371, x43719, x43723);
  nand n44372(x44372, x44371, x44370);
  nand n44374(x44374, x43732, x44373);
  nand n44375(x44375, x43731, x44372);
  nand n44376(x44376, x44375, x44374);
  nand n44378(x44378, x44370, x44374);
  nand n44379(x44379, x85087, x85088);
  nand n44380(x44380, x43710, x43716);
  nand n44381(x44381, x44380, x44379);
  nand n44383(x44383, x85090, x44382);
  nand n44384(x44384, x43721, x44381);
  nand n44385(x44385, x44384, x44383);
  nand n44387(x44387, x44379, x44383);
  nand n44388(x44388, x43733, x85092);
  nand n44390(x44390, x44389, x43734);
  nand n44391(x44391, x44390, x44388);
  nand n44393(x44393, x43746, x44392);
  nand n44394(x44394, x43745, x44391);
  nand n44395(x44395, x44394, x44393);
  nand n44397(x44397, x44388, x44393);
  nand n44398(x44398, x43753, x43757);
  nand n44399(x44399, x43752, x43756);
  nand n44400(x44400, x44399, x44398);
  nand n44402(x44402, x43765, x44401);
  nand n44403(x44403, x43764, x44400);
  nand n44404(x44404, x44403, x44402);
  nand n44406(x44406, x44398, x44402);
  nand n44407(x44407, x43747, x85093);
  nand n44409(x44409, x44408, x43749);
  nand n44410(x44410, x44409, x44407);
  nand n44412(x44412, x85095, x44411);
  nand n44413(x44413, x43754, x44410);
  nand n44414(x44414, x44413, x44412);
  nand n44416(x44416, x44407, x44412);
  nand n44417(x44417, x43766, x85097);
  nand n44419(x44419, x44418, x43767);
  nand n44420(x44420, x44419, x44417);
  nand n44422(x44422, x43779, x44421);
  nand n44423(x44423, x43778, x44420);
  nand n44424(x44424, x44423, x44422);
  nand n44426(x44426, x44417, x44422);
  nand n44427(x44427, x43786, x43794);
  nand n44428(x44428, x43785, x43793);
  nand n44429(x44429, x44428, x44427);
  nand n44431(x44431, x43803, x44430);
  nand n44432(x44432, x43802, x44429);
  nand n44433(x44433, x44432, x44431);
  nand n44435(x44435, x44427, x44431);
  nand n44436(x44436, x43780, x85098);
  nand n44438(x44438, x44437, x43782);
  nand n44439(x44439, x44438, x44436);
  nand n44441(x44441, x43795, x44440);
  nand n44443(x44443, x44442, x44439);
  nand n44444(x44444, x44443, x44441);
  nand n44446(x44446, x44436, x44441);
  nand n44447(x44447, x43804, x85100);
  nand n44449(x44449, x44448, x43805);
  nand n44450(x44450, x44449, x44447);
  nand n44452(x44452, x43817, x44451);
  nand n44453(x44453, x43816, x44450);
  nand n44454(x44454, x44453, x44452);
  nand n44456(x44456, x44447, x44452);
  nand n44457(x44457, x43824, x43832);
  nand n44458(x44458, x43823, x43831);
  nand n44459(x44459, x44458, x44457);
  nand n44461(x44461, x43841, x44460);
  nand n44462(x44462, x43840, x44459);
  nand n44463(x44463, x44462, x44461);
  nand n44465(x44465, x44457, x44461);
  nand n44466(x44466, x43818, x85101);
  nand n44468(x44468, x44467, x43820);
  nand n44469(x44469, x44468, x44466);
  nand n44471(x44471, x43833, x44470);
  nand n44473(x44473, x44472, x44469);
  nand n44474(x44474, x44473, x44471);
  nand n44476(x44476, x44466, x44471);
  nand n44477(x44477, x43842, x85103);
  nand n44479(x44479, x44478, x43843);
  nand n44480(x44480, x44479, x44477);
  nand n44482(x44482, x43856, x44481);
  nand n44483(x44483, x43855, x44480);
  nand n44484(x44484, x44483, x44482);
  nand n44486(x44486, x44477, x44482);
  nand n44487(x44487, x43863, x43871);
  nand n44488(x44488, x43862, x43870);
  nand n44489(x44489, x44488, x44487);
  nand n44491(x44491, x43880, x44490);
  nand n44492(x44492, x43879, x44489);
  nand n44493(x44493, x44492, x44491);
  nand n44495(x44495, x44487, x44491);
  nand n44496(x44496, x43857, x85104);
  nand n44498(x44498, x44497, x43859);
  nand n44499(x44499, x44498, x44496);
  nand n44501(x44501, x43872, x44500);
  nand n44503(x44503, x44502, x44499);
  nand n44504(x44504, x44503, x44501);
  nand n44506(x44506, x44496, x44501);
  nand n44507(x44507, x43881, x85106);
  nand n44509(x44509, x44508, x43882);
  nand n44510(x44510, x44509, x44507);
  nand n44512(x44512, x43895, x44511);
  nand n44513(x44513, x43894, x44510);
  nand n44514(x44514, x44513, x44512);
  nand n44516(x44516, x44507, x44512);
  nand n44517(x44517, x43902, x43911);
  nand n44518(x44518, x43901, x43910);
  nand n44519(x44519, x44518, x44517);
  nand n44521(x44521, x43920, x44520);
  nand n44522(x44522, x43919, x44519);
  nand n44523(x44523, x44522, x44521);
  nand n44525(x44525, x44517, x44521);
  nand n44526(x44526, x43896, x85107);
  nand n44528(x44528, x44527, x43898);
  nand n44529(x44529, x44528, x44526);
  nand n44531(x44531, x43912, x44530);
  nand n44533(x44533, x44532, x44529);
  nand n44534(x44534, x44533, x44531);
  nand n44536(x44536, x44526, x44531);
  nand n44537(x44537, x43921, x85109);
  nand n44539(x44539, x44538, x43922);
  nand n44540(x44540, x44539, x44537);
  nand n44542(x44542, x43935, x44541);
  nand n44543(x44543, x43934, x44540);
  nand n44544(x44544, x44543, x44542);
  nand n44546(x44546, x44537, x44542);
  nand n44547(x44547, x43942, x43951);
  nand n44548(x44548, x43941, x43950);
  nand n44549(x44549, x44548, x44547);
  nand n44551(x44551, x43960, x44550);
  nand n44552(x44552, x43959, x44549);
  nand n44553(x44553, x44552, x44551);
  nand n44555(x44555, x44547, x44551);
  nand n44556(x44556, x43936, x85110);
  nand n44558(x44558, x44557, x43938);
  nand n44559(x44559, x44558, x44556);
  nand n44561(x44561, x43952, x44560);
  nand n44563(x44563, x44562, x44559);
  nand n44564(x44564, x44563, x44561);
  nand n44566(x44566, x44556, x44561);
  nand n44567(x44567, x43961, x85112);
  nand n44569(x44569, x44568, x43962);
  nand n44570(x44570, x44569, x44567);
  nand n44572(x44572, x43975, x44571);
  nand n44573(x44573, x43974, x44570);
  nand n44574(x44574, x44573, x44572);
  nand n44576(x44576, x44567, x44572);
  nand n44577(x44577, x43986, x43996);
  nand n44578(x44578, x43985, x43995);
  nand n44579(x44579, x44578, x44577);
  nand n44581(x44581, x44005, x44580);
  nand n44582(x44582, x44004, x44579);
  nand n44583(x44583, x44582, x44581);
  nand n44585(x44585, x44577, x44581);
  nand n44586(x44586, x43976, x43987);
  nand n44589(x44589, x44588, x44587);
  nand n44590(x44590, x44589, x44586);
  nand n44592(x44592, x43997, x44591);
  nand n44594(x44594, x44593, x44590);
  nand n44595(x44595, x44594, x44592);
  nand n44597(x44597, x44006, x44015);
  nand n44600(x44600, x44599, x44598);
  nand n44601(x44601, x44600, x44597);
  nand n44603(x44603, x44026, x44602);
  nand n44604(x44604, x44025, x44601);
  nand n44605(x44605, x44604, x44603);
  nand n44607(x44607, x44036, x44045);
  nand n44608(x44608, x44035, x44044);
  nand n44609(x44609, x44608, x44607);
  nand n44611(x44611, x44053, x44610);
  nand n44612(x44612, x44052, x44609);
  nand n44613(x44613, x44612, x44611);
  nand n44615(x44615, x44071, x85143);
  nand n44616(x44616, x44070, x43473);
  nand n44617(x44617, x44616, x44615);
  nand n44618(x44618, x44075, x85145);
  nand n44619(x44619, x44074, x43477);
  nand n44620(x44620, x44619, x44618);
  nand n44621(x44621, x44082, x85147);
  nand n44622(x44622, x44081, x44078);
  nand n44623(x44623, x44622, x44621);
  nand n44624(x44624, x85116, x85148);
  nand n44625(x44625, x44079, x44076);
  nand n44626(x44626, x44625, x44624);
  nand n44628(x44628, x44093, x85150);
  nand n44629(x44629, x44092, x44085);
  nand n44630(x44630, x44629, x44628);
  nand n44631(x44631, x44094, x85152);
  nand n44633(x44633, x44632, x44083);
  nand n44634(x44634, x44633, x44631);
  nand n44636(x44636, x44105, x85154);
  nand n44637(x44637, x44104, x44097);
  nand n44638(x44638, x44637, x44636);
  nand n44639(x44639, x44106, x85156);
  nand n44641(x44641, x44640, x44095);
  nand n44642(x44642, x44641, x44639);
  nand n44644(x44644, x44117, x85158);
  nand n44645(x44645, x44116, x44109);
  nand n44646(x44646, x44645, x44644);
  nand n44647(x44647, x44118, x85160);
  nand n44649(x44649, x44648, x44107);
  nand n44650(x44650, x44649, x44647);
  nand n44652(x44652, x44129, x85162);
  nand n44653(x44653, x44128, x44121);
  nand n44654(x44654, x44653, x44652);
  nand n44655(x44655, x44130, x85164);
  nand n44657(x44657, x44656, x44119);
  nand n44658(x44658, x44657, x44655);
  nand n44660(x44660, x44141, x85166);
  nand n44661(x44661, x44140, x44133);
  nand n44662(x44662, x44661, x44660);
  nand n44663(x44663, x44142, x85168);
  nand n44665(x44665, x44664, x44131);
  nand n44666(x44666, x44665, x44663);
  nand n44668(x44668, x85122, x44146);
  nand n44669(x44669, x43510, x44145);
  nand n44670(x44670, x44669, x44668);
  nand n44672(x44672, x44154, x44671);
  nand n44673(x44673, x44153, x44670);
  nand n44674(x44674, x44673, x44672);
  nand n44676(x44676, x44668, x44672);
  nand n44677(x44677, x44155, x85170);
  nand n44679(x44679, x44678, x44143);
  nand n44680(x44680, x44679, x44677);
  nand n44682(x44682, x85124, x44159);
  nand n44683(x44683, x43520, x44158);
  nand n44684(x44684, x44683, x44682);
  nand n44686(x44686, x44167, x44685);
  nand n44687(x44687, x44166, x44684);
  nand n44688(x44688, x44687, x44686);
  nand n44690(x44690, x44682, x44686);
  nand n44691(x44691, x44168, x85172);
  nand n44693(x44693, x44692, x44156);
  nand n44694(x44694, x44693, x44691);
  nand n44696(x44696, x85126, x44172);
  nand n44697(x44697, x43530, x44171);
  nand n44698(x44698, x44697, x44696);
  nand n44700(x44700, x44180, x44699);
  nand n44701(x44701, x44179, x44698);
  nand n44702(x44702, x44701, x44700);
  nand n44704(x44704, x44696, x44700);
  nand n44705(x44705, x44181, x85174);
  nand n44707(x44707, x44706, x44169);
  nand n44708(x44708, x44707, x44705);
  nand n44710(x44710, x85128, x44185);
  nand n44711(x44711, x43540, x44184);
  nand n44712(x44712, x44711, x44710);
  nand n44714(x44714, x44193, x44713);
  nand n44715(x44715, x44192, x44712);
  nand n44716(x44716, x44715, x44714);
  nand n44718(x44718, x44710, x44714);
  nand n44719(x44719, x44194, x85176);
  nand n44721(x44721, x44720, x44182);
  nand n44722(x44722, x44721, x44719);
  nand n44724(x44724, x44198, x44202);
  nand n44725(x44725, x44197, x44201);
  nand n44726(x44726, x44725, x44724);
  nand n44728(x44728, x44210, x44727);
  nand n44729(x44729, x44209, x44726);
  nand n44730(x44730, x44729, x44728);
  nand n44732(x44732, x44724, x44728);
  nand n44733(x44733, x85131, x85133);
  nand n44734(x44734, x44195, x44199);
  nand n44735(x44735, x44734, x44733);
  nand n44737(x44737, x44211, x44736);
  nand n44739(x44739, x44738, x44735);
  nand n44740(x44740, x44739, x44737);
  nand n44742(x44742, x44733, x44737);
  nand n44743(x44743, x44219, x44224);
  nand n44744(x44744, x44218, x44223);
  nand n44745(x44745, x44744, x44743);
  nand n44747(x44747, x44232, x44746);
  nand n44748(x44748, x44231, x44745);
  nand n44749(x44749, x44748, x44747);
  nand n44751(x44751, x44743, x44747);
  nand n44752(x44752, x44220, x85135);
  nand n44754(x44754, x44753, x44221);
  nand n44755(x44755, x44754, x44752);
  nand n44757(x44757, x44233, x44756);
  nand n44759(x44759, x44758, x44755);
  nand n44760(x44760, x44759, x44757);
  nand n44762(x44762, x44752, x44757);
  nand n44763(x44763, x44241, x44246);
  nand n44764(x44764, x44240, x44245);
  nand n44765(x44765, x44764, x44763);
  nand n44767(x44767, x44254, x44766);
  nand n44768(x44768, x44253, x44765);
  nand n44769(x44769, x44768, x44767);
  nand n44771(x44771, x44763, x44767);
  nand n44772(x44772, x44242, x85137);
  nand n44774(x44774, x44773, x44243);
  nand n44775(x44775, x44774, x44772);
  nand n44777(x44777, x44255, x44776);
  nand n44779(x44779, x44778, x44775);
  nand n44780(x44780, x44779, x44777);
  nand n44782(x44782, x44772, x44777);
  nand n44783(x44783, x44263, x44268);
  nand n44784(x44784, x44262, x44267);
  nand n44785(x44785, x44784, x44783);
  nand n44787(x44787, x44276, x44786);
  nand n44788(x44788, x44275, x44785);
  nand n44789(x44789, x44788, x44787);
  nand n44791(x44791, x44783, x44787);
  nand n44792(x44792, x44264, x85139);
  nand n44794(x44794, x44793, x44265);
  nand n44795(x44795, x44794, x44792);
  nand n44797(x44797, x44277, x44796);
  nand n44799(x44799, x44798, x44795);
  nand n44800(x44800, x44799, x44797);
  nand n44802(x44802, x44792, x44797);
  nand n44803(x44803, x44285, x44290);
  nand n44804(x44804, x44284, x44289);
  nand n44805(x44805, x44804, x44803);
  nand n44807(x44807, x44298, x44806);
  nand n44808(x44808, x44297, x44805);
  nand n44809(x44809, x44808, x44807);
  nand n44811(x44811, x44803, x44807);
  nand n44812(x44812, x44286, x85141);
  nand n44814(x44814, x44813, x44287);
  nand n44815(x44815, x44814, x44812);
  nand n44817(x44817, x44299, x44816);
  nand n44819(x44819, x44818, x44815);
  nand n44820(x44820, x44819, x44817);
  nand n44822(x44822, x44812, x44817);
  nand n44823(x44823, x44307, x44313);
  nand n44824(x44824, x44306, x44312);
  nand n44825(x44825, x44824, x44823);
  nand n44827(x44827, x44321, x44826);
  nand n44828(x44828, x44320, x44825);
  nand n44829(x44829, x44828, x44827);
  nand n44831(x44831, x44823, x44827);
  nand n44832(x44832, x44308, x85142);
  nand n44834(x44834, x44833, x44310);
  nand n44835(x44835, x44834, x44832);
  nand n44837(x44837, x44322, x44836);
  nand n44839(x44839, x44838, x44835);
  nand n44840(x44840, x44839, x44837);
  nand n44842(x44842, x44832, x44837);
  nand n44843(x44843, x44330, x44340);
  nand n44844(x44844, x44329, x44339);
  nand n44845(x44845, x44844, x44843);
  nand n44847(x44847, x44349, x44846);
  nand n44848(x44848, x44348, x44845);
  nand n44849(x44849, x44848, x44847);
  nand n44851(x44851, x44843, x44847);
  nand n44852(x44852, x44331, x44341);
  nand n44855(x44855, x44854, x44853);
  nand n44856(x44856, x44855, x44852);
  nand n44858(x44858, x44350, x44857);
  nand n44860(x44860, x44859, x44856);
  nand n44861(x44861, x44860, x44858);
  nand n44863(x44863, x44852, x44858);
  nand n44864(x44864, x44358, x44368);
  nand n44865(x44865, x44357, x44367);
  nand n44866(x44866, x44865, x44864);
  nand n44868(x44868, x44377, x44867);
  nand n44869(x44869, x44376, x44866);
  nand n44870(x44870, x44869, x44868);
  nand n44872(x44872, x44864, x44868);
  nand n44873(x44873, x44359, x44369);
  nand n44876(x44876, x44875, x44874);
  nand n44877(x44877, x44876, x44873);
  nand n44879(x44879, x44378, x44878);
  nand n44881(x44881, x44880, x44877);
  nand n44882(x44882, x44881, x44879);
  nand n44884(x44884, x44873, x44879);
  nand n44885(x44885, x44386, x44396);
  nand n44886(x44886, x44385, x44395);
  nand n44887(x44887, x44886, x44885);
  nand n44889(x44889, x44405, x44888);
  nand n44890(x44890, x44404, x44887);
  nand n44891(x44891, x44890, x44889);
  nand n44893(x44893, x44885, x44889);
  nand n44894(x44894, x44387, x44397);
  nand n44897(x44897, x44896, x44895);
  nand n44898(x44898, x44897, x44894);
  nand n44900(x44900, x44406, x44899);
  nand n44902(x44902, x44901, x44898);
  nand n44903(x44903, x44902, x44900);
  nand n44905(x44905, x44894, x44900);
  nand n44906(x44906, x44415, x44425);
  nand n44907(x44907, x44414, x44424);
  nand n44908(x44908, x44907, x44906);
  nand n44910(x44910, x44434, x44909);
  nand n44911(x44911, x44433, x44908);
  nand n44912(x44912, x44911, x44910);
  nand n44914(x44914, x44906, x44910);
  nand n44915(x44915, x44416, x44426);
  nand n44918(x44918, x44917, x44916);
  nand n44919(x44919, x44918, x44915);
  nand n44921(x44921, x44435, x44920);
  nand n44923(x44923, x44922, x44919);
  nand n44924(x44924, x44923, x44921);
  nand n44926(x44926, x44915, x44921);
  nand n44927(x44927, x44445, x44455);
  nand n44928(x44928, x44444, x44454);
  nand n44929(x44929, x44928, x44927);
  nand n44931(x44931, x44464, x44930);
  nand n44932(x44932, x44463, x44929);
  nand n44933(x44933, x44932, x44931);
  nand n44935(x44935, x44927, x44931);
  nand n44936(x44936, x44446, x44456);
  nand n44939(x44939, x44938, x44937);
  nand n44940(x44940, x44939, x44936);
  nand n44942(x44942, x44465, x44941);
  nand n44944(x44944, x44943, x44940);
  nand n44945(x44945, x44944, x44942);
  nand n44947(x44947, x44936, x44942);
  nand n44948(x44948, x44475, x44485);
  nand n44949(x44949, x44474, x44484);
  nand n44950(x44950, x44949, x44948);
  nand n44952(x44952, x44494, x44951);
  nand n44953(x44953, x44493, x44950);
  nand n44954(x44954, x44953, x44952);
  nand n44956(x44956, x44948, x44952);
  nand n44957(x44957, x44476, x44486);
  nand n44960(x44960, x44959, x44958);
  nand n44961(x44961, x44960, x44957);
  nand n44963(x44963, x44495, x44962);
  nand n44965(x44965, x44964, x44961);
  nand n44966(x44966, x44965, x44963);
  nand n44968(x44968, x44957, x44963);
  nand n44969(x44969, x44505, x44515);
  nand n44970(x44970, x44504, x44514);
  nand n44971(x44971, x44970, x44969);
  nand n44973(x44973, x44524, x44972);
  nand n44974(x44974, x44523, x44971);
  nand n44975(x44975, x44974, x44973);
  nand n44977(x44977, x44969, x44973);
  nand n44978(x44978, x44506, x44516);
  nand n44981(x44981, x44980, x44979);
  nand n44982(x44982, x44981, x44978);
  nand n44984(x44984, x44525, x44983);
  nand n44986(x44986, x44985, x44982);
  nand n44987(x44987, x44986, x44984);
  nand n44989(x44989, x44978, x44984);
  nand n44990(x44990, x44535, x44545);
  nand n44991(x44991, x44534, x44544);
  nand n44992(x44992, x44991, x44990);
  nand n44994(x44994, x44554, x44993);
  nand n44995(x44995, x44553, x44992);
  nand n44996(x44996, x44995, x44994);
  nand n44998(x44998, x44990, x44994);
  nand n44999(x44999, x44536, x44546);
  nand n45002(x45002, x45001, x45000);
  nand n45003(x45003, x45002, x44999);
  nand n45005(x45005, x44555, x45004);
  nand n45007(x45007, x45006, x45003);
  nand n45008(x45008, x45007, x45005);
  nand n45010(x45010, x44999, x45005);
  nand n45011(x45011, x44565, x44575);
  nand n45012(x45012, x44564, x44574);
  nand n45013(x45013, x45012, x45011);
  nand n45015(x45015, x44584, x45014);
  nand n45016(x45016, x44583, x45013);
  nand n45017(x45017, x45016, x45015);
  nand n45019(x45019, x45011, x45015);
  nand n45020(x45020, x44566, x44576);
  nand n45023(x45023, x45022, x45021);
  nand n45024(x45024, x45023, x45020);
  nand n45026(x45026, x44585, x45025);
  nand n45028(x45028, x45027, x45024);
  nand n45029(x45029, x45028, x45026);
  nand n45031(x45031, x44596, x44606);
  nand n45032(x45032, x44595, x44605);
  nand n45033(x45033, x45032, x45031);
  nand n45035(x45035, x44614, x45034);
  nand n45036(x45036, x44613, x45033);
  nand n45037(x45037, x45036, x45035);
  nand n45039(x45039, x85144, x85180);
  nand n45040(x45040, x44068, x44615);
  nand n45041(x45041, x45040, x45039);
  nand n45042(x45042, x85146, x85182);
  nand n45043(x45043, x44072, x44618);
  nand n45044(x45044, x45043, x45042);
  nand n45046(x45046, x44627, x85184);
  nand n45047(x45047, x44626, x44621);
  nand n45048(x45048, x45047, x45046);
  nand n45050(x45050, x85149, x85151);
  nand n45051(x45051, x44624, x44628);
  nand n45052(x45052, x45051, x45050);
  nand n45054(x45054, x44635, x45053);
  nand n45055(x45055, x44634, x45052);
  nand n45056(x45056, x45055, x45054);
  nand n45058(x45058, x45050, x45054);
  nand n45059(x45059, x85153, x85155);
  nand n45060(x45060, x44631, x44636);
  nand n45061(x45061, x45060, x45059);
  nand n45063(x45063, x44643, x45062);
  nand n45064(x45064, x44642, x45061);
  nand n45065(x45065, x45064, x45063);
  nand n45067(x45067, x45059, x45063);
  nand n45068(x45068, x85157, x85159);
  nand n45069(x45069, x44639, x44644);
  nand n45070(x45070, x45069, x45068);
  nand n45072(x45072, x44651, x45071);
  nand n45073(x45073, x44650, x45070);
  nand n45074(x45074, x45073, x45072);
  nand n45076(x45076, x45068, x45072);
  nand n45077(x45077, x85161, x85163);
  nand n45078(x45078, x44647, x44652);
  nand n45079(x45079, x45078, x45077);
  nand n45081(x45081, x44659, x45080);
  nand n45082(x45082, x44658, x45079);
  nand n45083(x45083, x45082, x45081);
  nand n45085(x45085, x45077, x45081);
  nand n45086(x45086, x85165, x85167);
  nand n45087(x45087, x44655, x44660);
  nand n45088(x45088, x45087, x45086);
  nand n45090(x45090, x44667, x45089);
  nand n45091(x45091, x44666, x45088);
  nand n45092(x45092, x45091, x45090);
  nand n45094(x45094, x45086, x45090);
  nand n45095(x45095, x44675, x85026);
  nand n45096(x45096, x44674, x40147);
  nand n45097(x45097, x45096, x45095);
  nand n45100(x45100, x85169, x44676);
  nand n45102(x45102, x44663, x45101);
  nand n45103(x45103, x45102, x45100);
  nand n45105(x45105, x44681, x45104);
  nand n45106(x45106, x44680, x45103);
  nand n45107(x45107, x45106, x45105);
  nand n45109(x45109, x45100, x45105);
  nand n45110(x45110, x44689, x85029);
  nand n45111(x45111, x44688, x41287);
  nand n45112(x45112, x45111, x45110);
  nand n45115(x45115, x85171, x44690);
  nand n45117(x45117, x44677, x45116);
  nand n45118(x45118, x45117, x45115);
  nand n45120(x45120, x44695, x45119);
  nand n45121(x45121, x44694, x45118);
  nand n45122(x45122, x45121, x45120);
  nand n45124(x45124, x45115, x45120);
  nand n45125(x45125, x44703, x85032);
  nand n45126(x45126, x44702, x41329);
  nand n45127(x45127, x45126, x45125);
  nand n45130(x45130, x85173, x44704);
  nand n45132(x45132, x44691, x45131);
  nand n45133(x45133, x45132, x45130);
  nand n45135(x45135, x44709, x45134);
  nand n45136(x45136, x44708, x45133);
  nand n45137(x45137, x45136, x45135);
  nand n45139(x45139, x45130, x45135);
  nand n45140(x45140, x44717, x85037);
  nand n45141(x45141, x44716, x42683);
  nand n45142(x45142, x45141, x45140);
  nand n45145(x45145, x85175, x44718);
  nand n45147(x45147, x44705, x45146);
  nand n45148(x45148, x45147, x45145);
  nand n45150(x45150, x44723, x45149);
  nand n45151(x45151, x44722, x45148);
  nand n45152(x45152, x45151, x45150);
  nand n45154(x45154, x45145, x45150);
  nand n45155(x45155, x44731, x85044);
  nand n45156(x45156, x44730, x42711);
  nand n45157(x45157, x45156, x45155);
  nand n45160(x45160, x85177, x44732);
  nand n45162(x45162, x44719, x45161);
  nand n45163(x45163, x45162, x45160);
  nand n45165(x45165, x44741, x45164);
  nand n45166(x45166, x44740, x45163);
  nand n45167(x45167, x45166, x45165);
  nand n45169(x45169, x45160, x45165);
  nand n45170(x45170, x44750, x85051);
  nand n45171(x45171, x44749, x42745);
  nand n45172(x45172, x45171, x45170);
  nand n45175(x45175, x44742, x44751);
  nand n45178(x45178, x45177, x45176);
  nand n45179(x45179, x45178, x45175);
  nand n45181(x45181, x44761, x45180);
  nand n45182(x45182, x44760, x45179);
  nand n45183(x45183, x45182, x45181);
  nand n45185(x45185, x45175, x45181);
  nand n45186(x45186, x44770, x85058);
  nand n45187(x45187, x44769, x42784);
  nand n45188(x45188, x45187, x45186);
  nand n45191(x45191, x44762, x44771);
  nand n45194(x45194, x45193, x45192);
  nand n45195(x45195, x45194, x45191);
  nand n45197(x45197, x44781, x45196);
  nand n45198(x45198, x44780, x45195);
  nand n45199(x45199, x45198, x45197);
  nand n45201(x45201, x45191, x45197);
  nand n45202(x45202, x44790, x85065);
  nand n45203(x45203, x44789, x42824);
  nand n45204(x45204, x45203, x45202);
  nand n45207(x45207, x44782, x44791);
  nand n45210(x45210, x45209, x45208);
  nand n45211(x45211, x45210, x45207);
  nand n45213(x45213, x44801, x45212);
  nand n45214(x45214, x44800, x45211);
  nand n45215(x45215, x45214, x45213);
  nand n45217(x45217, x45207, x45213);
  nand n45218(x45218, x44810, x85071);
  nand n45219(x45219, x44809, x42864);
  nand n45220(x45220, x45219, x45218);
  nand n45223(x45223, x44802, x44811);
  nand n45226(x45226, x45225, x45224);
  nand n45227(x45227, x45226, x45223);
  nand n45229(x45229, x44821, x45228);
  nand n45230(x45230, x44820, x45227);
  nand n45231(x45231, x45230, x45229);
  nand n45233(x45233, x45223, x45229);
  nand n45234(x45234, x44830, x85077);
  nand n45235(x45235, x44829, x43682);
  nand n45236(x45236, x45235, x45234);
  nand n45239(x45239, x44822, x44831);
  nand n45242(x45242, x45241, x45240);
  nand n45243(x45243, x45242, x45239);
  nand n45245(x45245, x44841, x45244);
  nand n45246(x45246, x44840, x45243);
  nand n45247(x45247, x45246, x45245);
  nand n45249(x45249, x45239, x45245);
  nand n45250(x45250, x44850, x85084);
  nand n45251(x45251, x44849, x43709);
  nand n45252(x45252, x45251, x45250);
  nand n45255(x45255, x44842, x44851);
  nand n45258(x45258, x45257, x45256);
  nand n45259(x45259, x45258, x45255);
  nand n45261(x45261, x44862, x45260);
  nand n45262(x45262, x44861, x45259);
  nand n45263(x45263, x45262, x45261);
  nand n45265(x45265, x45255, x45261);
  nand n45266(x45266, x44871, x85091);
  nand n45267(x45267, x44870, x43736);
  nand n45268(x45268, x45267, x45266);
  nand n45271(x45271, x44863, x44872);
  nand n45274(x45274, x45273, x45272);
  nand n45275(x45275, x45274, x45271);
  nand n45277(x45277, x44883, x45276);
  nand n45278(x45278, x44882, x45275);
  nand n45279(x45279, x45278, x45277);
  nand n45281(x45281, x45271, x45277);
  nand n45282(x45282, x44892, x85096);
  nand n45283(x45283, x44891, x43769);
  nand n45284(x45284, x45283, x45282);
  nand n45287(x45287, x44884, x44893);
  nand n45290(x45290, x45289, x45288);
  nand n45291(x45291, x45290, x45287);
  nand n45293(x45293, x44904, x45292);
  nand n45294(x45294, x44903, x45291);
  nand n45295(x45295, x45294, x45293);
  nand n45297(x45297, x45287, x45293);
  nand n45298(x45298, x44913, x85099);
  nand n45299(x45299, x44912, x43807);
  nand n45300(x45300, x45299, x45298);
  nand n45303(x45303, x44905, x44914);
  nand n45306(x45306, x45305, x45304);
  nand n45307(x45307, x45306, x45303);
  nand n45309(x45309, x44925, x45308);
  nand n45310(x45310, x44924, x45307);
  nand n45311(x45311, x45310, x45309);
  nand n45313(x45313, x45303, x45309);
  nand n45314(x45314, x44934, x85102);
  nand n45315(x45315, x44933, x43845);
  nand n45316(x45316, x45315, x45314);
  nand n45319(x45319, x44926, x44935);
  nand n45322(x45322, x45321, x45320);
  nand n45323(x45323, x45322, x45319);
  nand n45325(x45325, x44946, x45324);
  nand n45326(x45326, x44945, x45323);
  nand n45327(x45327, x45326, x45325);
  nand n45329(x45329, x45319, x45325);
  nand n45330(x45330, x44955, x85105);
  nand n45331(x45331, x44954, x43884);
  nand n45332(x45332, x45331, x45330);
  nand n45335(x45335, x44947, x44956);
  nand n45338(x45338, x45337, x45336);
  nand n45339(x45339, x45338, x45335);
  nand n45341(x45341, x44967, x45340);
  nand n45342(x45342, x44966, x45339);
  nand n45343(x45343, x45342, x45341);
  nand n45345(x45345, x45335, x45341);
  nand n45346(x45346, x44976, x85108);
  nand n45347(x45347, x44975, x43924);
  nand n45348(x45348, x45347, x45346);
  nand n45351(x45351, x44968, x44977);
  nand n45354(x45354, x45353, x45352);
  nand n45355(x45355, x45354, x45351);
  nand n45357(x45357, x44988, x45356);
  nand n45358(x45358, x44987, x45355);
  nand n45359(x45359, x45358, x45357);
  nand n45361(x45361, x45351, x45357);
  nand n45362(x45362, x44997, x85111);
  nand n45363(x45363, x44996, x43964);
  nand n45364(x45364, x45363, x45362);
  nand n45367(x45367, x44989, x44998);
  nand n45370(x45370, x45369, x45368);
  nand n45371(x45371, x45370, x45367);
  nand n45373(x45373, x45009, x45372);
  nand n45374(x45374, x45008, x45371);
  nand n45375(x45375, x45374, x45373);
  nand n45377(x45377, x45367, x45373);
  nand n45378(x45378, x45018, x44014);
  nand n45379(x45379, x45017, x44013);
  nand n45380(x45380, x45379, x45378);
  nand n45383(x45383, x45010, x45019);
  nand n45386(x45386, x45385, x45384);
  nand n45387(x45387, x45386, x45383);
  nand n45389(x45389, x45030, x45388);
  nand n45390(x45390, x45029, x45387);
  nand n45391(x45391, x45390, x45389);
  nand n45393(x45393, x45038, x44061);
  nand n45394(x45394, x45037, x44060);
  nand n45395(x45395, x45394, x45393);
  nand n45397(x45397, x85178, x85190);
  nand n45398(x45398, x44067, x44062);
  nand n45399(x45399, x45398, x45397);
  nand n45400(x45400, x45045, x85193);
  nand n45401(x45401, x45044, x45039);
  nand n45402(x45402, x45401, x45400);
  nand n45403(x45403, x45049, x85195);
  nand n45404(x45404, x45048, x45042);
  nand n45405(x45405, x45404, x45403);
  nand n45407(x45407, x45057, x85197);
  nand n45408(x45408, x45056, x45046);
  nand n45409(x45409, x45408, x45407);
  nand n45412(x45412, x45066, x45058);
  nand n45413(x45413, x45065, x45411);
  nand n45414(x45414, x45413, x45412);
  nand n45417(x45417, x45075, x45067);
  nand n45418(x45418, x45074, x45416);
  nand n45419(x45419, x45418, x45417);
  nand n45422(x45422, x45084, x45076);
  nand n45423(x45423, x45083, x45421);
  nand n45424(x45424, x45423, x45422);
  nand n45427(x45427, x45093, x45085);
  nand n45428(x45428, x45092, x45426);
  nand n45429(x45429, x45428, x45427);
  nand n45431(x45431, x45094, x45099);
  nand n45433(x45433, x45432, x45095);
  nand n45434(x45434, x45433, x45431);
  nand n45436(x45436, x45108, x45435);
  nand n45437(x45437, x45107, x45434);
  nand n45438(x45438, x45437, x45436);
  nand n45440(x45440, x45431, x45436);
  nand n45441(x45441, x45109, x45114);
  nand n45443(x45443, x45442, x45110);
  nand n45444(x45444, x45443, x45441);
  nand n45446(x45446, x45123, x45445);
  nand n45447(x45447, x45122, x45444);
  nand n45448(x45448, x45447, x45446);
  nand n45450(x45450, x45441, x45446);
  nand n45451(x45451, x45124, x45129);
  nand n45453(x45453, x45452, x45125);
  nand n45454(x45454, x45453, x45451);
  nand n45456(x45456, x45138, x45455);
  nand n45457(x45457, x45137, x45454);
  nand n45458(x45458, x45457, x45456);
  nand n45460(x45460, x45451, x45456);
  nand n45461(x45461, x45139, x45144);
  nand n45463(x45463, x45462, x45140);
  nand n45464(x45464, x45463, x45461);
  nand n45466(x45466, x45153, x45465);
  nand n45467(x45467, x45152, x45464);
  nand n45468(x45468, x45467, x45466);
  nand n45470(x45470, x45461, x45466);
  nand n45471(x45471, x45154, x45159);
  nand n45473(x45473, x45472, x45155);
  nand n45474(x45474, x45473, x45471);
  nand n45476(x45476, x45168, x45475);
  nand n45477(x45477, x45167, x45474);
  nand n45478(x45478, x45477, x45476);
  nand n45480(x45480, x45471, x45476);
  nand n45481(x45481, x45169, x45174);
  nand n45483(x45483, x45482, x45170);
  nand n45484(x45484, x45483, x45481);
  nand n45486(x45486, x45184, x45485);
  nand n45487(x45487, x45183, x45484);
  nand n45488(x45488, x45487, x45486);
  nand n45490(x45490, x45481, x45486);
  nand n45491(x45491, x45185, x45190);
  nand n45493(x45493, x45492, x45186);
  nand n45494(x45494, x45493, x45491);
  nand n45496(x45496, x45200, x45495);
  nand n45497(x45497, x45199, x45494);
  nand n45498(x45498, x45497, x45496);
  nand n45500(x45500, x45491, x45496);
  nand n45501(x45501, x45201, x45206);
  nand n45503(x45503, x45502, x45202);
  nand n45504(x45504, x45503, x45501);
  nand n45506(x45506, x45216, x45505);
  nand n45507(x45507, x45215, x45504);
  nand n45508(x45508, x45507, x45506);
  nand n45510(x45510, x45501, x45506);
  nand n45511(x45511, x45217, x45222);
  nand n45513(x45513, x45512, x45218);
  nand n45514(x45514, x45513, x45511);
  nand n45516(x45516, x45232, x45515);
  nand n45517(x45517, x45231, x45514);
  nand n45518(x45518, x45517, x45516);
  nand n45520(x45520, x45511, x45516);
  nand n45521(x45521, x45233, x45238);
  nand n45523(x45523, x45522, x45234);
  nand n45524(x45524, x45523, x45521);
  nand n45526(x45526, x45248, x45525);
  nand n45527(x45527, x45247, x45524);
  nand n45528(x45528, x45527, x45526);
  nand n45530(x45530, x45521, x45526);
  nand n45531(x45531, x45249, x45254);
  nand n45533(x45533, x45532, x45250);
  nand n45534(x45534, x45533, x45531);
  nand n45536(x45536, x45264, x45535);
  nand n45537(x45537, x45263, x45534);
  nand n45538(x45538, x45537, x45536);
  nand n45540(x45540, x45531, x45536);
  nand n45541(x45541, x45265, x45270);
  nand n45543(x45543, x45542, x45266);
  nand n45544(x45544, x45543, x45541);
  nand n45546(x45546, x45280, x45545);
  nand n45547(x45547, x45279, x45544);
  nand n45548(x45548, x45547, x45546);
  nand n45550(x45550, x45541, x45546);
  nand n45551(x45551, x45281, x45286);
  nand n45553(x45553, x45552, x45282);
  nand n45554(x45554, x45553, x45551);
  nand n45556(x45556, x45296, x45555);
  nand n45557(x45557, x45295, x45554);
  nand n45558(x45558, x45557, x45556);
  nand n45560(x45560, x45551, x45556);
  nand n45561(x45561, x45297, x45302);
  nand n45563(x45563, x45562, x45298);
  nand n45564(x45564, x45563, x45561);
  nand n45566(x45566, x45312, x45565);
  nand n45567(x45567, x45311, x45564);
  nand n45568(x45568, x45567, x45566);
  nand n45570(x45570, x45561, x45566);
  nand n45571(x45571, x45313, x45318);
  nand n45573(x45573, x45572, x45314);
  nand n45574(x45574, x45573, x45571);
  nand n45576(x45576, x45328, x45575);
  nand n45577(x45577, x45327, x45574);
  nand n45578(x45578, x45577, x45576);
  nand n45580(x45580, x45571, x45576);
  nand n45581(x45581, x45329, x45334);
  nand n45583(x45583, x45582, x45330);
  nand n45584(x45584, x45583, x45581);
  nand n45586(x45586, x45344, x45585);
  nand n45587(x45587, x45343, x45584);
  nand n45588(x45588, x45587, x45586);
  nand n45590(x45590, x45581, x45586);
  nand n45591(x45591, x45345, x45350);
  nand n45593(x45593, x45592, x45346);
  nand n45594(x45594, x45593, x45591);
  nand n45596(x45596, x45360, x45595);
  nand n45597(x45597, x45359, x45594);
  nand n45598(x45598, x45597, x45596);
  nand n45600(x45600, x45591, x45596);
  nand n45601(x45601, x45361, x45366);
  nand n45603(x45603, x45602, x45362);
  nand n45604(x45604, x45603, x45601);
  nand n45606(x45606, x45376, x45605);
  nand n45607(x45607, x45375, x45604);
  nand n45608(x45608, x45607, x45606);
  nand n45610(x45610, x45601, x45606);
  nand n45611(x45611, x45377, x45382);
  nand n45613(x45613, x45612, x45378);
  nand n45614(x45614, x45613, x45611);
  nand n45616(x45616, x45392, x45615);
  nand n45617(x45617, x45391, x45614);
  nand n45618(x45618, x45617, x45616);
  nand n45620(x45620, x85191, x85192);
  nand n45621(x45621, x45397, x44065);
  nand n45622(x45622, x45621, x45620);
  nand n45624(x45624, x85179, x45623);
  nand n45625(x45625, x44617, x45622);
  nand n45626(x45626, x45625, x45624);
  nand n45627(x45627, x45620, x45624);
  nand n45628(x45628, x85181, x85203);
  nand n45629(x45629, x44620, x45041);
  nand n45630(x45630, x45629, x45628);
  nand n45632(x45632, x85183, x85205);
  nand n45633(x45633, x44623, x45402);
  nand n45634(x45634, x45633, x45632);
  nand n45636(x45636, x85194, x45406);
  nand n45637(x45637, x45400, x45405);
  nand n45638(x45638, x45637, x45636);
  nand n45640(x45640, x85185, x45639);
  nand n45641(x45641, x44630, x45638);
  nand n45642(x45642, x45641, x45640);
  nand n45644(x45644, x45636, x45640);
  nand n45645(x45645, x85196, x45410);
  nand n45646(x45646, x45403, x45409);
  nand n45647(x45647, x45646, x45645);
  nand n45649(x45649, x85186, x45648);
  nand n45650(x45650, x44638, x45647);
  nand n45651(x45651, x45650, x45649);
  nand n45653(x45653, x45645, x45649);
  nand n45654(x45654, x85198, x45415);
  nand n45655(x45655, x45407, x45414);
  nand n45656(x45656, x45655, x45654);
  nand n45658(x45658, x85187, x45657);
  nand n45659(x45659, x44646, x45656);
  nand n45660(x45660, x45659, x45658);
  nand n45662(x45662, x45654, x45658);
  nand n45663(x45663, x85199, x45420);
  nand n45664(x45664, x45412, x45419);
  nand n45665(x45665, x45664, x45663);
  nand n45667(x45667, x85188, x45666);
  nand n45668(x45668, x44654, x45665);
  nand n45669(x45669, x45668, x45667);
  nand n45671(x45671, x45663, x45667);
  nand n45672(x45672, x85200, x45425);
  nand n45673(x45673, x45417, x45424);
  nand n45674(x45674, x45673, x45672);
  nand n45676(x45676, x85189, x45675);
  nand n45677(x45677, x44662, x45674);
  nand n45678(x45678, x45677, x45676);
  nand n45680(x45680, x45672, x45676);
  nand n45681(x45681, x85201, x45430);
  nand n45682(x45682, x45422, x45429);
  nand n45683(x45683, x45682, x45681);
  nand n45685(x45685, x45098, x45684);
  nand n45686(x45686, x45097, x45683);
  nand n45687(x45687, x45686, x45685);
  nand n45689(x45689, x45681, x45685);
  nand n45690(x45690, x85202, x45439);
  nand n45691(x45691, x45427, x45438);
  nand n45692(x45692, x45691, x45690);
  nand n45694(x45694, x45113, x45693);
  nand n45695(x45695, x45112, x45692);
  nand n45696(x45696, x45695, x45694);
  nand n45698(x45698, x45690, x45694);
  nand n45699(x45699, x45440, x45449);
  nand n45701(x45701, x45700, x45448);
  nand n45702(x45702, x45701, x45699);
  nand n45704(x45704, x45128, x45703);
  nand n45705(x45705, x45127, x45702);
  nand n45706(x45706, x45705, x45704);
  nand n45708(x45708, x45699, x45704);
  nand n45709(x45709, x45450, x45459);
  nand n45711(x45711, x45710, x45458);
  nand n45712(x45712, x45711, x45709);
  nand n45714(x45714, x45143, x45713);
  nand n45715(x45715, x45142, x45712);
  nand n45716(x45716, x45715, x45714);
  nand n45718(x45718, x45709, x45714);
  nand n45719(x45719, x45460, x45469);
  nand n45721(x45721, x45720, x45468);
  nand n45722(x45722, x45721, x45719);
  nand n45724(x45724, x45158, x45723);
  nand n45725(x45725, x45157, x45722);
  nand n45726(x45726, x45725, x45724);
  nand n45728(x45728, x45719, x45724);
  nand n45729(x45729, x45470, x45479);
  nand n45731(x45731, x45730, x45478);
  nand n45732(x45732, x45731, x45729);
  nand n45734(x45734, x45173, x45733);
  nand n45735(x45735, x45172, x45732);
  nand n45736(x45736, x45735, x45734);
  nand n45738(x45738, x45729, x45734);
  nand n45739(x45739, x45480, x45489);
  nand n45741(x45741, x45740, x45488);
  nand n45742(x45742, x45741, x45739);
  nand n45744(x45744, x45189, x45743);
  nand n45745(x45745, x45188, x45742);
  nand n45746(x45746, x45745, x45744);
  nand n45748(x45748, x45739, x45744);
  nand n45749(x45749, x45490, x45499);
  nand n45751(x45751, x45750, x45498);
  nand n45752(x45752, x45751, x45749);
  nand n45754(x45754, x45205, x45753);
  nand n45755(x45755, x45204, x45752);
  nand n45756(x45756, x45755, x45754);
  nand n45758(x45758, x45749, x45754);
  nand n45759(x45759, x45500, x45509);
  nand n45761(x45761, x45760, x45508);
  nand n45762(x45762, x45761, x45759);
  nand n45764(x45764, x45221, x45763);
  nand n45765(x45765, x45220, x45762);
  nand n45766(x45766, x45765, x45764);
  nand n45768(x45768, x45759, x45764);
  nand n45769(x45769, x45510, x45519);
  nand n45771(x45771, x45770, x45518);
  nand n45772(x45772, x45771, x45769);
  nand n45774(x45774, x45237, x45773);
  nand n45775(x45775, x45236, x45772);
  nand n45776(x45776, x45775, x45774);
  nand n45778(x45778, x45769, x45774);
  nand n45779(x45779, x45520, x45529);
  nand n45781(x45781, x45780, x45528);
  nand n45782(x45782, x45781, x45779);
  nand n45784(x45784, x45253, x45783);
  nand n45785(x45785, x45252, x45782);
  nand n45786(x45786, x45785, x45784);
  nand n45788(x45788, x45779, x45784);
  nand n45789(x45789, x45530, x45539);
  nand n45791(x45791, x45790, x45538);
  nand n45792(x45792, x45791, x45789);
  nand n45794(x45794, x45269, x45793);
  nand n45795(x45795, x45268, x45792);
  nand n45796(x45796, x45795, x45794);
  nand n45798(x45798, x45789, x45794);
  nand n45799(x45799, x45540, x45549);
  nand n45801(x45801, x45800, x45548);
  nand n45802(x45802, x45801, x45799);
  nand n45804(x45804, x45285, x45803);
  nand n45805(x45805, x45284, x45802);
  nand n45806(x45806, x45805, x45804);
  nand n45808(x45808, x45799, x45804);
  nand n45809(x45809, x45550, x45559);
  nand n45811(x45811, x45810, x45558);
  nand n45812(x45812, x45811, x45809);
  nand n45814(x45814, x45301, x45813);
  nand n45815(x45815, x45300, x45812);
  nand n45816(x45816, x45815, x45814);
  nand n45818(x45818, x45809, x45814);
  nand n45819(x45819, x45560, x45569);
  nand n45821(x45821, x45820, x45568);
  nand n45822(x45822, x45821, x45819);
  nand n45824(x45824, x45317, x45823);
  nand n45825(x45825, x45316, x45822);
  nand n45826(x45826, x45825, x45824);
  nand n45828(x45828, x45819, x45824);
  nand n45829(x45829, x45570, x45579);
  nand n45831(x45831, x45830, x45578);
  nand n45832(x45832, x45831, x45829);
  nand n45834(x45834, x45333, x45833);
  nand n45835(x45835, x45332, x45832);
  nand n45836(x45836, x45835, x45834);
  nand n45838(x45838, x45829, x45834);
  nand n45839(x45839, x45580, x45589);
  nand n45841(x45841, x45840, x45588);
  nand n45842(x45842, x45841, x45839);
  nand n45844(x45844, x45349, x45843);
  nand n45845(x45845, x45348, x45842);
  nand n45846(x45846, x45845, x45844);
  nand n45848(x45848, x45839, x45844);
  nand n45849(x45849, x45590, x45599);
  nand n45851(x45851, x45850, x45598);
  nand n45852(x45852, x45851, x45849);
  nand n45854(x45854, x45365, x45853);
  nand n45855(x45855, x45364, x45852);
  nand n45856(x45856, x45855, x45854);
  nand n45858(x45858, x45849, x45854);
  nand n45859(x45859, x45600, x45609);
  nand n45861(x45861, x45860, x45608);
  nand n45862(x45862, x45861, x45859);
  nand n45864(x45864, x45381, x45863);
  nand n45865(x45865, x45380, x45862);
  nand n45866(x45866, x45865, x45864);
  nand n45868(x45868, x45859, x45864);
  nand n45869(x45869, x45610, x45619);
  nand n45871(x45871, x45870, x45618);
  nand n45872(x45872, x45871, x45869);
  nand n45874(x45874, x45396, x45873);
  nand n45875(x45875, x45395, x45872);
  nand n45876(x45876, x45875, x45874);
  nand n45878(x45878, x45627, x45631);
  nand n45880(x45880, x45879, x45630);
  nand n45881(x45881, x45880, x45878);
  nand n45882(x45882, x85204, x45635);
  nand n45883(x45883, x45628, x45634);
  nand n45884(x45884, x45883, x45882);
  nand n45886(x45886, x85206, x45643);
  nand n45887(x45887, x45632, x45642);
  nand n45888(x45888, x45887, x45886);
  nand n45890(x45890, x45644, x45652);
  nand n45892(x45892, x45891, x45651);
  nand n45893(x45893, x45892, x45890);
  nand n45895(x45895, x45653, x45661);
  nand n45897(x45897, x45896, x45660);
  nand n45898(x45898, x45897, x45895);
  nand n45900(x45900, x45662, x45670);
  nand n45902(x45902, x45901, x45669);
  nand n45903(x45903, x45902, x45900);
  nand n45905(x45905, x45671, x45679);
  nand n45907(x45907, x45906, x45678);
  nand n45908(x45908, x45907, x45905);
  nand n45910(x45910, x45680, x45688);
  nand n45912(x45912, x45911, x45687);
  nand n45913(x45913, x45912, x45910);
  nand n45915(x45915, x45689, x45697);
  nand n45917(x45917, x45916, x45696);
  nand n45918(x45918, x45917, x45915);
  nand n45920(x45920, x45698, x45707);
  nand n45922(x45922, x45921, x45706);
  nand n45923(x45923, x45922, x45920);
  nand n45925(x45925, x45708, x45717);
  nand n45927(x45927, x45926, x45716);
  nand n45928(x45928, x45927, x45925);
  nand n45930(x45930, x45718, x45727);
  nand n45932(x45932, x45931, x45726);
  nand n45933(x45933, x45932, x45930);
  nand n45935(x45935, x45728, x45737);
  nand n45937(x45937, x45936, x45736);
  nand n45938(x45938, x45937, x45935);
  nand n45940(x45940, x45738, x45747);
  nand n45942(x45942, x45941, x45746);
  nand n45943(x45943, x45942, x45940);
  nand n45945(x45945, x45748, x45757);
  nand n45947(x45947, x45946, x45756);
  nand n45948(x45948, x45947, x45945);
  nand n45950(x45950, x45758, x45767);
  nand n45952(x45952, x45951, x45766);
  nand n45953(x45953, x45952, x45950);
  nand n45955(x45955, x45768, x45777);
  nand n45957(x45957, x45956, x45776);
  nand n45958(x45958, x45957, x45955);
  nand n45960(x45960, x45778, x45787);
  nand n45962(x45962, x45961, x45786);
  nand n45963(x45963, x45962, x45960);
  nand n45965(x45965, x45788, x45797);
  nand n45967(x45967, x45966, x45796);
  nand n45968(x45968, x45967, x45965);
  nand n45970(x45970, x45798, x45807);
  nand n45972(x45972, x45971, x45806);
  nand n45973(x45973, x45972, x45970);
  nand n45975(x45975, x45808, x45817);
  nand n45977(x45977, x45976, x45816);
  nand n45978(x45978, x45977, x45975);
  nand n45980(x45980, x45818, x45827);
  nand n45982(x45982, x45981, x45826);
  nand n45983(x45983, x45982, x45980);
  nand n45985(x45985, x45828, x45837);
  nand n45987(x45987, x45986, x45836);
  nand n45988(x45988, x45987, x45985);
  nand n45990(x45990, x45838, x45847);
  nand n45992(x45992, x45991, x45846);
  nand n45993(x45993, x45992, x45990);
  nand n45995(x45995, x45848, x45857);
  nand n45997(x45997, x45996, x45856);
  nand n45998(x45998, x45997, x45995);
  nand n46000(x46000, x45858, x45867);
  nand n46002(x46002, x46001, x45866);
  nand n46003(x46003, x46002, x46000);
  nand n46005(x46005, x45868, x45877);
  nand n46007(x46007, x46006, x45876);
  nand n46008(x46008, x46007, x46005);
  nand n46035(x46035, x45885, x46010);
  nand n46036(x46036, x46035, x45882);
  nand n46037(x46037, x45889, x46011);
  nand n46038(x46038, x46037, x45886);
  nand n46039(x46039, x45889, x45885);
  nand n46041(x46041, x45894, x46012);
  nand n46042(x46042, x46041, x45890);
  nand n46043(x46043, x45894, x45889);
  nand n46045(x46045, x45899, x46013);
  nand n46046(x46046, x46045, x45895);
  nand n46047(x46047, x45899, x45894);
  nand n46049(x46049, x45904, x46014);
  nand n46050(x46050, x46049, x45900);
  nand n46051(x46051, x45904, x45899);
  nand n46053(x46053, x45909, x46015);
  nand n46054(x46054, x46053, x45905);
  nand n46055(x46055, x45909, x45904);
  nand n46057(x46057, x45914, x46016);
  nand n46058(x46058, x46057, x45910);
  nand n46059(x46059, x45914, x45909);
  nand n46061(x46061, x45919, x46017);
  nand n46062(x46062, x46061, x45915);
  nand n46063(x46063, x45919, x45914);
  nand n46065(x46065, x45924, x46018);
  nand n46066(x46066, x46065, x45920);
  nand n46067(x46067, x45924, x45919);
  nand n46069(x46069, x45929, x46019);
  nand n46070(x46070, x46069, x45925);
  nand n46071(x46071, x45929, x45924);
  nand n46073(x46073, x45934, x46020);
  nand n46074(x46074, x46073, x45930);
  nand n46075(x46075, x45934, x45929);
  nand n46077(x46077, x45939, x46021);
  nand n46078(x46078, x46077, x45935);
  nand n46079(x46079, x45939, x45934);
  nand n46081(x46081, x45944, x46022);
  nand n46082(x46082, x46081, x45940);
  nand n46083(x46083, x45944, x45939);
  nand n46085(x46085, x45949, x46023);
  nand n46086(x46086, x46085, x45945);
  nand n46087(x46087, x45949, x45944);
  nand n46089(x46089, x45954, x46024);
  nand n46090(x46090, x46089, x45950);
  nand n46091(x46091, x45954, x45949);
  nand n46093(x46093, x45959, x46025);
  nand n46094(x46094, x46093, x45955);
  nand n46095(x46095, x45959, x45954);
  nand n46097(x46097, x45964, x46026);
  nand n46098(x46098, x46097, x45960);
  nand n46099(x46099, x45964, x45959);
  nand n46101(x46101, x45969, x46027);
  nand n46102(x46102, x46101, x45965);
  nand n46103(x46103, x45969, x45964);
  nand n46105(x46105, x45974, x46028);
  nand n46106(x46106, x46105, x45970);
  nand n46107(x46107, x45974, x45969);
  nand n46109(x46109, x45979, x46029);
  nand n46110(x46110, x46109, x45975);
  nand n46111(x46111, x45979, x45974);
  nand n46113(x46113, x45984, x46030);
  nand n46114(x46114, x46113, x45980);
  nand n46115(x46115, x45984, x45979);
  nand n46117(x46117, x45989, x46031);
  nand n46118(x46118, x46117, x45985);
  nand n46119(x46119, x45989, x45984);
  nand n46121(x46121, x45994, x46032);
  nand n46122(x46122, x46121, x45990);
  nand n46123(x46123, x45994, x45989);
  nand n46125(x46125, x45999, x46033);
  nand n46126(x46126, x46125, x45995);
  nand n46127(x46127, x45999, x45994);
  nand n46129(x46129, x46004, x46034);
  nand n46130(x46130, x46129, x46000);
  nand n46131(x46131, x46004, x45999);
  nand n46134(x46134, x46040, x46010);
  nand n46136(x46136, x46134, x46135);
  nand n46137(x46137, x46044, x46036);
  nand n46139(x46139, x46137, x46138);
  nand n46140(x46140, x46048, x46038);
  nand n46142(x46142, x46140, x46141);
  nand n46143(x46143, x46048, x46040);
  nand n46145(x46145, x46052, x46042);
  nand n46147(x46147, x46145, x46146);
  nand n46148(x46148, x46052, x46044);
  nand n46150(x46150, x46056, x46046);
  nand n46152(x46152, x46150, x46151);
  nand n46153(x46153, x46056, x46048);
  nand n46155(x46155, x46060, x46050);
  nand n46157(x46157, x46155, x46156);
  nand n46158(x46158, x46060, x46052);
  nand n46160(x46160, x46064, x46054);
  nand n46162(x46162, x46160, x46161);
  nand n46163(x46163, x46064, x46056);
  nand n46165(x46165, x46068, x46058);
  nand n46167(x46167, x46165, x46166);
  nand n46168(x46168, x46068, x46060);
  nand n46170(x46170, x46072, x46062);
  nand n46172(x46172, x46170, x46171);
  nand n46173(x46173, x46072, x46064);
  nand n46175(x46175, x46076, x46066);
  nand n46177(x46177, x46175, x46176);
  nand n46178(x46178, x46076, x46068);
  nand n46180(x46180, x46080, x46070);
  nand n46182(x46182, x46180, x46181);
  nand n46183(x46183, x46080, x46072);
  nand n46185(x46185, x46084, x46074);
  nand n46187(x46187, x46185, x46186);
  nand n46188(x46188, x46084, x46076);
  nand n46190(x46190, x46088, x46078);
  nand n46192(x46192, x46190, x46191);
  nand n46193(x46193, x46088, x46080);
  nand n46195(x46195, x46092, x46082);
  nand n46197(x46197, x46195, x46196);
  nand n46198(x46198, x46092, x46084);
  nand n46200(x46200, x46096, x46086);
  nand n46202(x46202, x46200, x46201);
  nand n46203(x46203, x46096, x46088);
  nand n46205(x46205, x46100, x46090);
  nand n46207(x46207, x46205, x46206);
  nand n46208(x46208, x46100, x46092);
  nand n46210(x46210, x46104, x46094);
  nand n46212(x46212, x46210, x46211);
  nand n46213(x46213, x46104, x46096);
  nand n46215(x46215, x46108, x46098);
  nand n46217(x46217, x46215, x46216);
  nand n46218(x46218, x46108, x46100);
  nand n46220(x46220, x46112, x46102);
  nand n46222(x46222, x46220, x46221);
  nand n46223(x46223, x46112, x46104);
  nand n46225(x46225, x46116, x46106);
  nand n46227(x46227, x46225, x46226);
  nand n46228(x46228, x46116, x46108);
  nand n46230(x46230, x46120, x46110);
  nand n46232(x46232, x46230, x46231);
  nand n46233(x46233, x46120, x46112);
  nand n46235(x46235, x46124, x46114);
  nand n46237(x46237, x46235, x46236);
  nand n46238(x46238, x46124, x46116);
  nand n46240(x46240, x46128, x46118);
  nand n46242(x46242, x46240, x46241);
  nand n46243(x46243, x46128, x46120);
  nand n46245(x46245, x46132, x46122);
  nand n46247(x46247, x46245, x46246);
  nand n46248(x46248, x46132, x46124);
  nand n46252(x46252, x46144, x46010);
  nand n46254(x46254, x46252, x46253);
  nand n46255(x46255, x46149, x46036);
  nand n46257(x46257, x46255, x46256);
  nand n46258(x46258, x46154, x46136);
  nand n46260(x46260, x46258, x46259);
  nand n46261(x46261, x46159, x46139);
  nand n46263(x46263, x46261, x46262);
  nand n46264(x46264, x46164, x46142);
  nand n46266(x46266, x46264, x46265);
  nand n46267(x46267, x46164, x46144);
  nand n46269(x46269, x46169, x46147);
  nand n46271(x46271, x46269, x46270);
  nand n46272(x46272, x46169, x46149);
  nand n46274(x46274, x46174, x46152);
  nand n46276(x46276, x46274, x46275);
  nand n46277(x46277, x46174, x46154);
  nand n46279(x46279, x46179, x46157);
  nand n46281(x46281, x46279, x46280);
  nand n46282(x46282, x46179, x46159);
  nand n46284(x46284, x46184, x46162);
  nand n46286(x46286, x46284, x46285);
  nand n46287(x46287, x46184, x46164);
  nand n46289(x46289, x46189, x46167);
  nand n46291(x46291, x46289, x46290);
  nand n46292(x46292, x46189, x46169);
  nand n46294(x46294, x46194, x46172);
  nand n46296(x46296, x46294, x46295);
  nand n46297(x46297, x46194, x46174);
  nand n46299(x46299, x46199, x46177);
  nand n46301(x46301, x46299, x46300);
  nand n46302(x46302, x46199, x46179);
  nand n46304(x46304, x46204, x46182);
  nand n46306(x46306, x46304, x46305);
  nand n46307(x46307, x46204, x46184);
  nand n46309(x46309, x46209, x46187);
  nand n46311(x46311, x46309, x46310);
  nand n46312(x46312, x46209, x46189);
  nand n46314(x46314, x46214, x46192);
  nand n46316(x46316, x46314, x46315);
  nand n46317(x46317, x46214, x46194);
  nand n46319(x46319, x46219, x46197);
  nand n46321(x46321, x46319, x46320);
  nand n46322(x46322, x46219, x46199);
  nand n46324(x46324, x46224, x46202);
  nand n46326(x46326, x46324, x46325);
  nand n46327(x46327, x46224, x46204);
  nand n46329(x46329, x46229, x46207);
  nand n46331(x46331, x46329, x46330);
  nand n46332(x46332, x46229, x46209);
  nand n46334(x46334, x46234, x46212);
  nand n46336(x46336, x46334, x46335);
  nand n46337(x46337, x46234, x46214);
  nand n46339(x46339, x46239, x46217);
  nand n46341(x46341, x46339, x46340);
  nand n46342(x46342, x46239, x46219);
  nand n46344(x46344, x46244, x46222);
  nand n46346(x46346, x46344, x46345);
  nand n46347(x46347, x46244, x46224);
  nand n46349(x46349, x46249, x46227);
  nand n46351(x46351, x46349, x46350);
  nand n46352(x46352, x46249, x46229);
  nand n46358(x46358, x46268, x46010);
  nand n46360(x46360, x46358, x46359);
  nand n46361(x46361, x46273, x46036);
  nand n46363(x46363, x46361, x46362);
  nand n46364(x46364, x46278, x46136);
  nand n46366(x46366, x46364, x46365);
  nand n46367(x46367, x46283, x46139);
  nand n46369(x46369, x46367, x46368);
  nand n46370(x46370, x46288, x46254);
  nand n46372(x46372, x46370, x46371);
  nand n46373(x46373, x46293, x46257);
  nand n46375(x46375, x46373, x46374);
  nand n46376(x46376, x46298, x46260);
  nand n46378(x46378, x46376, x46377);
  nand n46379(x46379, x46303, x46263);
  nand n46381(x46381, x46379, x46380);
  nand n46382(x46382, x46308, x46266);
  nand n46384(x46384, x46382, x46383);
  nand n46385(x46385, x46308, x46268);
  nand n46387(x46387, x46313, x46271);
  nand n46389(x46389, x46387, x46388);
  nand n46390(x46390, x46313, x46273);
  nand n46392(x46392, x46318, x46276);
  nand n46394(x46394, x46392, x46393);
  nand n46395(x46395, x46318, x46278);
  nand n46397(x46397, x46323, x46281);
  nand n46399(x46399, x46397, x46398);
  nand n46400(x46400, x46323, x46283);
  nand n46402(x46402, x46328, x46286);
  nand n46404(x46404, x46402, x46403);
  nand n46405(x46405, x46328, x46288);
  nand n46407(x46407, x46333, x46291);
  nand n46409(x46409, x46407, x46408);
  nand n46410(x46410, x46333, x46293);
  nand n46412(x46412, x46338, x46296);
  nand n46414(x46414, x46412, x46413);
  nand n46415(x46415, x46338, x46298);
  nand n46417(x46417, x46343, x46301);
  nand n46419(x46419, x46417, x46418);
  nand n46420(x46420, x46343, x46303);
  nand n46422(x46422, x46348, x46306);
  nand n46424(x46424, x46422, x46423);
  nand n46425(x46425, x46348, x46308);
  nand n46427(x46427, x46353, x46311);
  nand n46429(x46429, x46427, x46428);
  nand n46430(x46430, x46353, x46313);
  nand n46438(x46438, x46386, x46010);
  nand n46440(x46440, x46438, x46439);
  nand n46441(x46441, x46391, x46036);
  nand n46443(x46443, x46441, x46442);
  nand n46444(x46444, x46396, x46136);
  nand n46446(x46446, x46444, x46445);
  nand n46447(x46447, x46401, x46139);
  nand n46449(x46449, x46447, x46448);
  nand n46450(x46450, x46406, x46254);
  nand n46452(x46452, x46450, x46451);
  nand n46453(x46453, x46411, x46257);
  nand n46455(x46455, x46453, x46454);
  nand n46456(x46456, x46416, x46260);
  nand n46458(x46458, x46456, x46457);
  nand n46459(x46459, x46421, x46263);
  nand n46461(x46461, x46459, x46460);
  nand n46462(x46462, x46426, x46360);
  nand n46464(x46464, x46462, x46463);
  nand n46465(x46465, x46431, x46363);
  nand n46467(x46467, x46465, x46466);
  nand n46468(x46468, x45884, x45878);
  nand n46469(x46469, x46468, x46035);
  nand n46471(x46471, x45889, x46036);
  nand n46472(x46472, x45888, x46133);
  nand n46473(x46473, x46472, x46471);
  nand n46475(x46475, x45894, x46136);
  nand n46476(x46476, x45893, x46250);
  nand n46477(x46477, x46476, x46475);
  nand n46479(x46479, x45899, x46139);
  nand n46480(x46480, x45898, x46251);
  nand n46481(x46481, x46480, x46479);
  nand n46483(x46483, x45904, x46254);
  nand n46484(x46484, x45903, x46354);
  nand n46485(x46485, x46484, x46483);
  nand n46487(x46487, x45909, x46257);
  nand n46488(x46488, x45908, x46355);
  nand n46489(x46489, x46488, x46487);
  nand n46491(x46491, x45914, x46260);
  nand n46492(x46492, x45913, x46356);
  nand n46493(x46493, x46492, x46491);
  nand n46495(x46495, x45919, x46263);
  nand n46496(x46496, x45918, x46357);
  nand n46497(x46497, x46496, x46495);
  nand n46499(x46499, x45924, x46360);
  nand n46501(x46501, x45923, x46500);
  nand n46502(x46502, x46501, x46499);
  nand n46504(x46504, x45929, x46363);
  nand n46506(x46506, x45928, x46505);
  nand n46507(x46507, x46506, x46504);
  nand n46509(x46509, x45934, x46366);
  nand n46510(x46510, x45933, x46432);
  nand n46511(x46511, x46510, x46509);
  nand n46513(x46513, x45939, x46369);
  nand n46514(x46514, x45938, x46433);
  nand n46515(x46515, x46514, x46513);
  nand n46517(x46517, x45944, x46372);
  nand n46518(x46518, x45943, x46434);
  nand n46519(x46519, x46518, x46517);
  nand n46521(x46521, x45949, x46375);
  nand n46522(x46522, x45948, x46435);
  nand n46523(x46523, x46522, x46521);
  nand n46525(x46525, x45954, x46378);
  nand n46526(x46526, x45953, x46436);
  nand n46527(x46527, x46526, x46525);
  nand n46529(x46529, x45959, x46381);
  nand n46530(x46530, x45958, x46437);
  nand n46531(x46531, x46530, x46529);
  nand n46533(x46533, x45964, x46440);
  nand n46535(x46535, x45963, x46534);
  nand n46536(x46536, x46535, x46533);
  nand n46538(x46538, x45969, x46443);
  nand n46540(x46540, x45968, x46539);
  nand n46541(x46541, x46540, x46538);
  nand n46543(x46543, x45974, x46446);
  nand n46545(x46545, x45973, x46544);
  nand n46546(x46546, x46545, x46543);
  nand n46548(x46548, x45979, x46449);
  nand n46550(x46550, x45978, x46549);
  nand n46551(x46551, x46550, x46548);
  nand n46553(x46553, x45984, x46452);
  nand n46555(x46555, x45983, x46554);
  nand n46556(x46556, x46555, x46553);
  nand n46558(x46558, x45989, x46455);
  nand n46560(x46560, x45988, x46559);
  nand n46561(x46561, x46560, x46558);
  nand n46563(x46563, x45994, x46458);
  nand n46565(x46565, x45993, x46564);
  nand n46566(x46566, x46565, x46563);
  nand n46568(x46568, x45999, x46461);
  nand n46570(x46570, x45998, x46569);
  nand n46571(x46571, x46570, x46568);
  nand n46573(x46573, x46004, x46464);
  nand n46575(x46575, x46003, x46574);
  nand n46576(x46576, x46575, x46573);
  nand n46578(x46578, x46009, x46467);
  nand n46580(x46580, x46008, x46579);
  nand n46581(x46581, x46580, x46578);
  nand n46583(x46583, x39047, x39041);
  nand n46585(x46585, x39053, x39047);
  nand n46587(x46587, x39059, x39053);
  nand n46589(x46589, x39065, x39059);
  nand n46591(x46591, x39071, x39065);
  nand n46593(x46593, x39077, x39071);
  nand n46595(x46595, x39083, x39077);
  nand n46597(x46597, x39089, x39083);
  nand n46599(x46599, x39095, x39089);
  nand n46601(x46601, x39101, x39095);
  nand n46603(x46603, x39107, x39101);
  nand n46605(x46605, x39113, x39107);
  nand n46607(x46607, x39119, x39113);
  nand n46609(x46609, x39125, x39119);
  nand n46611(x46611, x39131, x39125);
  nand n46613(x46613, x39137, x39131);
  nand n46615(x46615, x39143, x39137);
  nand n46617(x46617, x39149, x39143);
  nand n46619(x46619, x39155, x39149);
  nand n46621(x46621, x39161, x39155);
  nand n46623(x46623, x39167, x39161);
  nand n46625(x46625, x39173, x39167);
  nand n46627(x46627, x39179, x39173);
  nand n46629(x46629, x39185, x39179);
  nand n46631(x46631, x39191, x39185);
  nand n46633(x46633, x39197, x39191);
  nand n46635(x46635, x39203, x39197);
  nand n46637(x46637, x39209, x39203);
  nand n46639(x46639, x39215, x39209);
  nand n46641(x46641, x39221, x39215);
  nand n46643(x46643, x46586, x39041);
  nand n46644(x46644, x46588, x46584);
  nand n46646(x46646, x46590, x46586);
  nand n46648(x46648, x46592, x46588);
  nand n46650(x46650, x46594, x46590);
  nand n46652(x46652, x46596, x46592);
  nand n46654(x46654, x46598, x46594);
  nand n46656(x46656, x46600, x46596);
  nand n46658(x46658, x46602, x46598);
  nand n46660(x46660, x46604, x46600);
  nand n46662(x46662, x46606, x46602);
  nand n46664(x46664, x46608, x46604);
  nand n46666(x46666, x46610, x46606);
  nand n46668(x46668, x46612, x46608);
  nand n46670(x46670, x46614, x46610);
  nand n46672(x46672, x46616, x46612);
  nand n46674(x46674, x46618, x46614);
  nand n46676(x46676, x46620, x46616);
  nand n46678(x46678, x46622, x46618);
  nand n46680(x46680, x46624, x46620);
  nand n46682(x46682, x46626, x46622);
  nand n46684(x46684, x46628, x46624);
  nand n46686(x46686, x46630, x46626);
  nand n46688(x46688, x46632, x46628);
  nand n46690(x46690, x46634, x46630);
  nand n46692(x46692, x46636, x46632);
  nand n46694(x46694, x46638, x46634);
  nand n46696(x46696, x46640, x46636);
  nand n46698(x46698, x46642, x46638);
  nand n46700(x46700, x46647, x39041);
  nand n46701(x46701, x46649, x46584);
  nand n46702(x46702, x46651, x85212);
  nand n46703(x46703, x46653, x46645);
  nand n46705(x46705, x46655, x46647);
  nand n46707(x46707, x46657, x46649);
  nand n46709(x46709, x46659, x46651);
  nand n46711(x46711, x46661, x46653);
  nand n46713(x46713, x46663, x46655);
  nand n46715(x46715, x46665, x46657);
  nand n46717(x46717, x46667, x46659);
  nand n46719(x46719, x46669, x46661);
  nand n46721(x46721, x46671, x46663);
  nand n46723(x46723, x46673, x46665);
  nand n46725(x46725, x46675, x46667);
  nand n46727(x46727, x46677, x46669);
  nand n46729(x46729, x46679, x46671);
  nand n46731(x46731, x46681, x46673);
  nand n46733(x46733, x46683, x46675);
  nand n46735(x46735, x46685, x46677);
  nand n46737(x46737, x46687, x46679);
  nand n46739(x46739, x46689, x46681);
  nand n46741(x46741, x46691, x46683);
  nand n46743(x46743, x46693, x46685);
  nand n46745(x46745, x46695, x46687);
  nand n46747(x46747, x46697, x46689);
  nand n46749(x46749, x46699, x46691);
  nand n46751(x46751, x46706, x39041);
  nand n46752(x46752, x46708, x46584);
  nand n46753(x46753, x46710, x85212);
  nand n46754(x46754, x46712, x46645);
  nand n46755(x46755, x46714, x85213);
  nand n46756(x46756, x46716, x85214);
  nand n46757(x46757, x46718, x85215);
  nand n46758(x46758, x46720, x46704);
  nand n46759(x46759, x46722, x46706);
  nand n46761(x46761, x46724, x46708);
  nand n46763(x46763, x46726, x46710);
  nand n46765(x46765, x46728, x46712);
  nand n46767(x46767, x46730, x46714);
  nand n46769(x46769, x46732, x46716);
  nand n46771(x46771, x46734, x46718);
  nand n46773(x46773, x46736, x46720);
  nand n46775(x46775, x46738, x46722);
  nand n46777(x46777, x46740, x46724);
  nand n46779(x46779, x46742, x46726);
  nand n46781(x46781, x46744, x46728);
  nand n46783(x46783, x46746, x46730);
  nand n46785(x46785, x46748, x46732);
  nand n46787(x46787, x46750, x46734);
  nand n46789(x46789, x46760, x39041);
  nand n46790(x46790, x46762, x46584);
  nand n46791(x46791, x46764, x85212);
  nand n46792(x46792, x46766, x46645);
  nand n46793(x46793, x46768, x85213);
  nand n46794(x46794, x46770, x85214);
  nand n46795(x46795, x46772, x85215);
  nand n46796(x46796, x46774, x46704);
  nand n46797(x46797, x46776, x85216);
  nand n46798(x46798, x46778, x85217);
  nand n46799(x46799, x46780, x85218);
  nand n46800(x46800, x46782, x85219);
  nand n46801(x46801, x46784, x85220);
  nand n46802(x46802, x46786, x85221);
  nand n46803(x46803, x46788, x85222);
  nand n46804(x46804, x73032, x73027);
  nand n46805(x46805, x46804, x46583);
  nand n46807(x46807, x39053, x46584);
  nand n46808(x46808, x73037, x46583);
  nand n46809(x46809, x46808, x46807);
  nand n46811(x46811, x39059, x85212);
  nand n46812(x46812, x73042, x46643);
  nand n46813(x46813, x46812, x46811);
  nand n46815(x46815, x39065, x46645);
  nand n46816(x46816, x73047, x46644);
  nand n46817(x46817, x46816, x46815);
  nand n46819(x46819, x39071, x85213);
  nand n46820(x46820, x73052, x46700);
  nand n46821(x46821, x46820, x46819);
  nand n46823(x46823, x39077, x85214);
  nand n46824(x46824, x73057, x46701);
  nand n46825(x46825, x46824, x46823);
  nand n46827(x46827, x39083, x85215);
  nand n46828(x46828, x73062, x46702);
  nand n46829(x46829, x46828, x46827);
  nand n46831(x46831, x39089, x46704);
  nand n46832(x46832, x73067, x46703);
  nand n46833(x46833, x46832, x46831);
  nand n46835(x46835, x39095, x85216);
  nand n46836(x46836, x73072, x46751);
  nand n46837(x46837, x46836, x46835);
  nand n46839(x46839, x39101, x85217);
  nand n46840(x46840, x73077, x46752);
  nand n46841(x46841, x46840, x46839);
  nand n46843(x46843, x39107, x85218);
  nand n46844(x46844, x73082, x46753);
  nand n46845(x46845, x46844, x46843);
  nand n46847(x46847, x39113, x85219);
  nand n46848(x46848, x73087, x46754);
  nand n46849(x46849, x46848, x46847);
  nand n46851(x46851, x39119, x85220);
  nand n46852(x46852, x73092, x46755);
  nand n46853(x46853, x46852, x46851);
  nand n46855(x46855, x39125, x85221);
  nand n46856(x46856, x73097, x46756);
  nand n46857(x46857, x46856, x46855);
  nand n46859(x46859, x39131, x85222);
  nand n46860(x46860, x73102, x46757);
  nand n46861(x46861, x46860, x46859);
  nand n46863(x46863, x39137, x85223);
  nand n46864(x46864, x73107, x46758);
  nand n46865(x46865, x46864, x46863);
  nand n46867(x46867, x39143, x85224);
  nand n46868(x46868, x73112, x46789);
  nand n46869(x46869, x46868, x46867);
  nand n46871(x46871, x39149, x85225);
  nand n46872(x46872, x73117, x46790);
  nand n46873(x46873, x46872, x46871);
  nand n46875(x46875, x39155, x85226);
  nand n46876(x46876, x73122, x46791);
  nand n46877(x46877, x46876, x46875);
  nand n46879(x46879, x39161, x85227);
  nand n46880(x46880, x73127, x46792);
  nand n46881(x46881, x46880, x46879);
  nand n46883(x46883, x39167, x85228);
  nand n46884(x46884, x73132, x46793);
  nand n46885(x46885, x46884, x46883);
  nand n46887(x46887, x39173, x85229);
  nand n46888(x46888, x73137, x46794);
  nand n46889(x46889, x46888, x46887);
  nand n46891(x46891, x39179, x85230);
  nand n46892(x46892, x73142, x46795);
  nand n46893(x46893, x46892, x46891);
  nand n46895(x46895, x39185, x85231);
  nand n46896(x46896, x73147, x46796);
  nand n46897(x46897, x46896, x46895);
  nand n46899(x46899, x39191, x85232);
  nand n46900(x46900, x73152, x46797);
  nand n46901(x46901, x46900, x46899);
  nand n46903(x46903, x39197, x85233);
  nand n46904(x46904, x73157, x46798);
  nand n46905(x46905, x46904, x46903);
  nand n46907(x46907, x39203, x85234);
  nand n46908(x46908, x73162, x46799);
  nand n46909(x46909, x46908, x46907);
  nand n46911(x46911, x39209, x85235);
  nand n46912(x46912, x73167, x46800);
  nand n46913(x46913, x46912, x46911);
  nand n46915(x46915, x39215, x85236);
  nand n46916(x46916, x73172, x46801);
  nand n46917(x46917, x46916, x46915);
  nand n46919(x46919, x39221, x85237);
  nand n46920(x46920, x73177, x46802);
  nand n46921(x46921, x46920, x46919);
  nand n46923(x46923, x39227, x85238);
  nand n46924(x46924, x73182, x46803);
  nand n46925(x46925, x46924, x46923);
  nand n46928(x46928, x73107, x38880);
  nand n46930(x46930, x73112, x38882);
  nand n46932(x46932, x73117, x38884);
  nand n46934(x46934, x73122, x38886);
  nand n46936(x46936, x73127, x38888);
  nand n46938(x46938, x73132, x38890);
  nand n46940(x46940, x73137, x38892);
  nand n46942(x46942, x73142, x38894);
  nand n46944(x46944, x73147, x38896);
  nand n46946(x46946, x73152, x38898);
  nand n46948(x46948, x73157, x38900);
  nand n46950(x46950, x73162, x38902);
  nand n46952(x46952, x73167, x38904);
  nand n46954(x46954, x73172, x38906);
  nand n46956(x46956, x73177, x38908);
  nand n46958(x46958, x73182, x38910);
  nand n46960(x46960, x39041, x38911);
  nand n46961(x46961, x39047, x38912);
  nand n46962(x46962, x39053, x38913);
  nand n46963(x46963, x39059, x38914);
  nand n46964(x46964, x39065, x38915);
  nand n46965(x46965, x39071, x38916);
  nand n46966(x46966, x39077, x38917);
  nand n46967(x46967, x39083, x38918);
  nand n46968(x46968, x39089, x38919);
  nand n46969(x46969, x39095, x38920);
  nand n46970(x46970, x39101, x38921);
  nand n46971(x46971, x39107, x38922);
  nand n46972(x46972, x39113, x38923);
  nand n46973(x46973, x39119, x38924);
  nand n46974(x46974, x39125, x38925);
  nand n46975(x46975, x39131, x38926);
  nand n46976(x46976, x39137, x38927);
  nand n46977(x46977, x39143, x38928);
  nand n46978(x46978, x39149, x38929);
  nand n46979(x46979, x39155, x38930);
  nand n46980(x46980, x39161, x38931);
  nand n46981(x46981, x39167, x38932);
  nand n46982(x46982, x39173, x38933);
  nand n46983(x46983, x39179, x38934);
  nand n46984(x46984, x39185, x38935);
  nand n46985(x46985, x39191, x38936);
  nand n46986(x46986, x39197, x38937);
  nand n46987(x46987, x39203, x38938);
  nand n46988(x46988, x39209, x38939);
  nand n46989(x46989, x39215, x38940);
  nand n46990(x46990, x39221, x38941);
  nand n46991(x46991, x39227, x38942);
  nand n46992(x46992, x46960, x39971);
  nand n46994(x46994, x46961, x39978);
  nand n46996(x46996, x46962, x39993);
  nand n46998(x46998, x46963, x40017);
  nand n47000(x47000, x46964, x40048);
  nand n47002(x47002, x46965, x40087);
  nand n47004(x47004, x46966, x40135);
  nand n47006(x47006, x46967, x40190);
  nand n47008(x47008, x46968, x40253);
  nand n47010(x47010, x46969, x40325);
  nand n47012(x47012, x46970, x40404);
  nand n47014(x47014, x46971, x40491);
  nand n47016(x47016, x46972, x40587);
  nand n47018(x47018, x46973, x40690);
  nand n47020(x47020, x46974, x40801);
  nand n47022(x47022, x46975, x40921);
  nand n47024(x47024, x46976, x46928);
  nand n47026(x47026, x46977, x46930);
  nand n47028(x47028, x46978, x46932);
  nand n47030(x47030, x46979, x46934);
  nand n47032(x47032, x46980, x46936);
  nand n47034(x47034, x46981, x46938);
  nand n47036(x47036, x46982, x46940);
  nand n47038(x47038, x46983, x46942);
  nand n47040(x47040, x46984, x46944);
  nand n47042(x47042, x46985, x46946);
  nand n47044(x47044, x46986, x46948);
  nand n47046(x47046, x46987, x46950);
  nand n47048(x47048, x46988, x46952);
  nand n47050(x47050, x46989, x46954);
  nand n47052(x47052, x46990, x46956);
  nand n47054(x47054, x46991, x46958);
  nand n47056(x47056, x38911, x73027);
  nand n47057(x47057, x38911, x73032);
  nand n47058(x47058, x47057, x39971);
  nand n47059(x47059, x38911, x73037);
  nand n47060(x47060, x47059, x39972);
  nand n47061(x47061, x38911, x73042);
  nand n47062(x47062, x47061, x39976);
  nand n47063(x47063, x38911, x73047);
  nand n47064(x47064, x47063, x39982);
  nand n47065(x47065, x38911, x73052);
  nand n47066(x47066, x47065, x39989);
  nand n47067(x47067, x38911, x73057);
  nand n47068(x47068, x47067, x39999);
  nand n47069(x47069, x38911, x73062);
  nand n47070(x47070, x47069, x40011);
  nand n47071(x47071, x38911, x73067);
  nand n47072(x47072, x47071, x40024);
  nand n47073(x47073, x38911, x73072);
  nand n47074(x47074, x47073, x40040);
  nand n47075(x47075, x38911, x73077);
  nand n47076(x47076, x47075, x40058);
  nand n47077(x47077, x38911, x73082);
  nand n47078(x47078, x47077, x40077);
  nand n47079(x47079, x38911, x73087);
  nand n47080(x47080, x47079, x40099);
  nand n47081(x47081, x38911, x73092);
  nand n47082(x47082, x47081, x40123);
  nand n47083(x47083, x38911, x73097);
  nand n47084(x47084, x47083, x40148);
  nand n47085(x47085, x38911, x73102);
  nand n47086(x47086, x47085, x40176);
  nand n47087(x47087, x38911, x73107);
  nand n47088(x47088, x47087, x40206);
  nand n47089(x47089, x38911, x73112);
  nand n47090(x47090, x47089, x40237);
  nand n47091(x47091, x38911, x73117);
  nand n47092(x47092, x47091, x40271);
  nand n47093(x47093, x38911, x73122);
  nand n47094(x47094, x47093, x40307);
  nand n47095(x47095, x38911, x73127);
  nand n47096(x47096, x47095, x40344);
  nand n47097(x47097, x38911, x73132);
  nand n47098(x47098, x47097, x40384);
  nand n47099(x47099, x38911, x73137);
  nand n47100(x47100, x47099, x40426);
  nand n47101(x47101, x38911, x73142);
  nand n47102(x47102, x47101, x40469);
  nand n47103(x47103, x38911, x73147);
  nand n47104(x47104, x47103, x40515);
  nand n47105(x47105, x38911, x73152);
  nand n47106(x47106, x47105, x40563);
  nand n47107(x47107, x38911, x73157);
  nand n47108(x47108, x47107, x40612);
  nand n47109(x47109, x38911, x73162);
  nand n47110(x47110, x47109, x40664);
  nand n47111(x47111, x38911, x73167);
  nand n47112(x47112, x47111, x40718);
  nand n47113(x47113, x38911, x73172);
  nand n47114(x47114, x47113, x40773);
  nand n47115(x47115, x38911, x73177);
  nand n47116(x47116, x47115, x40831);
  nand n47117(x47117, x38911, x73182);
  nand n47118(x47118, x47117, x40891);
  nand n47119(x47119, x38912, x85239);
  nand n47120(x47120, x38912, x47058);
  nand n47121(x47121, x38850, x85239);
  nand n47122(x47122, x38912, x47060);
  nand n47123(x47123, x47122, x47121);
  nand n47124(x47124, x38850, x47058);
  nand n47125(x47125, x38912, x47062);
  nand n47126(x47126, x47125, x47124);
  nand n47127(x47127, x38850, x47060);
  nand n47128(x47128, x38912, x47064);
  nand n47129(x47129, x47128, x47127);
  nand n47130(x47130, x38850, x47062);
  nand n47131(x47131, x38912, x47066);
  nand n47132(x47132, x47131, x47130);
  nand n47133(x47133, x38850, x47064);
  nand n47134(x47134, x38912, x47068);
  nand n47135(x47135, x47134, x47133);
  nand n47136(x47136, x38850, x47066);
  nand n47137(x47137, x38912, x47070);
  nand n47138(x47138, x47137, x47136);
  nand n47139(x47139, x38850, x47068);
  nand n47140(x47140, x38912, x47072);
  nand n47141(x47141, x47140, x47139);
  nand n47142(x47142, x38850, x47070);
  nand n47143(x47143, x38912, x47074);
  nand n47144(x47144, x47143, x47142);
  nand n47145(x47145, x38850, x47072);
  nand n47146(x47146, x38912, x47076);
  nand n47147(x47147, x47146, x47145);
  nand n47148(x47148, x38850, x47074);
  nand n47149(x47149, x38912, x47078);
  nand n47150(x47150, x47149, x47148);
  nand n47151(x47151, x38850, x47076);
  nand n47152(x47152, x38912, x47080);
  nand n47153(x47153, x47152, x47151);
  nand n47154(x47154, x38850, x47078);
  nand n47155(x47155, x38912, x47082);
  nand n47156(x47156, x47155, x47154);
  nand n47157(x47157, x38850, x47080);
  nand n47158(x47158, x38912, x47084);
  nand n47159(x47159, x47158, x47157);
  nand n47160(x47160, x38850, x47082);
  nand n47161(x47161, x38912, x47086);
  nand n47162(x47162, x47161, x47160);
  nand n47163(x47163, x38850, x47084);
  nand n47164(x47164, x38912, x47088);
  nand n47165(x47165, x47164, x47163);
  nand n47166(x47166, x38850, x47086);
  nand n47167(x47167, x38912, x47090);
  nand n47168(x47168, x47167, x47166);
  nand n47169(x47169, x38850, x47088);
  nand n47170(x47170, x38912, x47092);
  nand n47171(x47171, x47170, x47169);
  nand n47172(x47172, x38850, x47090);
  nand n47173(x47173, x38912, x47094);
  nand n47174(x47174, x47173, x47172);
  nand n47175(x47175, x38850, x47092);
  nand n47176(x47176, x38912, x47096);
  nand n47177(x47177, x47176, x47175);
  nand n47178(x47178, x38850, x47094);
  nand n47179(x47179, x38912, x47098);
  nand n47180(x47180, x47179, x47178);
  nand n47181(x47181, x38850, x47096);
  nand n47182(x47182, x38912, x47100);
  nand n47183(x47183, x47182, x47181);
  nand n47184(x47184, x38850, x47098);
  nand n47185(x47185, x38912, x47102);
  nand n47186(x47186, x47185, x47184);
  nand n47187(x47187, x38850, x47100);
  nand n47188(x47188, x38912, x47104);
  nand n47189(x47189, x47188, x47187);
  nand n47190(x47190, x38850, x47102);
  nand n47191(x47191, x38912, x47106);
  nand n47192(x47192, x47191, x47190);
  nand n47193(x47193, x38850, x47104);
  nand n47194(x47194, x38912, x47108);
  nand n47195(x47195, x47194, x47193);
  nand n47196(x47196, x38850, x47106);
  nand n47197(x47197, x38912, x47110);
  nand n47198(x47198, x47197, x47196);
  nand n47199(x47199, x38850, x47108);
  nand n47200(x47200, x38912, x47112);
  nand n47201(x47201, x47200, x47199);
  nand n47202(x47202, x38850, x47110);
  nand n47203(x47203, x38912, x47114);
  nand n47204(x47204, x47203, x47202);
  nand n47205(x47205, x38850, x47112);
  nand n47206(x47206, x38912, x47116);
  nand n47207(x47207, x47206, x47205);
  nand n47208(x47208, x38850, x47114);
  nand n47209(x47209, x38912, x47118);
  nand n47210(x47210, x47209, x47208);
  nand n47211(x47211, x38913, x85240);
  nand n47212(x47212, x38913, x85241);
  nand n47213(x47213, x38913, x47123);
  nand n47214(x47214, x38913, x47126);
  nand n47215(x47215, x38852, x85240);
  nand n47216(x47216, x38913, x47129);
  nand n47217(x47217, x47216, x47215);
  nand n47218(x47218, x38852, x85241);
  nand n47219(x47219, x38913, x47132);
  nand n47220(x47220, x47219, x47218);
  nand n47221(x47221, x38852, x47123);
  nand n47222(x47222, x38913, x47135);
  nand n47223(x47223, x47222, x47221);
  nand n47224(x47224, x38852, x47126);
  nand n47225(x47225, x38913, x47138);
  nand n47226(x47226, x47225, x47224);
  nand n47227(x47227, x38852, x47129);
  nand n47228(x47228, x38913, x47141);
  nand n47229(x47229, x47228, x47227);
  nand n47230(x47230, x38852, x47132);
  nand n47231(x47231, x38913, x47144);
  nand n47232(x47232, x47231, x47230);
  nand n47233(x47233, x38852, x47135);
  nand n47234(x47234, x38913, x47147);
  nand n47235(x47235, x47234, x47233);
  nand n47236(x47236, x38852, x47138);
  nand n47237(x47237, x38913, x47150);
  nand n47238(x47238, x47237, x47236);
  nand n47239(x47239, x38852, x47141);
  nand n47240(x47240, x38913, x47153);
  nand n47241(x47241, x47240, x47239);
  nand n47242(x47242, x38852, x47144);
  nand n47243(x47243, x38913, x47156);
  nand n47244(x47244, x47243, x47242);
  nand n47245(x47245, x38852, x47147);
  nand n47246(x47246, x38913, x47159);
  nand n47247(x47247, x47246, x47245);
  nand n47248(x47248, x38852, x47150);
  nand n47249(x47249, x38913, x47162);
  nand n47250(x47250, x47249, x47248);
  nand n47251(x47251, x38852, x47153);
  nand n47252(x47252, x38913, x47165);
  nand n47253(x47253, x47252, x47251);
  nand n47254(x47254, x38852, x47156);
  nand n47255(x47255, x38913, x47168);
  nand n47256(x47256, x47255, x47254);
  nand n47257(x47257, x38852, x47159);
  nand n47258(x47258, x38913, x47171);
  nand n47259(x47259, x47258, x47257);
  nand n47260(x47260, x38852, x47162);
  nand n47261(x47261, x38913, x47174);
  nand n47262(x47262, x47261, x47260);
  nand n47263(x47263, x38852, x47165);
  nand n47264(x47264, x38913, x47177);
  nand n47265(x47265, x47264, x47263);
  nand n47266(x47266, x38852, x47168);
  nand n47267(x47267, x38913, x47180);
  nand n47268(x47268, x47267, x47266);
  nand n47269(x47269, x38852, x47171);
  nand n47270(x47270, x38913, x47183);
  nand n47271(x47271, x47270, x47269);
  nand n47272(x47272, x38852, x47174);
  nand n47273(x47273, x38913, x47186);
  nand n47274(x47274, x47273, x47272);
  nand n47275(x47275, x38852, x47177);
  nand n47276(x47276, x38913, x47189);
  nand n47277(x47277, x47276, x47275);
  nand n47278(x47278, x38852, x47180);
  nand n47279(x47279, x38913, x47192);
  nand n47280(x47280, x47279, x47278);
  nand n47281(x47281, x38852, x47183);
  nand n47282(x47282, x38913, x47195);
  nand n47283(x47283, x47282, x47281);
  nand n47284(x47284, x38852, x47186);
  nand n47285(x47285, x38913, x47198);
  nand n47286(x47286, x47285, x47284);
  nand n47287(x47287, x38852, x47189);
  nand n47288(x47288, x38913, x47201);
  nand n47289(x47289, x47288, x47287);
  nand n47290(x47290, x38852, x47192);
  nand n47291(x47291, x38913, x47204);
  nand n47292(x47292, x47291, x47290);
  nand n47293(x47293, x38852, x47195);
  nand n47294(x47294, x38913, x47207);
  nand n47295(x47295, x47294, x47293);
  nand n47296(x47296, x38852, x47198);
  nand n47297(x47297, x38913, x47210);
  nand n47298(x47298, x47297, x47296);
  nand n47299(x47299, x38914, x85242);
  nand n47300(x47300, x38914, x85243);
  nand n47301(x47301, x38914, x85244);
  nand n47302(x47302, x38914, x85245);
  nand n47303(x47303, x38914, x47217);
  nand n47304(x47304, x38914, x47220);
  nand n47305(x47305, x38914, x47223);
  nand n47306(x47306, x38914, x47226);
  nand n47307(x47307, x38854, x85242);
  nand n47308(x47308, x38914, x47229);
  nand n47309(x47309, x47308, x47307);
  nand n47310(x47310, x38854, x85243);
  nand n47311(x47311, x38914, x47232);
  nand n47312(x47312, x47311, x47310);
  nand n47313(x47313, x38854, x85244);
  nand n47314(x47314, x38914, x47235);
  nand n47315(x47315, x47314, x47313);
  nand n47316(x47316, x38854, x85245);
  nand n47317(x47317, x38914, x47238);
  nand n47318(x47318, x47317, x47316);
  nand n47319(x47319, x38854, x47217);
  nand n47320(x47320, x38914, x47241);
  nand n47321(x47321, x47320, x47319);
  nand n47322(x47322, x38854, x47220);
  nand n47323(x47323, x38914, x47244);
  nand n47324(x47324, x47323, x47322);
  nand n47325(x47325, x38854, x47223);
  nand n47326(x47326, x38914, x47247);
  nand n47327(x47327, x47326, x47325);
  nand n47328(x47328, x38854, x47226);
  nand n47329(x47329, x38914, x47250);
  nand n47330(x47330, x47329, x47328);
  nand n47331(x47331, x38854, x47229);
  nand n47332(x47332, x38914, x47253);
  nand n47333(x47333, x47332, x47331);
  nand n47334(x47334, x38854, x47232);
  nand n47335(x47335, x38914, x47256);
  nand n47336(x47336, x47335, x47334);
  nand n47337(x47337, x38854, x47235);
  nand n47338(x47338, x38914, x47259);
  nand n47339(x47339, x47338, x47337);
  nand n47340(x47340, x38854, x47238);
  nand n47341(x47341, x38914, x47262);
  nand n47342(x47342, x47341, x47340);
  nand n47343(x47343, x38854, x47241);
  nand n47344(x47344, x38914, x47265);
  nand n47345(x47345, x47344, x47343);
  nand n47346(x47346, x38854, x47244);
  nand n47347(x47347, x38914, x47268);
  nand n47348(x47348, x47347, x47346);
  nand n47349(x47349, x38854, x47247);
  nand n47350(x47350, x38914, x47271);
  nand n47351(x47351, x47350, x47349);
  nand n47352(x47352, x38854, x47250);
  nand n47353(x47353, x38914, x47274);
  nand n47354(x47354, x47353, x47352);
  nand n47355(x47355, x38854, x47253);
  nand n47356(x47356, x38914, x47277);
  nand n47357(x47357, x47356, x47355);
  nand n47358(x47358, x38854, x47256);
  nand n47359(x47359, x38914, x47280);
  nand n47360(x47360, x47359, x47358);
  nand n47361(x47361, x38854, x47259);
  nand n47362(x47362, x38914, x47283);
  nand n47363(x47363, x47362, x47361);
  nand n47364(x47364, x38854, x47262);
  nand n47365(x47365, x38914, x47286);
  nand n47366(x47366, x47365, x47364);
  nand n47367(x47367, x38854, x47265);
  nand n47368(x47368, x38914, x47289);
  nand n47369(x47369, x47368, x47367);
  nand n47370(x47370, x38854, x47268);
  nand n47371(x47371, x38914, x47292);
  nand n47372(x47372, x47371, x47370);
  nand n47373(x47373, x38854, x47271);
  nand n47374(x47374, x38914, x47295);
  nand n47375(x47375, x47374, x47373);
  nand n47376(x47376, x38854, x47274);
  nand n47377(x47377, x38914, x47298);
  nand n47378(x47378, x47377, x47376);
  nand n47379(x47379, x38915, x85246);
  nand n47380(x47380, x38915, x85247);
  nand n47381(x47381, x38915, x85248);
  nand n47382(x47382, x38915, x85249);
  nand n47383(x47383, x38915, x85250);
  nand n47384(x47384, x38915, x85251);
  nand n47385(x47385, x38915, x85252);
  nand n47386(x47386, x38915, x85253);
  nand n47387(x47387, x38915, x47309);
  nand n47388(x47388, x38915, x47312);
  nand n47389(x47389, x38915, x47315);
  nand n47390(x47390, x38915, x47318);
  nand n47391(x47391, x38915, x47321);
  nand n47392(x47392, x38915, x47324);
  nand n47393(x47393, x38915, x47327);
  nand n47394(x47394, x38915, x47330);
  nand n47395(x47395, x38856, x85246);
  nand n47396(x47396, x38915, x47333);
  nand n47397(x47397, x47396, x47395);
  nand n47398(x47398, x38856, x85247);
  nand n47399(x47399, x38915, x47336);
  nand n47400(x47400, x47399, x47398);
  nand n47401(x47401, x38856, x85248);
  nand n47402(x47402, x38915, x47339);
  nand n47403(x47403, x47402, x47401);
  nand n47404(x47404, x38856, x85249);
  nand n47405(x47405, x38915, x47342);
  nand n47406(x47406, x47405, x47404);
  nand n47407(x47407, x38856, x85250);
  nand n47408(x47408, x38915, x47345);
  nand n47409(x47409, x47408, x47407);
  nand n47410(x47410, x38856, x85251);
  nand n47411(x47411, x38915, x47348);
  nand n47412(x47412, x47411, x47410);
  nand n47413(x47413, x38856, x85252);
  nand n47414(x47414, x38915, x47351);
  nand n47415(x47415, x47414, x47413);
  nand n47416(x47416, x38856, x85253);
  nand n47417(x47417, x38915, x47354);
  nand n47418(x47418, x47417, x47416);
  nand n47419(x47419, x38856, x47309);
  nand n47420(x47420, x38915, x47357);
  nand n47421(x47421, x47420, x47419);
  nand n47422(x47422, x38856, x47312);
  nand n47423(x47423, x38915, x47360);
  nand n47424(x47424, x47423, x47422);
  nand n47425(x47425, x38856, x47315);
  nand n47426(x47426, x38915, x47363);
  nand n47427(x47427, x47426, x47425);
  nand n47428(x47428, x38856, x47318);
  nand n47429(x47429, x38915, x47366);
  nand n47430(x47430, x47429, x47428);
  nand n47431(x47431, x38856, x47321);
  nand n47432(x47432, x38915, x47369);
  nand n47433(x47433, x47432, x47431);
  nand n47434(x47434, x38856, x47324);
  nand n47435(x47435, x38915, x47372);
  nand n47436(x47436, x47435, x47434);
  nand n47437(x47437, x38856, x47327);
  nand n47438(x47438, x38915, x47375);
  nand n47439(x47439, x47438, x47437);
  nand n47440(x47440, x38856, x47330);
  nand n47441(x47441, x38915, x47378);
  nand n47442(x47442, x47441, x47440);
  nand n47443(x47443, x47056, x39972);
  nand n47444(x47444, x47057, x39976);
  nand n47445(x47445, x47059, x39982);
  nand n47446(x47446, x47061, x39989);
  nand n47447(x47447, x47063, x39999);
  nand n47448(x47448, x47065, x40011);
  nand n47449(x47449, x47067, x40024);
  nand n47450(x47450, x47069, x40040);
  nand n47451(x47451, x47071, x40058);
  nand n47452(x47452, x47073, x40077);
  nand n47453(x47453, x47075, x40099);
  nand n47454(x47454, x47077, x40123);
  nand n47455(x47455, x47079, x40148);
  nand n47456(x47456, x47081, x40176);
  nand n47457(x47457, x47083, x40206);
  nand n47458(x47458, x47085, x40237);
  nand n47459(x47459, x47087, x40271);
  nand n47460(x47460, x47089, x40307);
  nand n47461(x47461, x47091, x40344);
  nand n47462(x47462, x47093, x40384);
  nand n47463(x47463, x47095, x40426);
  nand n47464(x47464, x47097, x40469);
  nand n47465(x47465, x47099, x40515);
  nand n47466(x47466, x47101, x40563);
  nand n47467(x47467, x47103, x40612);
  nand n47468(x47468, x47105, x40664);
  nand n47469(x47469, x47107, x40718);
  nand n47470(x47470, x47109, x40773);
  nand n47471(x47471, x47111, x40831);
  nand n47472(x47472, x47113, x40891);
  nand n47473(x47473, x47115, x40952);
  nand n47474(x47474, x38850, x47445);
  nand n47475(x47475, x38912, x47443);
  nand n47476(x47476, x47475, x47474);
  nand n47477(x47477, x38850, x47446);
  nand n47478(x47478, x38912, x47444);
  nand n47479(x47479, x47478, x47477);
  nand n47480(x47480, x38850, x47447);
  nand n47481(x47481, x38912, x47445);
  nand n47482(x47482, x47481, x47480);
  nand n47483(x47483, x38850, x47448);
  nand n47484(x47484, x38912, x47446);
  nand n47485(x47485, x47484, x47483);
  nand n47486(x47486, x38850, x47449);
  nand n47487(x47487, x38912, x47447);
  nand n47488(x47488, x47487, x47486);
  nand n47489(x47489, x38850, x47450);
  nand n47490(x47490, x38912, x47448);
  nand n47491(x47491, x47490, x47489);
  nand n47492(x47492, x38850, x47451);
  nand n47493(x47493, x38912, x47449);
  nand n47494(x47494, x47493, x47492);
  nand n47495(x47495, x38850, x47452);
  nand n47496(x47496, x38912, x47450);
  nand n47497(x47497, x47496, x47495);
  nand n47498(x47498, x38850, x47453);
  nand n47499(x47499, x38912, x47451);
  nand n47500(x47500, x47499, x47498);
  nand n47501(x47501, x38850, x47454);
  nand n47502(x47502, x38912, x47452);
  nand n47503(x47503, x47502, x47501);
  nand n47504(x47504, x38850, x47455);
  nand n47505(x47505, x38912, x47453);
  nand n47506(x47506, x47505, x47504);
  nand n47507(x47507, x38850, x47456);
  nand n47508(x47508, x38912, x47454);
  nand n47509(x47509, x47508, x47507);
  nand n47510(x47510, x38850, x47457);
  nand n47511(x47511, x38912, x47455);
  nand n47512(x47512, x47511, x47510);
  nand n47513(x47513, x38850, x47458);
  nand n47514(x47514, x38912, x47456);
  nand n47515(x47515, x47514, x47513);
  nand n47516(x47516, x38850, x47459);
  nand n47517(x47517, x38912, x47457);
  nand n47518(x47518, x47517, x47516);
  nand n47519(x47519, x38850, x47460);
  nand n47520(x47520, x38912, x47458);
  nand n47521(x47521, x47520, x47519);
  nand n47522(x47522, x38850, x47461);
  nand n47523(x47523, x38912, x47459);
  nand n47524(x47524, x47523, x47522);
  nand n47525(x47525, x38850, x47462);
  nand n47526(x47526, x38912, x47460);
  nand n47527(x47527, x47526, x47525);
  nand n47528(x47528, x38850, x47463);
  nand n47529(x47529, x38912, x47461);
  nand n47530(x47530, x47529, x47528);
  nand n47531(x47531, x38850, x47464);
  nand n47532(x47532, x38912, x47462);
  nand n47533(x47533, x47532, x47531);
  nand n47534(x47534, x38850, x47465);
  nand n47535(x47535, x38912, x47463);
  nand n47536(x47536, x47535, x47534);
  nand n47537(x47537, x38850, x47466);
  nand n47538(x47538, x38912, x47464);
  nand n47539(x47539, x47538, x47537);
  nand n47540(x47540, x38850, x47467);
  nand n47541(x47541, x38912, x47465);
  nand n47542(x47542, x47541, x47540);
  nand n47543(x47543, x38850, x47468);
  nand n47544(x47544, x38912, x47466);
  nand n47545(x47545, x47544, x47543);
  nand n47546(x47546, x38850, x47469);
  nand n47547(x47547, x38912, x47467);
  nand n47548(x47548, x47547, x47546);
  nand n47549(x47549, x38850, x47470);
  nand n47550(x47550, x38912, x47468);
  nand n47551(x47551, x47550, x47549);
  nand n47552(x47552, x38850, x47471);
  nand n47553(x47553, x38912, x47469);
  nand n47554(x47554, x47553, x47552);
  nand n47555(x47555, x38850, x47472);
  nand n47556(x47556, x38912, x47470);
  nand n47557(x47557, x47556, x47555);
  nand n47558(x47558, x38850, x47473);
  nand n47559(x47559, x38912, x47471);
  nand n47560(x47560, x47559, x47558);
  nand n47561(x47561, x38850, x85270);
  nand n47562(x47562, x38912, x47472);
  nand n47563(x47563, x47562, x47561);
  nand n47564(x47564, x38912, x47473);
  nand n47565(x47565, x38912, x85270);
  nand n47566(x47566, x38852, x47488);
  nand n47567(x47567, x38913, x47476);
  nand n47568(x47568, x47567, x47566);
  nand n47569(x47569, x38852, x47491);
  nand n47570(x47570, x38913, x47479);
  nand n47571(x47571, x47570, x47569);
  nand n47572(x47572, x38852, x47494);
  nand n47573(x47573, x38913, x47482);
  nand n47574(x47574, x47573, x47572);
  nand n47575(x47575, x38852, x47497);
  nand n47576(x47576, x38913, x47485);
  nand n47577(x47577, x47576, x47575);
  nand n47578(x47578, x38852, x47500);
  nand n47579(x47579, x38913, x47488);
  nand n47580(x47580, x47579, x47578);
  nand n47581(x47581, x38852, x47503);
  nand n47582(x47582, x38913, x47491);
  nand n47583(x47583, x47582, x47581);
  nand n47584(x47584, x38852, x47506);
  nand n47585(x47585, x38913, x47494);
  nand n47586(x47586, x47585, x47584);
  nand n47587(x47587, x38852, x47509);
  nand n47588(x47588, x38913, x47497);
  nand n47589(x47589, x47588, x47587);
  nand n47590(x47590, x38852, x47512);
  nand n47591(x47591, x38913, x47500);
  nand n47592(x47592, x47591, x47590);
  nand n47593(x47593, x38852, x47515);
  nand n47594(x47594, x38913, x47503);
  nand n47595(x47595, x47594, x47593);
  nand n47596(x47596, x38852, x47518);
  nand n47597(x47597, x38913, x47506);
  nand n47598(x47598, x47597, x47596);
  nand n47599(x47599, x38852, x47521);
  nand n47600(x47600, x38913, x47509);
  nand n47601(x47601, x47600, x47599);
  nand n47602(x47602, x38852, x47524);
  nand n47603(x47603, x38913, x47512);
  nand n47604(x47604, x47603, x47602);
  nand n47605(x47605, x38852, x47527);
  nand n47606(x47606, x38913, x47515);
  nand n47607(x47607, x47606, x47605);
  nand n47608(x47608, x38852, x47530);
  nand n47609(x47609, x38913, x47518);
  nand n47610(x47610, x47609, x47608);
  nand n47611(x47611, x38852, x47533);
  nand n47612(x47612, x38913, x47521);
  nand n47613(x47613, x47612, x47611);
  nand n47614(x47614, x38852, x47536);
  nand n47615(x47615, x38913, x47524);
  nand n47616(x47616, x47615, x47614);
  nand n47617(x47617, x38852, x47539);
  nand n47618(x47618, x38913, x47527);
  nand n47619(x47619, x47618, x47617);
  nand n47620(x47620, x38852, x47542);
  nand n47621(x47621, x38913, x47530);
  nand n47622(x47622, x47621, x47620);
  nand n47623(x47623, x38852, x47545);
  nand n47624(x47624, x38913, x47533);
  nand n47625(x47625, x47624, x47623);
  nand n47626(x47626, x38852, x47548);
  nand n47627(x47627, x38913, x47536);
  nand n47628(x47628, x47627, x47626);
  nand n47629(x47629, x38852, x47551);
  nand n47630(x47630, x38913, x47539);
  nand n47631(x47631, x47630, x47629);
  nand n47632(x47632, x38852, x47554);
  nand n47633(x47633, x38913, x47542);
  nand n47634(x47634, x47633, x47632);
  nand n47635(x47635, x38852, x47557);
  nand n47636(x47636, x38913, x47545);
  nand n47637(x47637, x47636, x47635);
  nand n47638(x47638, x38852, x47560);
  nand n47639(x47639, x38913, x47548);
  nand n47640(x47640, x47639, x47638);
  nand n47641(x47641, x38852, x47563);
  nand n47642(x47642, x38913, x47551);
  nand n47643(x47643, x47642, x47641);
  nand n47644(x47644, x38852, x85271);
  nand n47645(x47645, x38913, x47554);
  nand n47646(x47646, x47645, x47644);
  nand n47647(x47647, x38852, x85272);
  nand n47648(x47648, x38913, x47557);
  nand n47649(x47649, x47648, x47647);
  nand n47650(x47650, x38913, x47560);
  nand n47651(x47651, x38913, x47563);
  nand n47652(x47652, x38913, x85271);
  nand n47653(x47653, x38913, x85272);
  nand n47654(x47654, x38854, x47592);
  nand n47655(x47655, x38914, x47568);
  nand n47656(x47656, x47655, x47654);
  nand n47657(x47657, x38854, x47595);
  nand n47658(x47658, x38914, x47571);
  nand n47659(x47659, x47658, x47657);
  nand n47660(x47660, x38854, x47598);
  nand n47661(x47661, x38914, x47574);
  nand n47662(x47662, x47661, x47660);
  nand n47663(x47663, x38854, x47601);
  nand n47664(x47664, x38914, x47577);
  nand n47665(x47665, x47664, x47663);
  nand n47666(x47666, x38854, x47604);
  nand n47667(x47667, x38914, x47580);
  nand n47668(x47668, x47667, x47666);
  nand n47669(x47669, x38854, x47607);
  nand n47670(x47670, x38914, x47583);
  nand n47671(x47671, x47670, x47669);
  nand n47672(x47672, x38854, x47610);
  nand n47673(x47673, x38914, x47586);
  nand n47674(x47674, x47673, x47672);
  nand n47675(x47675, x38854, x47613);
  nand n47676(x47676, x38914, x47589);
  nand n47677(x47677, x47676, x47675);
  nand n47678(x47678, x38854, x47616);
  nand n47679(x47679, x38914, x47592);
  nand n47680(x47680, x47679, x47678);
  nand n47681(x47681, x38854, x47619);
  nand n47682(x47682, x38914, x47595);
  nand n47683(x47683, x47682, x47681);
  nand n47684(x47684, x38854, x47622);
  nand n47685(x47685, x38914, x47598);
  nand n47686(x47686, x47685, x47684);
  nand n47687(x47687, x38854, x47625);
  nand n47688(x47688, x38914, x47601);
  nand n47689(x47689, x47688, x47687);
  nand n47690(x47690, x38854, x47628);
  nand n47691(x47691, x38914, x47604);
  nand n47692(x47692, x47691, x47690);
  nand n47693(x47693, x38854, x47631);
  nand n47694(x47694, x38914, x47607);
  nand n47695(x47695, x47694, x47693);
  nand n47696(x47696, x38854, x47634);
  nand n47697(x47697, x38914, x47610);
  nand n47698(x47698, x47697, x47696);
  nand n47699(x47699, x38854, x47637);
  nand n47700(x47700, x38914, x47613);
  nand n47701(x47701, x47700, x47699);
  nand n47702(x47702, x38854, x47640);
  nand n47703(x47703, x38914, x47616);
  nand n47704(x47704, x47703, x47702);
  nand n47705(x47705, x38854, x47643);
  nand n47706(x47706, x38914, x47619);
  nand n47707(x47707, x47706, x47705);
  nand n47708(x47708, x38854, x47646);
  nand n47709(x47709, x38914, x47622);
  nand n47710(x47710, x47709, x47708);
  nand n47711(x47711, x38854, x47649);
  nand n47712(x47712, x38914, x47625);
  nand n47713(x47713, x47712, x47711);
  nand n47714(x47714, x38854, x85273);
  nand n47715(x47715, x38914, x47628);
  nand n47716(x47716, x47715, x47714);
  nand n47717(x47717, x38854, x85274);
  nand n47718(x47718, x38914, x47631);
  nand n47719(x47719, x47718, x47717);
  nand n47720(x47720, x38854, x85275);
  nand n47721(x47721, x38914, x47634);
  nand n47722(x47722, x47721, x47720);
  nand n47723(x47723, x38854, x85276);
  nand n47724(x47724, x38914, x47637);
  nand n47725(x47725, x47724, x47723);
  nand n47726(x47726, x38914, x47640);
  nand n47727(x47727, x38914, x47643);
  nand n47728(x47728, x38914, x47646);
  nand n47729(x47729, x38914, x47649);
  nand n47730(x47730, x38914, x85273);
  nand n47731(x47731, x38914, x85274);
  nand n47732(x47732, x38914, x85275);
  nand n47733(x47733, x38914, x85276);
  nand n47734(x47734, x38856, x47704);
  nand n47735(x47735, x38915, x47656);
  nand n47736(x47736, x47735, x47734);
  nand n47737(x47737, x38856, x47707);
  nand n47738(x47738, x38915, x47659);
  nand n47739(x47739, x47738, x47737);
  nand n47740(x47740, x38856, x47710);
  nand n47741(x47741, x38915, x47662);
  nand n47742(x47742, x47741, x47740);
  nand n47743(x47743, x38856, x47713);
  nand n47744(x47744, x38915, x47665);
  nand n47745(x47745, x47744, x47743);
  nand n47746(x47746, x38856, x47716);
  nand n47747(x47747, x38915, x47668);
  nand n47748(x47748, x47747, x47746);
  nand n47749(x47749, x38856, x47719);
  nand n47750(x47750, x38915, x47671);
  nand n47751(x47751, x47750, x47749);
  nand n47752(x47752, x38856, x47722);
  nand n47753(x47753, x38915, x47674);
  nand n47754(x47754, x47753, x47752);
  nand n47755(x47755, x38856, x47725);
  nand n47756(x47756, x38915, x47677);
  nand n47757(x47757, x47756, x47755);
  nand n47758(x47758, x38856, x85277);
  nand n47759(x47759, x38915, x47680);
  nand n47760(x47760, x47759, x47758);
  nand n47761(x47761, x38856, x85278);
  nand n47762(x47762, x38915, x47683);
  nand n47763(x47763, x47762, x47761);
  nand n47764(x47764, x38856, x85279);
  nand n47765(x47765, x38915, x47686);
  nand n47766(x47766, x47765, x47764);
  nand n47767(x47767, x38856, x85280);
  nand n47768(x47768, x38915, x47689);
  nand n47769(x47769, x47768, x47767);
  nand n47770(x47770, x38856, x85281);
  nand n47771(x47771, x38915, x47692);
  nand n47772(x47772, x47771, x47770);
  nand n47773(x47773, x38856, x85282);
  nand n47774(x47774, x38915, x47695);
  nand n47775(x47775, x47774, x47773);
  nand n47776(x47776, x38856, x85283);
  nand n47777(x47777, x38915, x47698);
  nand n47778(x47778, x47777, x47776);
  nand n47779(x47779, x38856, x85284);
  nand n47780(x47780, x38915, x47701);
  nand n47781(x47781, x47780, x47779);
  nand n47782(x47782, x38915, x47704);
  nand n47783(x47783, x38915, x47707);
  nand n47784(x47784, x38915, x47710);
  nand n47785(x47785, x38915, x47713);
  nand n47786(x47786, x38915, x47716);
  nand n47787(x47787, x38915, x47719);
  nand n47788(x47788, x38915, x47722);
  nand n47789(x47789, x38915, x47725);
  nand n47790(x47790, x38915, x85277);
  nand n47791(x47791, x38915, x85278);
  nand n47792(x47792, x38915, x85279);
  nand n47793(x47793, x38915, x85280);
  nand n47794(x47794, x38915, x85281);
  nand n47795(x47795, x38915, x85282);
  nand n47796(x47796, x38915, x85283);
  nand n47797(x47797, x38915, x85284);
  nand n47798(x47798, x71977, x38848);
  nand n47799(x47799, x16876, x47736);
  nand n47800(x47800, x47799, x25733);
  nand n47801(x47801, x71977, x85254);
  nand n47802(x47802, x16876, x46927);
  nand n47803(x47803, x71977, x39815);
  nand n47804(x47804, x16876, x39815);
  nand n47805(x47805, x47804, x47803);
  nand n47806(x47806, x71977, x46993);
  nand n47807(x47807, x16876, x46960);
  nand n47808(x47808, x47807, x47806);
  nand n47809(x47809, x71977, x46927);
  nand n47810(x47810, x47799, x47809);
  nand n47811(x47811, x16876, x39041);
  nand n47812(x47812, x47811, x47809);
  nand n47813(x47813, x71977, x73027);
  nand n47814(x47814, x25749, x85301);
  nand n47815(x47815, x71982, x47800);
  nand n47816(x47816, x25749, x85302);
  nand n47817(x47817, x47816, x47815);
  nand n47818(x47818, x71982, x85303);
  nand n47819(x47819, x25749, x47805);
  nand n47820(x47820, x47819, x47818);
  nand n47821(x47821, x71982, x47808);
  nand n47822(x47822, x25749, x47810);
  nand n47823(x47823, x47822, x47821);
  nand n47824(x47824, x71982, x85302);
  nand n47825(x47825, x25749, x85303);
  nand n47826(x47826, x47825, x47824);
  nand n47827(x47827, x71982, x47805);
  nand n47828(x47828, x25749, x47808);
  nand n47829(x47829, x47828, x47827);
  nand n47830(x47830, x71982, x47812);
  nand n47831(x47831, x25749, x85304);
  nand n47832(x47832, x47831, x47830);
  nand n47833(x47833, x71987, x85305);
  nand n47834(x47834, x25772, x47817);
  nand n47835(x47835, x47834, x25771);
  nand n47836(x47836, x71987, x47820);
  nand n47837(x47837, x25772, x47823);
  nand n47838(x47838, x47837, x47836);
  nand n47839(x47839, x71987, x47826);
  nand n47840(x47840, x25772, x47829);
  nand n47841(x47841, x47840, x47839);
  nand n47842(x47842, x71987, x47832);
  nand n47843(x47843, x25782, x85306);
  nand n47844(x47844, x71992, x47835);
  nand n47845(x47845, x25782, x47838);
  nand n47846(x47846, x47845, x47844);
  nand n47847(x47847, x71992, x47841);
  nand n47848(x47848, x25782, x85307);
  nand n47849(x47849, x47848, x47847);
  nand n47850(x47850, x25790, x85308);
  nand n47851(x47851, x71997, x47846);
  nand n47852(x47852, x25790, x47849);
  nand n47853(x47853, x47852, x47851);
  nand n47854(x47854, x72002, x85309);
  nand n47855(x47855, x25796, x47853);
  nand n47856(x47856, x47855, x47854);
  nand n47857(x47857, x71977, x38850);
  nand n47858(x47858, x16876, x47739);
  nand n47859(x47859, x47858, x25801);
  nand n47860(x47860, x71977, x85255);
  nand n47861(x47861, x16876, x85207);
  nand n47862(x47862, x71977, x39820);
  nand n47863(x47863, x16876, x39820);
  nand n47864(x47864, x47863, x47862);
  nand n47865(x47865, x71977, x46995);
  nand n47866(x47866, x16876, x46961);
  nand n47867(x47867, x47866, x47865);
  nand n47868(x47868, x71977, x39979);
  nand n47869(x47869, x47858, x47868);
  nand n47870(x47870, x16876, x39047);
  nand n47871(x47871, x47870, x47868);
  nand n47872(x47872, x71977, x46806);
  nand n47873(x47873, x25749, x85310);
  nand n47874(x47874, x71982, x47859);
  nand n47875(x47875, x25749, x85311);
  nand n47876(x47876, x47875, x47874);
  nand n47877(x47877, x71982, x85312);
  nand n47878(x47878, x25749, x47864);
  nand n47879(x47879, x47878, x47877);
  nand n47880(x47880, x71982, x47867);
  nand n47881(x47881, x25749, x47869);
  nand n47882(x47882, x47881, x47880);
  nand n47883(x47883, x71982, x85311);
  nand n47884(x47884, x25749, x85312);
  nand n47885(x47885, x47884, x47883);
  nand n47886(x47886, x71982, x47864);
  nand n47887(x47887, x25749, x47867);
  nand n47888(x47888, x47887, x47886);
  nand n47889(x47889, x71982, x47871);
  nand n47890(x47890, x25749, x85313);
  nand n47891(x47891, x47890, x47889);
  nand n47892(x47892, x71987, x85314);
  nand n47893(x47893, x25772, x47876);
  nand n47894(x47894, x47893, x25838);
  nand n47895(x47895, x71987, x47879);
  nand n47896(x47896, x25772, x47882);
  nand n47897(x47897, x47896, x47895);
  nand n47898(x47898, x71987, x47885);
  nand n47899(x47899, x25772, x47888);
  nand n47900(x47900, x47899, x47898);
  nand n47901(x47901, x71987, x47891);
  nand n47902(x47902, x25782, x85315);
  nand n47903(x47903, x71992, x47894);
  nand n47904(x47904, x25782, x47897);
  nand n47905(x47905, x47904, x47903);
  nand n47906(x47906, x71992, x47900);
  nand n47907(x47907, x25782, x85316);
  nand n47908(x47908, x47907, x47906);
  nand n47909(x47909, x25790, x85317);
  nand n47910(x47910, x71997, x47905);
  nand n47911(x47911, x25790, x47908);
  nand n47912(x47912, x47911, x47910);
  nand n47913(x47913, x72002, x85318);
  nand n47914(x47914, x25796, x47912);
  nand n47915(x47915, x47914, x47913);
  nand n47916(x47916, x71977, x38852);
  nand n47917(x47917, x16876, x47742);
  nand n47918(x47918, x47917, x25864);
  nand n47919(x47919, x71977, x85256);
  nand n47920(x47920, x16876, x85208);
  nand n47921(x47921, x71977, x39825);
  nand n47922(x47922, x16876, x39825);
  nand n47923(x47923, x47922, x47921);
  nand n47924(x47924, x71977, x46997);
  nand n47925(x47925, x16876, x46962);
  nand n47926(x47926, x47925, x47924);
  nand n47927(x47927, x71977, x39994);
  nand n47928(x47928, x47917, x47927);
  nand n47929(x47929, x16876, x39053);
  nand n47930(x47930, x47929, x47927);
  nand n47931(x47931, x71977, x46810);
  nand n47932(x47932, x25749, x85319);
  nand n47933(x47933, x71982, x47918);
  nand n47934(x47934, x25749, x85320);
  nand n47935(x47935, x47934, x47933);
  nand n47936(x47936, x71982, x85321);
  nand n47937(x47937, x25749, x47923);
  nand n47938(x47938, x47937, x47936);
  nand n47939(x47939, x71982, x47926);
  nand n47940(x47940, x25749, x47928);
  nand n47941(x47941, x47940, x47939);
  nand n47942(x47942, x71982, x85320);
  nand n47943(x47943, x25749, x85321);
  nand n47944(x47944, x47943, x47942);
  nand n47945(x47945, x71982, x47923);
  nand n47946(x47946, x25749, x47926);
  nand n47947(x47947, x47946, x47945);
  nand n47948(x47948, x71982, x47930);
  nand n47949(x47949, x25749, x85322);
  nand n47950(x47950, x47949, x47948);
  nand n47951(x47951, x71987, x85323);
  nand n47952(x47952, x25772, x47935);
  nand n47953(x47953, x47952, x25901);
  nand n47954(x47954, x71987, x47938);
  nand n47955(x47955, x25772, x47941);
  nand n47956(x47956, x47955, x47954);
  nand n47957(x47957, x71987, x47944);
  nand n47958(x47958, x25772, x47947);
  nand n47959(x47959, x47958, x47957);
  nand n47960(x47960, x71987, x47950);
  nand n47961(x47961, x25782, x85324);
  nand n47962(x47962, x71992, x47953);
  nand n47963(x47963, x25782, x47956);
  nand n47964(x47964, x47963, x47962);
  nand n47965(x47965, x71992, x47959);
  nand n47966(x47966, x25782, x85325);
  nand n47967(x47967, x47966, x47965);
  nand n47968(x47968, x25790, x85326);
  nand n47969(x47969, x71997, x47964);
  nand n47970(x47970, x25790, x47967);
  nand n47971(x47971, x47970, x47969);
  nand n47972(x47972, x72002, x85327);
  nand n47973(x47973, x25796, x47971);
  nand n47974(x47974, x47973, x47972);
  nand n47975(x47975, x71977, x38854);
  nand n47976(x47976, x16876, x47745);
  nand n47977(x47977, x47976, x25927);
  nand n47978(x47978, x71977, x85257);
  nand n47979(x47979, x16876, x85209);
  nand n47980(x47980, x71977, x39830);
  nand n47981(x47981, x16876, x39830);
  nand n47982(x47982, x47981, x47980);
  nand n47983(x47983, x71977, x46999);
  nand n47984(x47984, x16876, x46963);
  nand n47985(x47985, x47984, x47983);
  nand n47986(x47986, x71977, x40018);
  nand n47987(x47987, x47976, x47986);
  nand n47988(x47988, x16876, x39059);
  nand n47989(x47989, x47988, x47986);
  nand n47990(x47990, x71977, x46814);
  nand n47991(x47991, x25749, x85328);
  nand n47992(x47992, x71982, x47977);
  nand n47993(x47993, x25749, x85329);
  nand n47994(x47994, x47993, x47992);
  nand n47995(x47995, x71982, x85330);
  nand n47996(x47996, x25749, x47982);
  nand n47997(x47997, x47996, x47995);
  nand n47998(x47998, x71982, x47985);
  nand n47999(x47999, x25749, x47987);
  nand n48000(x48000, x47999, x47998);
  nand n48001(x48001, x71982, x85329);
  nand n48002(x48002, x25749, x85330);
  nand n48003(x48003, x48002, x48001);
  nand n48004(x48004, x71982, x47982);
  nand n48005(x48005, x25749, x47985);
  nand n48006(x48006, x48005, x48004);
  nand n48007(x48007, x71982, x47989);
  nand n48008(x48008, x25749, x85331);
  nand n48009(x48009, x48008, x48007);
  nand n48010(x48010, x71987, x85332);
  nand n48011(x48011, x25772, x47994);
  nand n48012(x48012, x48011, x25964);
  nand n48013(x48013, x71987, x47997);
  nand n48014(x48014, x25772, x48000);
  nand n48015(x48015, x48014, x48013);
  nand n48016(x48016, x71987, x48003);
  nand n48017(x48017, x25772, x48006);
  nand n48018(x48018, x48017, x48016);
  nand n48019(x48019, x71987, x48009);
  nand n48020(x48020, x25782, x85333);
  nand n48021(x48021, x71992, x48012);
  nand n48022(x48022, x25782, x48015);
  nand n48023(x48023, x48022, x48021);
  nand n48024(x48024, x71992, x48018);
  nand n48025(x48025, x25782, x85334);
  nand n48026(x48026, x48025, x48024);
  nand n48027(x48027, x25790, x85335);
  nand n48028(x48028, x71997, x48023);
  nand n48029(x48029, x25790, x48026);
  nand n48030(x48030, x48029, x48028);
  nand n48031(x48031, x72002, x85336);
  nand n48032(x48032, x25796, x48030);
  nand n48033(x48033, x48032, x48031);
  nand n48034(x48034, x71977, x38856);
  nand n48035(x48035, x16876, x47748);
  nand n48036(x48036, x48035, x25990);
  nand n48037(x48037, x71977, x85258);
  nand n48038(x48038, x16876, x85210);
  nand n48039(x48039, x71977, x39835);
  nand n48040(x48040, x16876, x39835);
  nand n48041(x48041, x48040, x48039);
  nand n48042(x48042, x71977, x47001);
  nand n48043(x48043, x16876, x46964);
  nand n48044(x48044, x48043, x48042);
  nand n48045(x48045, x71977, x40049);
  nand n48046(x48046, x48035, x48045);
  nand n48047(x48047, x16876, x39065);
  nand n48048(x48048, x48047, x48045);
  nand n48049(x48049, x71977, x46818);
  nand n48050(x48050, x25749, x85337);
  nand n48051(x48051, x71982, x48036);
  nand n48052(x48052, x25749, x85338);
  nand n48053(x48053, x48052, x48051);
  nand n48054(x48054, x71982, x85339);
  nand n48055(x48055, x25749, x48041);
  nand n48056(x48056, x48055, x48054);
  nand n48057(x48057, x71982, x48044);
  nand n48058(x48058, x25749, x48046);
  nand n48059(x48059, x48058, x48057);
  nand n48060(x48060, x71982, x85338);
  nand n48061(x48061, x25749, x85339);
  nand n48062(x48062, x48061, x48060);
  nand n48063(x48063, x71982, x48041);
  nand n48064(x48064, x25749, x48044);
  nand n48065(x48065, x48064, x48063);
  nand n48066(x48066, x71982, x48048);
  nand n48067(x48067, x25749, x85340);
  nand n48068(x48068, x48067, x48066);
  nand n48069(x48069, x71987, x85341);
  nand n48070(x48070, x25772, x48053);
  nand n48071(x48071, x48070, x26027);
  nand n48072(x48072, x71987, x48056);
  nand n48073(x48073, x25772, x48059);
  nand n48074(x48074, x48073, x48072);
  nand n48075(x48075, x71987, x48062);
  nand n48076(x48076, x25772, x48065);
  nand n48077(x48077, x48076, x48075);
  nand n48078(x48078, x71987, x48068);
  nand n48079(x48079, x25782, x85342);
  nand n48080(x48080, x71992, x48071);
  nand n48081(x48081, x25782, x48074);
  nand n48082(x48082, x48081, x48080);
  nand n48083(x48083, x71992, x48077);
  nand n48084(x48084, x25782, x85343);
  nand n48085(x48085, x48084, x48083);
  nand n48086(x48086, x25790, x85344);
  nand n48087(x48087, x71997, x48082);
  nand n48088(x48088, x25790, x48085);
  nand n48089(x48089, x48088, x48087);
  nand n48090(x48090, x72002, x85345);
  nand n48091(x48091, x25796, x48089);
  nand n48092(x48092, x48091, x48090);
  nand n48093(x48093, x71977, x38858);
  nand n48094(x48094, x16876, x47751);
  nand n48095(x48095, x48094, x26053);
  nand n48096(x48096, x71977, x85259);
  nand n48097(x48097, x16876, x85211);
  nand n48098(x48098, x71977, x39840);
  nand n48099(x48099, x16876, x39840);
  nand n48100(x48100, x48099, x48098);
  nand n48101(x48101, x71977, x47003);
  nand n48102(x48102, x16876, x46965);
  nand n48103(x48103, x48102, x48101);
  nand n48104(x48104, x71977, x40088);
  nand n48105(x48105, x48094, x48104);
  nand n48106(x48106, x16876, x39071);
  nand n48107(x48107, x48106, x48104);
  nand n48108(x48108, x71977, x46822);
  nand n48109(x48109, x25749, x85346);
  nand n48110(x48110, x71982, x48095);
  nand n48111(x48111, x25749, x85347);
  nand n48112(x48112, x48111, x48110);
  nand n48113(x48113, x71982, x85348);
  nand n48114(x48114, x25749, x48100);
  nand n48115(x48115, x48114, x48113);
  nand n48116(x48116, x71982, x48103);
  nand n48117(x48117, x25749, x48105);
  nand n48118(x48118, x48117, x48116);
  nand n48119(x48119, x71982, x85347);
  nand n48120(x48120, x25749, x85348);
  nand n48121(x48121, x48120, x48119);
  nand n48122(x48122, x71982, x48100);
  nand n48123(x48123, x25749, x48103);
  nand n48124(x48124, x48123, x48122);
  nand n48125(x48125, x71982, x48107);
  nand n48126(x48126, x25749, x85349);
  nand n48127(x48127, x48126, x48125);
  nand n48128(x48128, x71987, x85350);
  nand n48129(x48129, x25772, x48112);
  nand n48130(x48130, x48129, x26090);
  nand n48131(x48131, x71987, x48115);
  nand n48132(x48132, x25772, x48118);
  nand n48133(x48133, x48132, x48131);
  nand n48134(x48134, x71987, x48121);
  nand n48135(x48135, x25772, x48124);
  nand n48136(x48136, x48135, x48134);
  nand n48137(x48137, x71987, x48127);
  nand n48138(x48138, x25782, x85351);
  nand n48139(x48139, x71992, x48130);
  nand n48140(x48140, x25782, x48133);
  nand n48141(x48141, x48140, x48139);
  nand n48142(x48142, x71992, x48136);
  nand n48143(x48143, x25782, x85352);
  nand n48144(x48144, x48143, x48142);
  nand n48145(x48145, x25790, x85353);
  nand n48146(x48146, x71997, x48141);
  nand n48147(x48147, x25790, x48144);
  nand n48148(x48148, x48147, x48146);
  nand n48149(x48149, x72002, x85354);
  nand n48150(x48150, x25796, x48148);
  nand n48151(x48151, x48150, x48149);
  nand n48152(x48152, x71977, x38860);
  nand n48153(x48153, x16876, x47754);
  nand n48154(x48154, x48153, x26116);
  nand n48155(x48155, x71977, x85260);
  nand n48156(x48156, x16876, x46470);
  nand n48157(x48157, x71977, x39845);
  nand n48158(x48158, x16876, x39845);
  nand n48159(x48159, x48158, x48157);
  nand n48160(x48160, x71977, x47005);
  nand n48161(x48161, x16876, x46966);
  nand n48162(x48162, x48161, x48160);
  nand n48163(x48163, x71977, x40136);
  nand n48164(x48164, x48153, x48163);
  nand n48165(x48165, x16876, x39077);
  nand n48166(x48166, x48165, x48163);
  nand n48167(x48167, x71977, x46826);
  nand n48168(x48168, x25749, x85355);
  nand n48169(x48169, x71982, x48154);
  nand n48170(x48170, x25749, x85356);
  nand n48171(x48171, x48170, x48169);
  nand n48172(x48172, x71982, x85357);
  nand n48173(x48173, x25749, x48159);
  nand n48174(x48174, x48173, x48172);
  nand n48175(x48175, x71982, x48162);
  nand n48176(x48176, x25749, x48164);
  nand n48177(x48177, x48176, x48175);
  nand n48178(x48178, x71982, x85356);
  nand n48179(x48179, x25749, x85357);
  nand n48180(x48180, x48179, x48178);
  nand n48181(x48181, x71982, x48159);
  nand n48182(x48182, x25749, x48162);
  nand n48183(x48183, x48182, x48181);
  nand n48184(x48184, x71982, x48166);
  nand n48185(x48185, x25749, x85358);
  nand n48186(x48186, x48185, x48184);
  nand n48187(x48187, x71987, x85359);
  nand n48188(x48188, x25772, x48171);
  nand n48189(x48189, x48188, x26153);
  nand n48190(x48190, x71987, x48174);
  nand n48191(x48191, x25772, x48177);
  nand n48192(x48192, x48191, x48190);
  nand n48193(x48193, x71987, x48180);
  nand n48194(x48194, x25772, x48183);
  nand n48195(x48195, x48194, x48193);
  nand n48196(x48196, x71987, x48186);
  nand n48197(x48197, x25782, x85360);
  nand n48198(x48198, x71992, x48189);
  nand n48199(x48199, x25782, x48192);
  nand n48200(x48200, x48199, x48198);
  nand n48201(x48201, x71992, x48195);
  nand n48202(x48202, x25782, x85361);
  nand n48203(x48203, x48202, x48201);
  nand n48204(x48204, x25790, x85362);
  nand n48205(x48205, x71997, x48200);
  nand n48206(x48206, x25790, x48203);
  nand n48207(x48207, x48206, x48205);
  nand n48208(x48208, x72002, x85363);
  nand n48209(x48209, x25796, x48207);
  nand n48210(x48210, x48209, x48208);
  nand n48211(x48211, x71977, x38862);
  nand n48212(x48212, x16876, x47757);
  nand n48213(x48213, x48212, x26179);
  nand n48214(x48214, x71977, x85261);
  nand n48215(x48215, x16876, x46474);
  nand n48216(x48216, x71977, x39850);
  nand n48217(x48217, x16876, x39850);
  nand n48218(x48218, x48217, x48216);
  nand n48219(x48219, x71977, x47007);
  nand n48220(x48220, x16876, x46967);
  nand n48221(x48221, x48220, x48219);
  nand n48222(x48222, x71977, x40191);
  nand n48223(x48223, x48212, x48222);
  nand n48224(x48224, x16876, x39083);
  nand n48225(x48225, x48224, x48222);
  nand n48226(x48226, x71977, x46830);
  nand n48227(x48227, x25749, x85364);
  nand n48228(x48228, x71982, x48213);
  nand n48229(x48229, x25749, x85365);
  nand n48230(x48230, x48229, x48228);
  nand n48231(x48231, x71982, x85366);
  nand n48232(x48232, x25749, x48218);
  nand n48233(x48233, x48232, x48231);
  nand n48234(x48234, x71982, x48221);
  nand n48235(x48235, x25749, x48223);
  nand n48236(x48236, x48235, x48234);
  nand n48237(x48237, x71982, x85365);
  nand n48238(x48238, x25749, x85366);
  nand n48239(x48239, x48238, x48237);
  nand n48240(x48240, x71982, x48218);
  nand n48241(x48241, x25749, x48221);
  nand n48242(x48242, x48241, x48240);
  nand n48243(x48243, x71982, x48225);
  nand n48244(x48244, x25749, x85367);
  nand n48245(x48245, x48244, x48243);
  nand n48246(x48246, x71987, x85368);
  nand n48247(x48247, x25772, x48230);
  nand n48248(x48248, x48247, x26216);
  nand n48249(x48249, x71987, x48233);
  nand n48250(x48250, x25772, x48236);
  nand n48251(x48251, x48250, x48249);
  nand n48252(x48252, x71987, x48239);
  nand n48253(x48253, x25772, x48242);
  nand n48254(x48254, x48253, x48252);
  nand n48255(x48255, x71987, x48245);
  nand n48256(x48256, x25782, x85369);
  nand n48257(x48257, x71992, x48248);
  nand n48258(x48258, x25782, x48251);
  nand n48259(x48259, x48258, x48257);
  nand n48260(x48260, x71992, x48254);
  nand n48261(x48261, x25782, x85370);
  nand n48262(x48262, x48261, x48260);
  nand n48263(x48263, x25790, x85371);
  nand n48264(x48264, x71997, x48259);
  nand n48265(x48265, x25790, x48262);
  nand n48266(x48266, x48265, x48264);
  nand n48267(x48267, x72002, x85372);
  nand n48268(x48268, x25796, x48266);
  nand n48269(x48269, x48268, x48267);
  nand n48270(x48270, x71977, x38864);
  nand n48271(x48271, x16876, x47760);
  nand n48272(x48272, x48271, x26242);
  nand n48273(x48273, x71977, x85262);
  nand n48274(x48274, x16876, x46478);
  nand n48275(x48275, x71977, x39855);
  nand n48276(x48276, x16876, x39855);
  nand n48277(x48277, x48276, x48275);
  nand n48278(x48278, x71977, x47009);
  nand n48279(x48279, x16876, x46968);
  nand n48280(x48280, x48279, x48278);
  nand n48281(x48281, x71977, x40254);
  nand n48282(x48282, x48271, x48281);
  nand n48283(x48283, x16876, x39089);
  nand n48284(x48284, x48283, x48281);
  nand n48285(x48285, x71977, x46834);
  nand n48286(x48286, x25749, x85373);
  nand n48287(x48287, x71982, x48272);
  nand n48288(x48288, x25749, x85374);
  nand n48289(x48289, x48288, x48287);
  nand n48290(x48290, x71982, x85375);
  nand n48291(x48291, x25749, x48277);
  nand n48292(x48292, x48291, x48290);
  nand n48293(x48293, x71982, x48280);
  nand n48294(x48294, x25749, x48282);
  nand n48295(x48295, x48294, x48293);
  nand n48296(x48296, x71982, x85374);
  nand n48297(x48297, x25749, x85375);
  nand n48298(x48298, x48297, x48296);
  nand n48299(x48299, x71982, x48277);
  nand n48300(x48300, x25749, x48280);
  nand n48301(x48301, x48300, x48299);
  nand n48302(x48302, x71982, x48284);
  nand n48303(x48303, x25749, x85376);
  nand n48304(x48304, x48303, x48302);
  nand n48305(x48305, x71987, x85377);
  nand n48306(x48306, x25772, x48289);
  nand n48307(x48307, x48306, x26279);
  nand n48308(x48308, x71987, x48292);
  nand n48309(x48309, x25772, x48295);
  nand n48310(x48310, x48309, x48308);
  nand n48311(x48311, x71987, x48298);
  nand n48312(x48312, x25772, x48301);
  nand n48313(x48313, x48312, x48311);
  nand n48314(x48314, x71987, x48304);
  nand n48315(x48315, x25782, x85378);
  nand n48316(x48316, x71992, x48307);
  nand n48317(x48317, x25782, x48310);
  nand n48318(x48318, x48317, x48316);
  nand n48319(x48319, x71992, x48313);
  nand n48320(x48320, x25782, x85379);
  nand n48321(x48321, x48320, x48319);
  nand n48322(x48322, x25790, x85380);
  nand n48323(x48323, x71997, x48318);
  nand n48324(x48324, x25790, x48321);
  nand n48325(x48325, x48324, x48323);
  nand n48326(x48326, x72002, x85381);
  nand n48327(x48327, x25796, x48325);
  nand n48328(x48328, x48327, x48326);
  nand n48329(x48329, x71977, x38866);
  nand n48330(x48330, x16876, x47763);
  nand n48331(x48331, x48330, x26305);
  nand n48332(x48332, x71977, x85263);
  nand n48333(x48333, x16876, x46482);
  nand n48334(x48334, x71977, x39860);
  nand n48335(x48335, x16876, x39860);
  nand n48336(x48336, x48335, x48334);
  nand n48337(x48337, x71977, x47011);
  nand n48338(x48338, x16876, x46969);
  nand n48339(x48339, x48338, x48337);
  nand n48340(x48340, x71977, x40326);
  nand n48341(x48341, x48330, x48340);
  nand n48342(x48342, x16876, x39095);
  nand n48343(x48343, x48342, x48340);
  nand n48344(x48344, x71977, x46838);
  nand n48345(x48345, x25749, x85382);
  nand n48346(x48346, x71982, x48331);
  nand n48347(x48347, x25749, x85383);
  nand n48348(x48348, x48347, x48346);
  nand n48349(x48349, x71982, x85384);
  nand n48350(x48350, x25749, x48336);
  nand n48351(x48351, x48350, x48349);
  nand n48352(x48352, x71982, x48339);
  nand n48353(x48353, x25749, x48341);
  nand n48354(x48354, x48353, x48352);
  nand n48355(x48355, x71982, x85383);
  nand n48356(x48356, x25749, x85384);
  nand n48357(x48357, x48356, x48355);
  nand n48358(x48358, x71982, x48336);
  nand n48359(x48359, x25749, x48339);
  nand n48360(x48360, x48359, x48358);
  nand n48361(x48361, x71982, x48343);
  nand n48362(x48362, x25749, x85385);
  nand n48363(x48363, x48362, x48361);
  nand n48364(x48364, x71987, x85386);
  nand n48365(x48365, x25772, x48348);
  nand n48366(x48366, x48365, x26342);
  nand n48367(x48367, x71987, x48351);
  nand n48368(x48368, x25772, x48354);
  nand n48369(x48369, x48368, x48367);
  nand n48370(x48370, x71987, x48357);
  nand n48371(x48371, x25772, x48360);
  nand n48372(x48372, x48371, x48370);
  nand n48373(x48373, x71987, x48363);
  nand n48374(x48374, x25782, x85387);
  nand n48375(x48375, x71992, x48366);
  nand n48376(x48376, x25782, x48369);
  nand n48377(x48377, x48376, x48375);
  nand n48378(x48378, x71992, x48372);
  nand n48379(x48379, x25782, x85388);
  nand n48380(x48380, x48379, x48378);
  nand n48381(x48381, x25790, x85389);
  nand n48382(x48382, x71997, x48377);
  nand n48383(x48383, x25790, x48380);
  nand n48384(x48384, x48383, x48382);
  nand n48385(x48385, x72002, x85390);
  nand n48386(x48386, x25796, x48384);
  nand n48387(x48387, x48386, x48385);
  nand n48388(x48388, x71977, x38868);
  nand n48389(x48389, x16876, x47766);
  nand n48390(x48390, x48389, x26368);
  nand n48391(x48391, x71977, x85264);
  nand n48392(x48392, x16876, x46486);
  nand n48393(x48393, x71977, x39865);
  nand n48394(x48394, x16876, x39865);
  nand n48395(x48395, x48394, x48393);
  nand n48396(x48396, x71977, x47013);
  nand n48397(x48397, x16876, x46970);
  nand n48398(x48398, x48397, x48396);
  nand n48399(x48399, x71977, x40405);
  nand n48400(x48400, x48389, x48399);
  nand n48401(x48401, x16876, x39101);
  nand n48402(x48402, x48401, x48399);
  nand n48403(x48403, x71977, x46842);
  nand n48404(x48404, x25749, x85391);
  nand n48405(x48405, x71982, x48390);
  nand n48406(x48406, x25749, x85392);
  nand n48407(x48407, x48406, x48405);
  nand n48408(x48408, x71982, x85393);
  nand n48409(x48409, x25749, x48395);
  nand n48410(x48410, x48409, x48408);
  nand n48411(x48411, x71982, x48398);
  nand n48412(x48412, x25749, x48400);
  nand n48413(x48413, x48412, x48411);
  nand n48414(x48414, x71982, x85392);
  nand n48415(x48415, x25749, x85393);
  nand n48416(x48416, x48415, x48414);
  nand n48417(x48417, x71982, x48395);
  nand n48418(x48418, x25749, x48398);
  nand n48419(x48419, x48418, x48417);
  nand n48420(x48420, x71982, x48402);
  nand n48421(x48421, x25749, x85394);
  nand n48422(x48422, x48421, x48420);
  nand n48423(x48423, x71987, x85395);
  nand n48424(x48424, x25772, x48407);
  nand n48425(x48425, x48424, x26405);
  nand n48426(x48426, x71987, x48410);
  nand n48427(x48427, x25772, x48413);
  nand n48428(x48428, x48427, x48426);
  nand n48429(x48429, x71987, x48416);
  nand n48430(x48430, x25772, x48419);
  nand n48431(x48431, x48430, x48429);
  nand n48432(x48432, x71987, x48422);
  nand n48433(x48433, x25782, x85396);
  nand n48434(x48434, x71992, x48425);
  nand n48435(x48435, x25782, x48428);
  nand n48436(x48436, x48435, x48434);
  nand n48437(x48437, x71992, x48431);
  nand n48438(x48438, x25782, x85397);
  nand n48439(x48439, x48438, x48437);
  nand n48440(x48440, x25790, x85398);
  nand n48441(x48441, x71997, x48436);
  nand n48442(x48442, x25790, x48439);
  nand n48443(x48443, x48442, x48441);
  nand n48444(x48444, x72002, x85399);
  nand n48445(x48445, x25796, x48443);
  nand n48446(x48446, x48445, x48444);
  nand n48447(x48447, x71977, x38870);
  nand n48448(x48448, x16876, x47769);
  nand n48449(x48449, x48448, x26431);
  nand n48450(x48450, x71977, x85265);
  nand n48451(x48451, x16876, x46490);
  nand n48452(x48452, x71977, x39870);
  nand n48453(x48453, x16876, x39870);
  nand n48454(x48454, x48453, x48452);
  nand n48455(x48455, x71977, x47015);
  nand n48456(x48456, x16876, x46971);
  nand n48457(x48457, x48456, x48455);
  nand n48458(x48458, x71977, x40492);
  nand n48459(x48459, x48448, x48458);
  nand n48460(x48460, x16876, x39107);
  nand n48461(x48461, x48460, x48458);
  nand n48462(x48462, x71977, x46846);
  nand n48463(x48463, x25749, x85400);
  nand n48464(x48464, x71982, x48449);
  nand n48465(x48465, x25749, x85401);
  nand n48466(x48466, x48465, x48464);
  nand n48467(x48467, x71982, x85402);
  nand n48468(x48468, x25749, x48454);
  nand n48469(x48469, x48468, x48467);
  nand n48470(x48470, x71982, x48457);
  nand n48471(x48471, x25749, x48459);
  nand n48472(x48472, x48471, x48470);
  nand n48473(x48473, x71982, x85401);
  nand n48474(x48474, x25749, x85402);
  nand n48475(x48475, x48474, x48473);
  nand n48476(x48476, x71982, x48454);
  nand n48477(x48477, x25749, x48457);
  nand n48478(x48478, x48477, x48476);
  nand n48479(x48479, x71982, x48461);
  nand n48480(x48480, x25749, x85403);
  nand n48481(x48481, x48480, x48479);
  nand n48482(x48482, x71987, x85404);
  nand n48483(x48483, x25772, x48466);
  nand n48484(x48484, x48483, x26468);
  nand n48485(x48485, x71987, x48469);
  nand n48486(x48486, x25772, x48472);
  nand n48487(x48487, x48486, x48485);
  nand n48488(x48488, x71987, x48475);
  nand n48489(x48489, x25772, x48478);
  nand n48490(x48490, x48489, x48488);
  nand n48491(x48491, x71987, x48481);
  nand n48492(x48492, x25782, x85405);
  nand n48493(x48493, x71992, x48484);
  nand n48494(x48494, x25782, x48487);
  nand n48495(x48495, x48494, x48493);
  nand n48496(x48496, x71992, x48490);
  nand n48497(x48497, x25782, x85406);
  nand n48498(x48498, x48497, x48496);
  nand n48499(x48499, x25790, x85407);
  nand n48500(x48500, x71997, x48495);
  nand n48501(x48501, x25790, x48498);
  nand n48502(x48502, x48501, x48500);
  nand n48503(x48503, x72002, x85408);
  nand n48504(x48504, x25796, x48502);
  nand n48505(x48505, x48504, x48503);
  nand n48506(x48506, x71977, x38872);
  nand n48507(x48507, x16876, x47772);
  nand n48508(x48508, x48507, x26494);
  nand n48509(x48509, x71977, x85266);
  nand n48510(x48510, x16876, x46494);
  nand n48511(x48511, x71977, x39875);
  nand n48512(x48512, x16876, x39875);
  nand n48513(x48513, x48512, x48511);
  nand n48514(x48514, x71977, x47017);
  nand n48515(x48515, x16876, x46972);
  nand n48516(x48516, x48515, x48514);
  nand n48517(x48517, x71977, x40588);
  nand n48518(x48518, x48507, x48517);
  nand n48519(x48519, x16876, x39113);
  nand n48520(x48520, x48519, x48517);
  nand n48521(x48521, x71977, x46850);
  nand n48522(x48522, x25749, x85409);
  nand n48523(x48523, x71982, x48508);
  nand n48524(x48524, x25749, x85410);
  nand n48525(x48525, x48524, x48523);
  nand n48526(x48526, x71982, x85411);
  nand n48527(x48527, x25749, x48513);
  nand n48528(x48528, x48527, x48526);
  nand n48529(x48529, x71982, x48516);
  nand n48530(x48530, x25749, x48518);
  nand n48531(x48531, x48530, x48529);
  nand n48532(x48532, x71982, x85410);
  nand n48533(x48533, x25749, x85411);
  nand n48534(x48534, x48533, x48532);
  nand n48535(x48535, x71982, x48513);
  nand n48536(x48536, x25749, x48516);
  nand n48537(x48537, x48536, x48535);
  nand n48538(x48538, x71982, x48520);
  nand n48539(x48539, x25749, x85412);
  nand n48540(x48540, x48539, x48538);
  nand n48541(x48541, x71987, x85413);
  nand n48542(x48542, x25772, x48525);
  nand n48543(x48543, x48542, x26531);
  nand n48544(x48544, x71987, x48528);
  nand n48545(x48545, x25772, x48531);
  nand n48546(x48546, x48545, x48544);
  nand n48547(x48547, x71987, x48534);
  nand n48548(x48548, x25772, x48537);
  nand n48549(x48549, x48548, x48547);
  nand n48550(x48550, x71987, x48540);
  nand n48551(x48551, x25782, x85414);
  nand n48552(x48552, x71992, x48543);
  nand n48553(x48553, x25782, x48546);
  nand n48554(x48554, x48553, x48552);
  nand n48555(x48555, x71992, x48549);
  nand n48556(x48556, x25782, x85415);
  nand n48557(x48557, x48556, x48555);
  nand n48558(x48558, x25790, x85416);
  nand n48559(x48559, x71997, x48554);
  nand n48560(x48560, x25790, x48557);
  nand n48561(x48561, x48560, x48559);
  nand n48562(x48562, x72002, x85417);
  nand n48563(x48563, x25796, x48561);
  nand n48564(x48564, x48563, x48562);
  nand n48565(x48565, x71977, x38874);
  nand n48566(x48566, x16876, x47775);
  nand n48567(x48567, x48566, x26557);
  nand n48568(x48568, x71977, x85267);
  nand n48569(x48569, x16876, x46498);
  nand n48570(x48570, x71977, x39880);
  nand n48571(x48571, x16876, x39880);
  nand n48572(x48572, x48571, x48570);
  nand n48573(x48573, x71977, x47019);
  nand n48574(x48574, x16876, x46973);
  nand n48575(x48575, x48574, x48573);
  nand n48576(x48576, x71977, x40691);
  nand n48577(x48577, x48566, x48576);
  nand n48578(x48578, x16876, x39119);
  nand n48579(x48579, x48578, x48576);
  nand n48580(x48580, x71977, x46854);
  nand n48581(x48581, x25749, x85418);
  nand n48582(x48582, x71982, x48567);
  nand n48583(x48583, x25749, x85419);
  nand n48584(x48584, x48583, x48582);
  nand n48585(x48585, x71982, x85420);
  nand n48586(x48586, x25749, x48572);
  nand n48587(x48587, x48586, x48585);
  nand n48588(x48588, x71982, x48575);
  nand n48589(x48589, x25749, x48577);
  nand n48590(x48590, x48589, x48588);
  nand n48591(x48591, x71982, x85419);
  nand n48592(x48592, x25749, x85420);
  nand n48593(x48593, x48592, x48591);
  nand n48594(x48594, x71982, x48572);
  nand n48595(x48595, x25749, x48575);
  nand n48596(x48596, x48595, x48594);
  nand n48597(x48597, x71982, x48579);
  nand n48598(x48598, x25749, x85421);
  nand n48599(x48599, x48598, x48597);
  nand n48600(x48600, x71987, x85422);
  nand n48601(x48601, x25772, x48584);
  nand n48602(x48602, x48601, x26594);
  nand n48603(x48603, x71987, x48587);
  nand n48604(x48604, x25772, x48590);
  nand n48605(x48605, x48604, x48603);
  nand n48606(x48606, x71987, x48593);
  nand n48607(x48607, x25772, x48596);
  nand n48608(x48608, x48607, x48606);
  nand n48609(x48609, x71987, x48599);
  nand n48610(x48610, x25782, x85423);
  nand n48611(x48611, x71992, x48602);
  nand n48612(x48612, x25782, x48605);
  nand n48613(x48613, x48612, x48611);
  nand n48614(x48614, x71992, x48608);
  nand n48615(x48615, x25782, x85424);
  nand n48616(x48616, x48615, x48614);
  nand n48617(x48617, x25790, x85425);
  nand n48618(x48618, x71997, x48613);
  nand n48619(x48619, x25790, x48616);
  nand n48620(x48620, x48619, x48618);
  nand n48621(x48621, x72002, x85426);
  nand n48622(x48622, x25796, x48620);
  nand n48623(x48623, x48622, x48621);
  nand n48624(x48624, x71977, x38876);
  nand n48625(x48625, x16876, x47778);
  nand n48626(x48626, x48625, x26620);
  nand n48627(x48627, x71977, x85268);
  nand n48628(x48628, x16876, x46503);
  nand n48629(x48629, x71977, x39885);
  nand n48630(x48630, x16876, x39885);
  nand n48631(x48631, x48630, x48629);
  nand n48632(x48632, x71977, x47021);
  nand n48633(x48633, x16876, x46974);
  nand n48634(x48634, x48633, x48632);
  nand n48635(x48635, x71977, x40802);
  nand n48636(x48636, x48625, x48635);
  nand n48637(x48637, x16876, x39125);
  nand n48638(x48638, x48637, x48635);
  nand n48639(x48639, x71977, x46858);
  nand n48640(x48640, x25749, x85427);
  nand n48641(x48641, x71982, x48626);
  nand n48642(x48642, x25749, x85428);
  nand n48643(x48643, x48642, x48641);
  nand n48644(x48644, x71982, x85429);
  nand n48645(x48645, x25749, x48631);
  nand n48646(x48646, x48645, x48644);
  nand n48647(x48647, x71982, x48634);
  nand n48648(x48648, x25749, x48636);
  nand n48649(x48649, x48648, x48647);
  nand n48650(x48650, x71982, x85428);
  nand n48651(x48651, x25749, x85429);
  nand n48652(x48652, x48651, x48650);
  nand n48653(x48653, x71982, x48631);
  nand n48654(x48654, x25749, x48634);
  nand n48655(x48655, x48654, x48653);
  nand n48656(x48656, x71982, x48638);
  nand n48657(x48657, x25749, x85430);
  nand n48658(x48658, x48657, x48656);
  nand n48659(x48659, x71987, x85431);
  nand n48660(x48660, x25772, x48643);
  nand n48661(x48661, x48660, x26657);
  nand n48662(x48662, x71987, x48646);
  nand n48663(x48663, x25772, x48649);
  nand n48664(x48664, x48663, x48662);
  nand n48665(x48665, x71987, x48652);
  nand n48666(x48666, x25772, x48655);
  nand n48667(x48667, x48666, x48665);
  nand n48668(x48668, x71987, x48658);
  nand n48669(x48669, x25782, x85432);
  nand n48670(x48670, x71992, x48661);
  nand n48671(x48671, x25782, x48664);
  nand n48672(x48672, x48671, x48670);
  nand n48673(x48673, x71992, x48667);
  nand n48674(x48674, x25782, x85433);
  nand n48675(x48675, x48674, x48673);
  nand n48676(x48676, x25790, x85434);
  nand n48677(x48677, x71997, x48672);
  nand n48678(x48678, x25790, x48675);
  nand n48679(x48679, x48678, x48677);
  nand n48680(x48680, x72002, x85435);
  nand n48681(x48681, x25796, x48679);
  nand n48682(x48682, x48681, x48680);
  nand n48683(x48683, x71977, x38878);
  nand n48684(x48684, x16876, x47781);
  nand n48685(x48685, x48684, x26683);
  nand n48686(x48686, x71977, x85269);
  nand n48687(x48687, x16876, x46508);
  nand n48688(x48688, x71977, x39890);
  nand n48689(x48689, x16876, x39890);
  nand n48690(x48690, x48689, x48688);
  nand n48691(x48691, x71977, x47023);
  nand n48692(x48692, x16876, x46975);
  nand n48693(x48693, x48692, x48691);
  nand n48694(x48694, x71977, x40922);
  nand n48695(x48695, x48684, x48694);
  nand n48696(x48696, x16876, x39131);
  nand n48697(x48697, x48696, x48694);
  nand n48698(x48698, x71977, x46862);
  nand n48699(x48699, x25749, x85436);
  nand n48700(x48700, x71982, x48685);
  nand n48701(x48701, x25749, x85437);
  nand n48702(x48702, x48701, x48700);
  nand n48703(x48703, x71982, x85438);
  nand n48704(x48704, x25749, x48690);
  nand n48705(x48705, x48704, x48703);
  nand n48706(x48706, x71982, x48693);
  nand n48707(x48707, x25749, x48695);
  nand n48708(x48708, x48707, x48706);
  nand n48709(x48709, x71982, x85437);
  nand n48710(x48710, x25749, x85438);
  nand n48711(x48711, x48710, x48709);
  nand n48712(x48712, x71982, x48690);
  nand n48713(x48713, x25749, x48693);
  nand n48714(x48714, x48713, x48712);
  nand n48715(x48715, x71982, x48697);
  nand n48716(x48716, x25749, x85439);
  nand n48717(x48717, x48716, x48715);
  nand n48718(x48718, x71987, x85440);
  nand n48719(x48719, x25772, x48702);
  nand n48720(x48720, x48719, x26720);
  nand n48721(x48721, x71987, x48705);
  nand n48722(x48722, x25772, x48708);
  nand n48723(x48723, x48722, x48721);
  nand n48724(x48724, x71987, x48711);
  nand n48725(x48725, x25772, x48714);
  nand n48726(x48726, x48725, x48724);
  nand n48727(x48727, x71987, x48717);
  nand n48728(x48728, x25782, x85441);
  nand n48729(x48729, x71992, x48720);
  nand n48730(x48730, x25782, x48723);
  nand n48731(x48731, x48730, x48729);
  nand n48732(x48732, x71992, x48726);
  nand n48733(x48733, x25782, x85442);
  nand n48734(x48734, x48733, x48732);
  nand n48735(x48735, x25790, x85443);
  nand n48736(x48736, x71997, x48731);
  nand n48737(x48737, x25790, x48734);
  nand n48738(x48738, x48737, x48736);
  nand n48739(x48739, x72002, x85444);
  nand n48740(x48740, x25796, x48738);
  nand n48741(x48741, x48740, x48739);
  nand n48742(x48742, x71977, x38880);
  nand n48743(x48743, x16876, x85285);
  nand n48744(x48744, x48743, x26746);
  nand n48745(x48745, x71977, x47397);
  nand n48746(x48746, x16876, x46512);
  nand n48747(x48747, x71977, x39895);
  nand n48748(x48748, x16876, x39895);
  nand n48749(x48749, x48748, x48747);
  nand n48750(x48750, x71977, x47025);
  nand n48751(x48751, x16876, x46976);
  nand n48752(x48752, x48751, x48750);
  nand n48753(x48753, x71977, x46929);
  nand n48754(x48754, x48743, x48753);
  nand n48755(x48755, x16876, x39137);
  nand n48756(x48756, x48755, x48753);
  nand n48757(x48757, x71977, x46866);
  nand n48758(x48758, x25749, x85445);
  nand n48759(x48759, x71982, x48744);
  nand n48760(x48760, x25749, x85446);
  nand n48761(x48761, x48760, x48759);
  nand n48762(x48762, x71982, x85447);
  nand n48763(x48763, x25749, x48749);
  nand n48764(x48764, x48763, x48762);
  nand n48765(x48765, x71982, x48752);
  nand n48766(x48766, x25749, x48754);
  nand n48767(x48767, x48766, x48765);
  nand n48768(x48768, x71982, x85446);
  nand n48769(x48769, x25749, x85447);
  nand n48770(x48770, x48769, x48768);
  nand n48771(x48771, x71982, x48749);
  nand n48772(x48772, x25749, x48752);
  nand n48773(x48773, x48772, x48771);
  nand n48774(x48774, x71982, x48756);
  nand n48775(x48775, x25749, x85448);
  nand n48776(x48776, x48775, x48774);
  nand n48777(x48777, x71987, x85449);
  nand n48778(x48778, x25772, x48761);
  nand n48779(x48779, x48778, x26783);
  nand n48780(x48780, x71987, x48764);
  nand n48781(x48781, x25772, x48767);
  nand n48782(x48782, x48781, x48780);
  nand n48783(x48783, x71987, x48770);
  nand n48784(x48784, x25772, x48773);
  nand n48785(x48785, x48784, x48783);
  nand n48786(x48786, x71987, x48776);
  nand n48787(x48787, x25782, x85450);
  nand n48788(x48788, x71992, x48779);
  nand n48789(x48789, x25782, x48782);
  nand n48790(x48790, x48789, x48788);
  nand n48791(x48791, x71992, x48785);
  nand n48792(x48792, x25782, x85451);
  nand n48793(x48793, x48792, x48791);
  nand n48794(x48794, x25790, x85452);
  nand n48795(x48795, x71997, x48790);
  nand n48796(x48796, x25790, x48793);
  nand n48797(x48797, x48796, x48795);
  nand n48798(x48798, x72002, x85453);
  nand n48799(x48799, x25796, x48797);
  nand n48800(x48800, x48799, x48798);
  nand n48801(x48801, x71977, x38882);
  nand n48802(x48802, x16876, x85286);
  nand n48803(x48803, x48802, x26809);
  nand n48804(x48804, x71977, x47400);
  nand n48805(x48805, x16876, x46516);
  nand n48806(x48806, x71977, x39900);
  nand n48807(x48807, x16876, x39900);
  nand n48808(x48808, x48807, x48806);
  nand n48809(x48809, x71977, x47027);
  nand n48810(x48810, x16876, x46977);
  nand n48811(x48811, x48810, x48809);
  nand n48812(x48812, x71977, x46931);
  nand n48813(x48813, x48802, x48812);
  nand n48814(x48814, x16876, x39143);
  nand n48815(x48815, x48814, x48812);
  nand n48816(x48816, x71977, x46870);
  nand n48817(x48817, x25749, x85454);
  nand n48818(x48818, x71982, x48803);
  nand n48819(x48819, x25749, x85455);
  nand n48820(x48820, x48819, x48818);
  nand n48821(x48821, x71982, x85456);
  nand n48822(x48822, x25749, x48808);
  nand n48823(x48823, x48822, x48821);
  nand n48824(x48824, x71982, x48811);
  nand n48825(x48825, x25749, x48813);
  nand n48826(x48826, x48825, x48824);
  nand n48827(x48827, x71982, x85455);
  nand n48828(x48828, x25749, x85456);
  nand n48829(x48829, x48828, x48827);
  nand n48830(x48830, x71982, x48808);
  nand n48831(x48831, x25749, x48811);
  nand n48832(x48832, x48831, x48830);
  nand n48833(x48833, x71982, x48815);
  nand n48834(x48834, x25749, x85457);
  nand n48835(x48835, x48834, x48833);
  nand n48836(x48836, x71987, x85458);
  nand n48837(x48837, x25772, x48820);
  nand n48838(x48838, x48837, x26846);
  nand n48839(x48839, x71987, x48823);
  nand n48840(x48840, x25772, x48826);
  nand n48841(x48841, x48840, x48839);
  nand n48842(x48842, x71987, x48829);
  nand n48843(x48843, x25772, x48832);
  nand n48844(x48844, x48843, x48842);
  nand n48845(x48845, x71987, x48835);
  nand n48846(x48846, x25782, x85459);
  nand n48847(x48847, x71992, x48838);
  nand n48848(x48848, x25782, x48841);
  nand n48849(x48849, x48848, x48847);
  nand n48850(x48850, x71992, x48844);
  nand n48851(x48851, x25782, x85460);
  nand n48852(x48852, x48851, x48850);
  nand n48853(x48853, x25790, x85461);
  nand n48854(x48854, x71997, x48849);
  nand n48855(x48855, x25790, x48852);
  nand n48856(x48856, x48855, x48854);
  nand n48857(x48857, x72002, x85462);
  nand n48858(x48858, x25796, x48856);
  nand n48859(x48859, x48858, x48857);
  nand n48860(x48860, x71977, x38884);
  nand n48861(x48861, x16876, x85287);
  nand n48862(x48862, x48861, x26872);
  nand n48863(x48863, x71977, x47403);
  nand n48864(x48864, x16876, x46520);
  nand n48865(x48865, x71977, x39905);
  nand n48866(x48866, x16876, x39905);
  nand n48867(x48867, x48866, x48865);
  nand n48868(x48868, x71977, x47029);
  nand n48869(x48869, x16876, x46978);
  nand n48870(x48870, x48869, x48868);
  nand n48871(x48871, x71977, x46933);
  nand n48872(x48872, x48861, x48871);
  nand n48873(x48873, x16876, x39149);
  nand n48874(x48874, x48873, x48871);
  nand n48875(x48875, x71977, x46874);
  nand n48876(x48876, x25749, x85463);
  nand n48877(x48877, x71982, x48862);
  nand n48878(x48878, x25749, x85464);
  nand n48879(x48879, x48878, x48877);
  nand n48880(x48880, x71982, x85465);
  nand n48881(x48881, x25749, x48867);
  nand n48882(x48882, x48881, x48880);
  nand n48883(x48883, x71982, x48870);
  nand n48884(x48884, x25749, x48872);
  nand n48885(x48885, x48884, x48883);
  nand n48886(x48886, x71982, x85464);
  nand n48887(x48887, x25749, x85465);
  nand n48888(x48888, x48887, x48886);
  nand n48889(x48889, x71982, x48867);
  nand n48890(x48890, x25749, x48870);
  nand n48891(x48891, x48890, x48889);
  nand n48892(x48892, x71982, x48874);
  nand n48893(x48893, x25749, x85466);
  nand n48894(x48894, x48893, x48892);
  nand n48895(x48895, x71987, x85467);
  nand n48896(x48896, x25772, x48879);
  nand n48897(x48897, x48896, x26909);
  nand n48898(x48898, x71987, x48882);
  nand n48899(x48899, x25772, x48885);
  nand n48900(x48900, x48899, x48898);
  nand n48901(x48901, x71987, x48888);
  nand n48902(x48902, x25772, x48891);
  nand n48903(x48903, x48902, x48901);
  nand n48904(x48904, x71987, x48894);
  nand n48905(x48905, x25782, x85468);
  nand n48906(x48906, x71992, x48897);
  nand n48907(x48907, x25782, x48900);
  nand n48908(x48908, x48907, x48906);
  nand n48909(x48909, x71992, x48903);
  nand n48910(x48910, x25782, x85469);
  nand n48911(x48911, x48910, x48909);
  nand n48912(x48912, x25790, x85470);
  nand n48913(x48913, x71997, x48908);
  nand n48914(x48914, x25790, x48911);
  nand n48915(x48915, x48914, x48913);
  nand n48916(x48916, x72002, x85471);
  nand n48917(x48917, x25796, x48915);
  nand n48918(x48918, x48917, x48916);
  nand n48919(x48919, x71977, x38886);
  nand n48920(x48920, x16876, x85288);
  nand n48921(x48921, x48920, x26935);
  nand n48922(x48922, x71977, x47406);
  nand n48923(x48923, x16876, x46524);
  nand n48924(x48924, x71977, x39910);
  nand n48925(x48925, x16876, x39910);
  nand n48926(x48926, x48925, x48924);
  nand n48927(x48927, x71977, x47031);
  nand n48928(x48928, x16876, x46979);
  nand n48929(x48929, x48928, x48927);
  nand n48930(x48930, x71977, x46935);
  nand n48931(x48931, x48920, x48930);
  nand n48932(x48932, x16876, x39155);
  nand n48933(x48933, x48932, x48930);
  nand n48934(x48934, x71977, x46878);
  nand n48935(x48935, x25749, x85472);
  nand n48936(x48936, x71982, x48921);
  nand n48937(x48937, x25749, x85473);
  nand n48938(x48938, x48937, x48936);
  nand n48939(x48939, x71982, x85474);
  nand n48940(x48940, x25749, x48926);
  nand n48941(x48941, x48940, x48939);
  nand n48942(x48942, x71982, x48929);
  nand n48943(x48943, x25749, x48931);
  nand n48944(x48944, x48943, x48942);
  nand n48945(x48945, x71982, x85473);
  nand n48946(x48946, x25749, x85474);
  nand n48947(x48947, x48946, x48945);
  nand n48948(x48948, x71982, x48926);
  nand n48949(x48949, x25749, x48929);
  nand n48950(x48950, x48949, x48948);
  nand n48951(x48951, x71982, x48933);
  nand n48952(x48952, x25749, x85475);
  nand n48953(x48953, x48952, x48951);
  nand n48954(x48954, x71987, x85476);
  nand n48955(x48955, x25772, x48938);
  nand n48956(x48956, x48955, x26972);
  nand n48957(x48957, x71987, x48941);
  nand n48958(x48958, x25772, x48944);
  nand n48959(x48959, x48958, x48957);
  nand n48960(x48960, x71987, x48947);
  nand n48961(x48961, x25772, x48950);
  nand n48962(x48962, x48961, x48960);
  nand n48963(x48963, x71987, x48953);
  nand n48964(x48964, x25782, x85477);
  nand n48965(x48965, x71992, x48956);
  nand n48966(x48966, x25782, x48959);
  nand n48967(x48967, x48966, x48965);
  nand n48968(x48968, x71992, x48962);
  nand n48969(x48969, x25782, x85478);
  nand n48970(x48970, x48969, x48968);
  nand n48971(x48971, x25790, x85479);
  nand n48972(x48972, x71997, x48967);
  nand n48973(x48973, x25790, x48970);
  nand n48974(x48974, x48973, x48972);
  nand n48975(x48975, x72002, x85480);
  nand n48976(x48976, x25796, x48974);
  nand n48977(x48977, x48976, x48975);
  nand n48978(x48978, x71977, x38888);
  nand n48979(x48979, x16876, x85289);
  nand n48980(x48980, x48979, x26998);
  nand n48981(x48981, x71977, x47409);
  nand n48982(x48982, x16876, x46528);
  nand n48983(x48983, x71977, x39915);
  nand n48984(x48984, x16876, x39915);
  nand n48985(x48985, x48984, x48983);
  nand n48986(x48986, x71977, x47033);
  nand n48987(x48987, x16876, x46980);
  nand n48988(x48988, x48987, x48986);
  nand n48989(x48989, x71977, x46937);
  nand n48990(x48990, x48979, x48989);
  nand n48991(x48991, x16876, x39161);
  nand n48992(x48992, x48991, x48989);
  nand n48993(x48993, x71977, x46882);
  nand n48994(x48994, x25749, x85481);
  nand n48995(x48995, x71982, x48980);
  nand n48996(x48996, x25749, x85482);
  nand n48997(x48997, x48996, x48995);
  nand n48998(x48998, x71982, x85483);
  nand n48999(x48999, x25749, x48985);
  nand n49000(x49000, x48999, x48998);
  nand n49001(x49001, x71982, x48988);
  nand n49002(x49002, x25749, x48990);
  nand n49003(x49003, x49002, x49001);
  nand n49004(x49004, x71982, x85482);
  nand n49005(x49005, x25749, x85483);
  nand n49006(x49006, x49005, x49004);
  nand n49007(x49007, x71982, x48985);
  nand n49008(x49008, x25749, x48988);
  nand n49009(x49009, x49008, x49007);
  nand n49010(x49010, x71982, x48992);
  nand n49011(x49011, x25749, x85484);
  nand n49012(x49012, x49011, x49010);
  nand n49013(x49013, x71987, x85485);
  nand n49014(x49014, x25772, x48997);
  nand n49015(x49015, x49014, x27035);
  nand n49016(x49016, x71987, x49000);
  nand n49017(x49017, x25772, x49003);
  nand n49018(x49018, x49017, x49016);
  nand n49019(x49019, x71987, x49006);
  nand n49020(x49020, x25772, x49009);
  nand n49021(x49021, x49020, x49019);
  nand n49022(x49022, x71987, x49012);
  nand n49023(x49023, x25782, x85486);
  nand n49024(x49024, x71992, x49015);
  nand n49025(x49025, x25782, x49018);
  nand n49026(x49026, x49025, x49024);
  nand n49027(x49027, x71992, x49021);
  nand n49028(x49028, x25782, x85487);
  nand n49029(x49029, x49028, x49027);
  nand n49030(x49030, x25790, x85488);
  nand n49031(x49031, x71997, x49026);
  nand n49032(x49032, x25790, x49029);
  nand n49033(x49033, x49032, x49031);
  nand n49034(x49034, x72002, x85489);
  nand n49035(x49035, x25796, x49033);
  nand n49036(x49036, x49035, x49034);
  nand n49037(x49037, x71977, x38890);
  nand n49038(x49038, x16876, x85290);
  nand n49039(x49039, x49038, x27061);
  nand n49040(x49040, x71977, x47412);
  nand n49041(x49041, x16876, x46532);
  nand n49042(x49042, x71977, x39920);
  nand n49043(x49043, x16876, x39920);
  nand n49044(x49044, x49043, x49042);
  nand n49045(x49045, x71977, x47035);
  nand n49046(x49046, x16876, x46981);
  nand n49047(x49047, x49046, x49045);
  nand n49048(x49048, x71977, x46939);
  nand n49049(x49049, x49038, x49048);
  nand n49050(x49050, x16876, x39167);
  nand n49051(x49051, x49050, x49048);
  nand n49052(x49052, x71977, x46886);
  nand n49053(x49053, x25749, x85490);
  nand n49054(x49054, x71982, x49039);
  nand n49055(x49055, x25749, x85491);
  nand n49056(x49056, x49055, x49054);
  nand n49057(x49057, x71982, x85492);
  nand n49058(x49058, x25749, x49044);
  nand n49059(x49059, x49058, x49057);
  nand n49060(x49060, x71982, x49047);
  nand n49061(x49061, x25749, x49049);
  nand n49062(x49062, x49061, x49060);
  nand n49063(x49063, x71982, x85491);
  nand n49064(x49064, x25749, x85492);
  nand n49065(x49065, x49064, x49063);
  nand n49066(x49066, x71982, x49044);
  nand n49067(x49067, x25749, x49047);
  nand n49068(x49068, x49067, x49066);
  nand n49069(x49069, x71982, x49051);
  nand n49070(x49070, x25749, x85493);
  nand n49071(x49071, x49070, x49069);
  nand n49072(x49072, x71987, x85494);
  nand n49073(x49073, x25772, x49056);
  nand n49074(x49074, x49073, x27098);
  nand n49075(x49075, x71987, x49059);
  nand n49076(x49076, x25772, x49062);
  nand n49077(x49077, x49076, x49075);
  nand n49078(x49078, x71987, x49065);
  nand n49079(x49079, x25772, x49068);
  nand n49080(x49080, x49079, x49078);
  nand n49081(x49081, x71987, x49071);
  nand n49082(x49082, x25782, x85495);
  nand n49083(x49083, x71992, x49074);
  nand n49084(x49084, x25782, x49077);
  nand n49085(x49085, x49084, x49083);
  nand n49086(x49086, x71992, x49080);
  nand n49087(x49087, x25782, x85496);
  nand n49088(x49088, x49087, x49086);
  nand n49089(x49089, x25790, x85497);
  nand n49090(x49090, x71997, x49085);
  nand n49091(x49091, x25790, x49088);
  nand n49092(x49092, x49091, x49090);
  nand n49093(x49093, x72002, x85498);
  nand n49094(x49094, x25796, x49092);
  nand n49095(x49095, x49094, x49093);
  nand n49096(x49096, x71977, x38892);
  nand n49097(x49097, x16876, x85291);
  nand n49098(x49098, x49097, x27124);
  nand n49099(x49099, x71977, x47415);
  nand n49100(x49100, x16876, x46537);
  nand n49101(x49101, x71977, x39925);
  nand n49102(x49102, x16876, x39925);
  nand n49103(x49103, x49102, x49101);
  nand n49104(x49104, x71977, x47037);
  nand n49105(x49105, x16876, x46982);
  nand n49106(x49106, x49105, x49104);
  nand n49107(x49107, x71977, x46941);
  nand n49108(x49108, x49097, x49107);
  nand n49109(x49109, x16876, x39173);
  nand n49110(x49110, x49109, x49107);
  nand n49111(x49111, x71977, x46890);
  nand n49112(x49112, x25749, x85499);
  nand n49113(x49113, x71982, x49098);
  nand n49114(x49114, x25749, x85500);
  nand n49115(x49115, x49114, x49113);
  nand n49116(x49116, x71982, x85501);
  nand n49117(x49117, x25749, x49103);
  nand n49118(x49118, x49117, x49116);
  nand n49119(x49119, x71982, x49106);
  nand n49120(x49120, x25749, x49108);
  nand n49121(x49121, x49120, x49119);
  nand n49122(x49122, x71982, x85500);
  nand n49123(x49123, x25749, x85501);
  nand n49124(x49124, x49123, x49122);
  nand n49125(x49125, x71982, x49103);
  nand n49126(x49126, x25749, x49106);
  nand n49127(x49127, x49126, x49125);
  nand n49128(x49128, x71982, x49110);
  nand n49129(x49129, x25749, x85502);
  nand n49130(x49130, x49129, x49128);
  nand n49131(x49131, x71987, x85503);
  nand n49132(x49132, x25772, x49115);
  nand n49133(x49133, x49132, x27161);
  nand n49134(x49134, x71987, x49118);
  nand n49135(x49135, x25772, x49121);
  nand n49136(x49136, x49135, x49134);
  nand n49137(x49137, x71987, x49124);
  nand n49138(x49138, x25772, x49127);
  nand n49139(x49139, x49138, x49137);
  nand n49140(x49140, x71987, x49130);
  nand n49141(x49141, x25782, x85504);
  nand n49142(x49142, x71992, x49133);
  nand n49143(x49143, x25782, x49136);
  nand n49144(x49144, x49143, x49142);
  nand n49145(x49145, x71992, x49139);
  nand n49146(x49146, x25782, x85505);
  nand n49147(x49147, x49146, x49145);
  nand n49148(x49148, x25790, x85506);
  nand n49149(x49149, x71997, x49144);
  nand n49150(x49150, x25790, x49147);
  nand n49151(x49151, x49150, x49149);
  nand n49152(x49152, x72002, x85507);
  nand n49153(x49153, x25796, x49151);
  nand n49154(x49154, x49153, x49152);
  nand n49155(x49155, x71977, x38894);
  nand n49156(x49156, x16876, x85292);
  nand n49157(x49157, x49156, x27187);
  nand n49158(x49158, x71977, x47418);
  nand n49159(x49159, x16876, x46542);
  nand n49160(x49160, x71977, x39930);
  nand n49161(x49161, x16876, x39930);
  nand n49162(x49162, x49161, x49160);
  nand n49163(x49163, x71977, x47039);
  nand n49164(x49164, x16876, x46983);
  nand n49165(x49165, x49164, x49163);
  nand n49166(x49166, x71977, x46943);
  nand n49167(x49167, x49156, x49166);
  nand n49168(x49168, x16876, x39179);
  nand n49169(x49169, x49168, x49166);
  nand n49170(x49170, x71977, x46894);
  nand n49171(x49171, x25749, x85508);
  nand n49172(x49172, x71982, x49157);
  nand n49173(x49173, x25749, x85509);
  nand n49174(x49174, x49173, x49172);
  nand n49175(x49175, x71982, x85510);
  nand n49176(x49176, x25749, x49162);
  nand n49177(x49177, x49176, x49175);
  nand n49178(x49178, x71982, x49165);
  nand n49179(x49179, x25749, x49167);
  nand n49180(x49180, x49179, x49178);
  nand n49181(x49181, x71982, x85509);
  nand n49182(x49182, x25749, x85510);
  nand n49183(x49183, x49182, x49181);
  nand n49184(x49184, x71982, x49162);
  nand n49185(x49185, x25749, x49165);
  nand n49186(x49186, x49185, x49184);
  nand n49187(x49187, x71982, x49169);
  nand n49188(x49188, x25749, x85511);
  nand n49189(x49189, x49188, x49187);
  nand n49190(x49190, x71987, x85512);
  nand n49191(x49191, x25772, x49174);
  nand n49192(x49192, x49191, x27224);
  nand n49193(x49193, x71987, x49177);
  nand n49194(x49194, x25772, x49180);
  nand n49195(x49195, x49194, x49193);
  nand n49196(x49196, x71987, x49183);
  nand n49197(x49197, x25772, x49186);
  nand n49198(x49198, x49197, x49196);
  nand n49199(x49199, x71987, x49189);
  nand n49200(x49200, x25782, x85513);
  nand n49201(x49201, x71992, x49192);
  nand n49202(x49202, x25782, x49195);
  nand n49203(x49203, x49202, x49201);
  nand n49204(x49204, x71992, x49198);
  nand n49205(x49205, x25782, x85514);
  nand n49206(x49206, x49205, x49204);
  nand n49207(x49207, x25790, x85515);
  nand n49208(x49208, x71997, x49203);
  nand n49209(x49209, x25790, x49206);
  nand n49210(x49210, x49209, x49208);
  nand n49211(x49211, x72002, x85516);
  nand n49212(x49212, x25796, x49210);
  nand n49213(x49213, x49212, x49211);
  nand n49214(x49214, x71977, x38896);
  nand n49215(x49215, x16876, x85293);
  nand n49216(x49216, x49215, x27250);
  nand n49217(x49217, x71977, x47421);
  nand n49218(x49218, x16876, x46547);
  nand n49219(x49219, x71977, x39935);
  nand n49220(x49220, x16876, x39935);
  nand n49221(x49221, x49220, x49219);
  nand n49222(x49222, x71977, x47041);
  nand n49223(x49223, x16876, x46984);
  nand n49224(x49224, x49223, x49222);
  nand n49225(x49225, x71977, x46945);
  nand n49226(x49226, x49215, x49225);
  nand n49227(x49227, x16876, x39185);
  nand n49228(x49228, x49227, x49225);
  nand n49229(x49229, x71977, x46898);
  nand n49230(x49230, x25749, x85517);
  nand n49231(x49231, x71982, x49216);
  nand n49232(x49232, x25749, x85518);
  nand n49233(x49233, x49232, x49231);
  nand n49234(x49234, x71982, x85519);
  nand n49235(x49235, x25749, x49221);
  nand n49236(x49236, x49235, x49234);
  nand n49237(x49237, x71982, x49224);
  nand n49238(x49238, x25749, x49226);
  nand n49239(x49239, x49238, x49237);
  nand n49240(x49240, x71982, x85518);
  nand n49241(x49241, x25749, x85519);
  nand n49242(x49242, x49241, x49240);
  nand n49243(x49243, x71982, x49221);
  nand n49244(x49244, x25749, x49224);
  nand n49245(x49245, x49244, x49243);
  nand n49246(x49246, x71982, x49228);
  nand n49247(x49247, x25749, x85520);
  nand n49248(x49248, x49247, x49246);
  nand n49249(x49249, x71987, x85521);
  nand n49250(x49250, x25772, x49233);
  nand n49251(x49251, x49250, x27287);
  nand n49252(x49252, x71987, x49236);
  nand n49253(x49253, x25772, x49239);
  nand n49254(x49254, x49253, x49252);
  nand n49255(x49255, x71987, x49242);
  nand n49256(x49256, x25772, x49245);
  nand n49257(x49257, x49256, x49255);
  nand n49258(x49258, x71987, x49248);
  nand n49259(x49259, x25782, x85522);
  nand n49260(x49260, x71992, x49251);
  nand n49261(x49261, x25782, x49254);
  nand n49262(x49262, x49261, x49260);
  nand n49263(x49263, x71992, x49257);
  nand n49264(x49264, x25782, x85523);
  nand n49265(x49265, x49264, x49263);
  nand n49266(x49266, x25790, x85524);
  nand n49267(x49267, x71997, x49262);
  nand n49268(x49268, x25790, x49265);
  nand n49269(x49269, x49268, x49267);
  nand n49270(x49270, x72002, x85525);
  nand n49271(x49271, x25796, x49269);
  nand n49272(x49272, x49271, x49270);
  nand n49273(x49273, x71977, x38898);
  nand n49274(x49274, x16876, x85294);
  nand n49275(x49275, x49274, x27313);
  nand n49276(x49276, x71977, x47424);
  nand n49277(x49277, x16876, x46552);
  nand n49278(x49278, x71977, x39940);
  nand n49279(x49279, x16876, x39940);
  nand n49280(x49280, x49279, x49278);
  nand n49281(x49281, x71977, x47043);
  nand n49282(x49282, x16876, x46985);
  nand n49283(x49283, x49282, x49281);
  nand n49284(x49284, x71977, x46947);
  nand n49285(x49285, x49274, x49284);
  nand n49286(x49286, x16876, x39191);
  nand n49287(x49287, x49286, x49284);
  nand n49288(x49288, x71977, x46902);
  nand n49289(x49289, x25749, x85526);
  nand n49290(x49290, x71982, x49275);
  nand n49291(x49291, x25749, x85527);
  nand n49292(x49292, x49291, x49290);
  nand n49293(x49293, x71982, x85528);
  nand n49294(x49294, x25749, x49280);
  nand n49295(x49295, x49294, x49293);
  nand n49296(x49296, x71982, x49283);
  nand n49297(x49297, x25749, x49285);
  nand n49298(x49298, x49297, x49296);
  nand n49299(x49299, x71982, x85527);
  nand n49300(x49300, x25749, x85528);
  nand n49301(x49301, x49300, x49299);
  nand n49302(x49302, x71982, x49280);
  nand n49303(x49303, x25749, x49283);
  nand n49304(x49304, x49303, x49302);
  nand n49305(x49305, x71982, x49287);
  nand n49306(x49306, x25749, x85529);
  nand n49307(x49307, x49306, x49305);
  nand n49308(x49308, x71987, x85530);
  nand n49309(x49309, x25772, x49292);
  nand n49310(x49310, x49309, x27350);
  nand n49311(x49311, x71987, x49295);
  nand n49312(x49312, x25772, x49298);
  nand n49313(x49313, x49312, x49311);
  nand n49314(x49314, x71987, x49301);
  nand n49315(x49315, x25772, x49304);
  nand n49316(x49316, x49315, x49314);
  nand n49317(x49317, x71987, x49307);
  nand n49318(x49318, x25782, x85531);
  nand n49319(x49319, x71992, x49310);
  nand n49320(x49320, x25782, x49313);
  nand n49321(x49321, x49320, x49319);
  nand n49322(x49322, x71992, x49316);
  nand n49323(x49323, x25782, x85532);
  nand n49324(x49324, x49323, x49322);
  nand n49325(x49325, x25790, x85533);
  nand n49326(x49326, x71997, x49321);
  nand n49327(x49327, x25790, x49324);
  nand n49328(x49328, x49327, x49326);
  nand n49329(x49329, x72002, x85534);
  nand n49330(x49330, x25796, x49328);
  nand n49331(x49331, x49330, x49329);
  nand n49332(x49332, x71977, x38900);
  nand n49333(x49333, x16876, x85295);
  nand n49334(x49334, x49333, x27376);
  nand n49335(x49335, x71977, x47427);
  nand n49336(x49336, x16876, x46557);
  nand n49337(x49337, x71977, x39945);
  nand n49338(x49338, x16876, x39945);
  nand n49339(x49339, x49338, x49337);
  nand n49340(x49340, x71977, x47045);
  nand n49341(x49341, x16876, x46986);
  nand n49342(x49342, x49341, x49340);
  nand n49343(x49343, x71977, x46949);
  nand n49344(x49344, x49333, x49343);
  nand n49345(x49345, x16876, x39197);
  nand n49346(x49346, x49345, x49343);
  nand n49347(x49347, x71977, x46906);
  nand n49348(x49348, x25749, x85535);
  nand n49349(x49349, x71982, x49334);
  nand n49350(x49350, x25749, x85536);
  nand n49351(x49351, x49350, x49349);
  nand n49352(x49352, x71982, x85537);
  nand n49353(x49353, x25749, x49339);
  nand n49354(x49354, x49353, x49352);
  nand n49355(x49355, x71982, x49342);
  nand n49356(x49356, x25749, x49344);
  nand n49357(x49357, x49356, x49355);
  nand n49358(x49358, x71982, x85536);
  nand n49359(x49359, x25749, x85537);
  nand n49360(x49360, x49359, x49358);
  nand n49361(x49361, x71982, x49339);
  nand n49362(x49362, x25749, x49342);
  nand n49363(x49363, x49362, x49361);
  nand n49364(x49364, x71982, x49346);
  nand n49365(x49365, x25749, x85538);
  nand n49366(x49366, x49365, x49364);
  nand n49367(x49367, x71987, x85539);
  nand n49368(x49368, x25772, x49351);
  nand n49369(x49369, x49368, x27413);
  nand n49370(x49370, x71987, x49354);
  nand n49371(x49371, x25772, x49357);
  nand n49372(x49372, x49371, x49370);
  nand n49373(x49373, x71987, x49360);
  nand n49374(x49374, x25772, x49363);
  nand n49375(x49375, x49374, x49373);
  nand n49376(x49376, x71987, x49366);
  nand n49377(x49377, x25782, x85540);
  nand n49378(x49378, x71992, x49369);
  nand n49379(x49379, x25782, x49372);
  nand n49380(x49380, x49379, x49378);
  nand n49381(x49381, x71992, x49375);
  nand n49382(x49382, x25782, x85541);
  nand n49383(x49383, x49382, x49381);
  nand n49384(x49384, x25790, x85542);
  nand n49385(x49385, x71997, x49380);
  nand n49386(x49386, x25790, x49383);
  nand n49387(x49387, x49386, x49385);
  nand n49388(x49388, x72002, x85543);
  nand n49389(x49389, x25796, x49387);
  nand n49390(x49390, x49389, x49388);
  nand n49391(x49391, x71977, x38902);
  nand n49392(x49392, x16876, x85296);
  nand n49393(x49393, x49392, x27439);
  nand n49394(x49394, x71977, x47430);
  nand n49395(x49395, x16876, x46562);
  nand n49396(x49396, x71977, x39950);
  nand n49397(x49397, x16876, x39950);
  nand n49398(x49398, x49397, x49396);
  nand n49399(x49399, x71977, x47047);
  nand n49400(x49400, x16876, x46987);
  nand n49401(x49401, x49400, x49399);
  nand n49402(x49402, x71977, x46951);
  nand n49403(x49403, x49392, x49402);
  nand n49404(x49404, x16876, x39203);
  nand n49405(x49405, x49404, x49402);
  nand n49406(x49406, x71977, x46910);
  nand n49407(x49407, x25749, x85544);
  nand n49408(x49408, x71982, x49393);
  nand n49409(x49409, x25749, x85545);
  nand n49410(x49410, x49409, x49408);
  nand n49411(x49411, x71982, x85546);
  nand n49412(x49412, x25749, x49398);
  nand n49413(x49413, x49412, x49411);
  nand n49414(x49414, x71982, x49401);
  nand n49415(x49415, x25749, x49403);
  nand n49416(x49416, x49415, x49414);
  nand n49417(x49417, x71982, x85545);
  nand n49418(x49418, x25749, x85546);
  nand n49419(x49419, x49418, x49417);
  nand n49420(x49420, x71982, x49398);
  nand n49421(x49421, x25749, x49401);
  nand n49422(x49422, x49421, x49420);
  nand n49423(x49423, x71982, x49405);
  nand n49424(x49424, x25749, x85547);
  nand n49425(x49425, x49424, x49423);
  nand n49426(x49426, x71987, x85548);
  nand n49427(x49427, x25772, x49410);
  nand n49428(x49428, x49427, x27476);
  nand n49429(x49429, x71987, x49413);
  nand n49430(x49430, x25772, x49416);
  nand n49431(x49431, x49430, x49429);
  nand n49432(x49432, x71987, x49419);
  nand n49433(x49433, x25772, x49422);
  nand n49434(x49434, x49433, x49432);
  nand n49435(x49435, x71987, x49425);
  nand n49436(x49436, x25782, x85549);
  nand n49437(x49437, x71992, x49428);
  nand n49438(x49438, x25782, x49431);
  nand n49439(x49439, x49438, x49437);
  nand n49440(x49440, x71992, x49434);
  nand n49441(x49441, x25782, x85550);
  nand n49442(x49442, x49441, x49440);
  nand n49443(x49443, x25790, x85551);
  nand n49444(x49444, x71997, x49439);
  nand n49445(x49445, x25790, x49442);
  nand n49446(x49446, x49445, x49444);
  nand n49447(x49447, x72002, x85552);
  nand n49448(x49448, x25796, x49446);
  nand n49449(x49449, x49448, x49447);
  nand n49450(x49450, x71977, x38904);
  nand n49451(x49451, x16876, x85297);
  nand n49452(x49452, x49451, x27502);
  nand n49453(x49453, x71977, x47433);
  nand n49454(x49454, x16876, x46567);
  nand n49455(x49455, x71977, x39955);
  nand n49456(x49456, x16876, x39955);
  nand n49457(x49457, x49456, x49455);
  nand n49458(x49458, x71977, x47049);
  nand n49459(x49459, x16876, x46988);
  nand n49460(x49460, x49459, x49458);
  nand n49461(x49461, x71977, x46953);
  nand n49462(x49462, x49451, x49461);
  nand n49463(x49463, x16876, x39209);
  nand n49464(x49464, x49463, x49461);
  nand n49465(x49465, x71977, x46914);
  nand n49466(x49466, x25749, x85553);
  nand n49467(x49467, x71982, x49452);
  nand n49468(x49468, x25749, x85554);
  nand n49469(x49469, x49468, x49467);
  nand n49470(x49470, x71982, x85555);
  nand n49471(x49471, x25749, x49457);
  nand n49472(x49472, x49471, x49470);
  nand n49473(x49473, x71982, x49460);
  nand n49474(x49474, x25749, x49462);
  nand n49475(x49475, x49474, x49473);
  nand n49476(x49476, x71982, x85554);
  nand n49477(x49477, x25749, x85555);
  nand n49478(x49478, x49477, x49476);
  nand n49479(x49479, x71982, x49457);
  nand n49480(x49480, x25749, x49460);
  nand n49481(x49481, x49480, x49479);
  nand n49482(x49482, x71982, x49464);
  nand n49483(x49483, x25749, x85556);
  nand n49484(x49484, x49483, x49482);
  nand n49485(x49485, x71987, x85557);
  nand n49486(x49486, x25772, x49469);
  nand n49487(x49487, x49486, x27539);
  nand n49488(x49488, x71987, x49472);
  nand n49489(x49489, x25772, x49475);
  nand n49490(x49490, x49489, x49488);
  nand n49491(x49491, x71987, x49478);
  nand n49492(x49492, x25772, x49481);
  nand n49493(x49493, x49492, x49491);
  nand n49494(x49494, x71987, x49484);
  nand n49495(x49495, x25782, x85558);
  nand n49496(x49496, x71992, x49487);
  nand n49497(x49497, x25782, x49490);
  nand n49498(x49498, x49497, x49496);
  nand n49499(x49499, x71992, x49493);
  nand n49500(x49500, x25782, x85559);
  nand n49501(x49501, x49500, x49499);
  nand n49502(x49502, x25790, x85560);
  nand n49503(x49503, x71997, x49498);
  nand n49504(x49504, x25790, x49501);
  nand n49505(x49505, x49504, x49503);
  nand n49506(x49506, x72002, x85561);
  nand n49507(x49507, x25796, x49505);
  nand n49508(x49508, x49507, x49506);
  nand n49509(x49509, x71977, x38906);
  nand n49510(x49510, x16876, x85298);
  nand n49511(x49511, x49510, x27565);
  nand n49512(x49512, x71977, x47436);
  nand n49513(x49513, x16876, x46572);
  nand n49514(x49514, x71977, x39960);
  nand n49515(x49515, x16876, x39960);
  nand n49516(x49516, x49515, x49514);
  nand n49517(x49517, x71977, x47051);
  nand n49518(x49518, x16876, x46989);
  nand n49519(x49519, x49518, x49517);
  nand n49520(x49520, x71977, x46955);
  nand n49521(x49521, x49510, x49520);
  nand n49522(x49522, x16876, x39215);
  nand n49523(x49523, x49522, x49520);
  nand n49524(x49524, x71977, x46918);
  nand n49525(x49525, x25749, x85562);
  nand n49526(x49526, x71982, x49511);
  nand n49527(x49527, x25749, x85563);
  nand n49528(x49528, x49527, x49526);
  nand n49529(x49529, x71982, x85564);
  nand n49530(x49530, x25749, x49516);
  nand n49531(x49531, x49530, x49529);
  nand n49532(x49532, x71982, x49519);
  nand n49533(x49533, x25749, x49521);
  nand n49534(x49534, x49533, x49532);
  nand n49535(x49535, x71982, x85563);
  nand n49536(x49536, x25749, x85564);
  nand n49537(x49537, x49536, x49535);
  nand n49538(x49538, x71982, x49516);
  nand n49539(x49539, x25749, x49519);
  nand n49540(x49540, x49539, x49538);
  nand n49541(x49541, x71982, x49523);
  nand n49542(x49542, x25749, x85565);
  nand n49543(x49543, x49542, x49541);
  nand n49544(x49544, x71987, x85566);
  nand n49545(x49545, x25772, x49528);
  nand n49546(x49546, x49545, x27602);
  nand n49547(x49547, x71987, x49531);
  nand n49548(x49548, x25772, x49534);
  nand n49549(x49549, x49548, x49547);
  nand n49550(x49550, x71987, x49537);
  nand n49551(x49551, x25772, x49540);
  nand n49552(x49552, x49551, x49550);
  nand n49553(x49553, x71987, x49543);
  nand n49554(x49554, x25782, x85567);
  nand n49555(x49555, x71992, x49546);
  nand n49556(x49556, x25782, x49549);
  nand n49557(x49557, x49556, x49555);
  nand n49558(x49558, x71992, x49552);
  nand n49559(x49559, x25782, x85568);
  nand n49560(x49560, x49559, x49558);
  nand n49561(x49561, x25790, x85569);
  nand n49562(x49562, x71997, x49557);
  nand n49563(x49563, x25790, x49560);
  nand n49564(x49564, x49563, x49562);
  nand n49565(x49565, x72002, x85570);
  nand n49566(x49566, x25796, x49564);
  nand n49567(x49567, x49566, x49565);
  nand n49568(x49568, x71977, x38908);
  nand n49569(x49569, x16876, x85299);
  nand n49570(x49570, x49569, x27628);
  nand n49571(x49571, x71977, x47439);
  nand n49572(x49572, x16876, x46577);
  nand n49573(x49573, x71977, x39965);
  nand n49574(x49574, x16876, x39965);
  nand n49575(x49575, x49574, x49573);
  nand n49576(x49576, x71977, x47053);
  nand n49577(x49577, x16876, x46990);
  nand n49578(x49578, x49577, x49576);
  nand n49579(x49579, x71977, x46957);
  nand n49580(x49580, x49569, x49579);
  nand n49581(x49581, x16876, x39221);
  nand n49582(x49582, x49581, x49579);
  nand n49583(x49583, x71977, x46922);
  nand n49584(x49584, x25749, x85571);
  nand n49585(x49585, x71982, x49570);
  nand n49586(x49586, x25749, x85572);
  nand n49587(x49587, x49586, x49585);
  nand n49588(x49588, x71982, x85573);
  nand n49589(x49589, x25749, x49575);
  nand n49590(x49590, x49589, x49588);
  nand n49591(x49591, x71982, x49578);
  nand n49592(x49592, x25749, x49580);
  nand n49593(x49593, x49592, x49591);
  nand n49594(x49594, x71982, x85572);
  nand n49595(x49595, x25749, x85573);
  nand n49596(x49596, x49595, x49594);
  nand n49597(x49597, x71982, x49575);
  nand n49598(x49598, x25749, x49578);
  nand n49599(x49599, x49598, x49597);
  nand n49600(x49600, x71982, x49582);
  nand n49601(x49601, x25749, x85574);
  nand n49602(x49602, x49601, x49600);
  nand n49603(x49603, x71987, x85575);
  nand n49604(x49604, x25772, x49587);
  nand n49605(x49605, x49604, x27665);
  nand n49606(x49606, x71987, x49590);
  nand n49607(x49607, x25772, x49593);
  nand n49608(x49608, x49607, x49606);
  nand n49609(x49609, x71987, x49596);
  nand n49610(x49610, x25772, x49599);
  nand n49611(x49611, x49610, x49609);
  nand n49612(x49612, x71987, x49602);
  nand n49613(x49613, x25782, x85576);
  nand n49614(x49614, x71992, x49605);
  nand n49615(x49615, x25782, x49608);
  nand n49616(x49616, x49615, x49614);
  nand n49617(x49617, x71992, x49611);
  nand n49618(x49618, x25782, x85577);
  nand n49619(x49619, x49618, x49617);
  nand n49620(x49620, x25790, x85578);
  nand n49621(x49621, x71997, x49616);
  nand n49622(x49622, x25790, x49619);
  nand n49623(x49623, x49622, x49621);
  nand n49624(x49624, x72002, x85579);
  nand n49625(x49625, x25796, x49623);
  nand n49626(x49626, x49625, x49624);
  nand n49627(x49627, x71977, x38910);
  nand n49628(x49628, x16876, x85300);
  nand n49629(x49629, x49628, x27691);
  nand n49630(x49630, x71977, x47442);
  nand n49631(x49631, x16876, x46582);
  nand n49632(x49632, x71977, x39970);
  nand n49633(x49633, x16876, x39970);
  nand n49634(x49634, x49633, x49632);
  nand n49635(x49635, x71977, x47055);
  nand n49636(x49636, x16876, x46991);
  nand n49637(x49637, x49636, x49635);
  nand n49638(x49638, x71977, x46959);
  nand n49639(x49639, x49628, x49638);
  nand n49640(x49640, x16876, x39227);
  nand n49641(x49641, x49640, x49638);
  nand n49642(x49642, x71977, x46926);
  nand n49643(x49643, x25749, x85580);
  nand n49644(x49644, x71982, x49629);
  nand n49645(x49645, x25749, x85581);
  nand n49646(x49646, x49645, x49644);
  nand n49647(x49647, x71982, x85582);
  nand n49648(x49648, x25749, x49634);
  nand n49649(x49649, x49648, x49647);
  nand n49650(x49650, x71982, x49637);
  nand n49651(x49651, x25749, x49639);
  nand n49652(x49652, x49651, x49650);
  nand n49653(x49653, x71982, x85581);
  nand n49654(x49654, x25749, x85582);
  nand n49655(x49655, x49654, x49653);
  nand n49656(x49656, x71982, x49634);
  nand n49657(x49657, x25749, x49637);
  nand n49658(x49658, x49657, x49656);
  nand n49659(x49659, x71982, x49641);
  nand n49660(x49660, x25749, x85583);
  nand n49661(x49661, x49660, x49659);
  nand n49662(x49662, x71987, x85584);
  nand n49663(x49663, x25772, x49646);
  nand n49664(x49664, x49663, x27728);
  nand n49665(x49665, x71987, x49649);
  nand n49666(x49666, x25772, x49652);
  nand n49667(x49667, x49666, x49665);
  nand n49668(x49668, x71987, x49655);
  nand n49669(x49669, x25772, x49658);
  nand n49670(x49670, x49669, x49668);
  nand n49671(x49671, x71987, x49661);
  nand n49672(x49672, x25782, x85585);
  nand n49673(x49673, x71992, x49664);
  nand n49674(x49674, x25782, x49667);
  nand n49675(x49675, x49674, x49673);
  nand n49676(x49676, x71992, x49670);
  nand n49677(x49677, x25782, x85586);
  nand n49678(x49678, x49677, x49676);
  nand n49679(x49679, x25790, x85587);
  nand n49680(x49680, x71997, x49675);
  nand n49681(x49681, x25790, x49678);
  nand n49682(x49682, x49681, x49680);
  nand n49683(x49683, x72002, x85588);
  nand n49684(x49684, x25796, x49682);
  nand n49685(x49685, x49684, x49683);
  nand n49686(x49686, x16745, x47856);
  nand n49687(x49687, x68738, x49689);
  nand n49688(x49688, x49687, x49686);
  nand n49690(x49690, x16745, x47915);
  nand n49691(x49691, x68738, x49693);
  nand n49692(x49692, x49691, x49690);
  nand n49694(x49694, x16745, x47974);
  nand n49695(x49695, x68738, x49697);
  nand n49696(x49696, x49695, x49694);
  nand n49698(x49698, x16745, x48033);
  nand n49699(x49699, x68738, x49701);
  nand n49700(x49700, x49699, x49698);
  nand n49702(x49702, x16745, x48092);
  nand n49703(x49703, x68738, x49705);
  nand n49704(x49704, x49703, x49702);
  nand n49706(x49706, x16745, x48151);
  nand n49707(x49707, x68738, x49709);
  nand n49708(x49708, x49707, x49706);
  nand n49710(x49710, x16745, x48210);
  nand n49711(x49711, x68738, x49713);
  nand n49712(x49712, x49711, x49710);
  nand n49714(x49714, x16745, x48269);
  nand n49715(x49715, x68738, x49717);
  nand n49716(x49716, x49715, x49714);
  nand n49718(x49718, x16745, x48328);
  nand n49719(x49719, x68738, x49721);
  nand n49720(x49720, x49719, x49718);
  nand n49722(x49722, x16745, x48387);
  nand n49723(x49723, x68738, x49725);
  nand n49724(x49724, x49723, x49722);
  nand n49726(x49726, x16745, x48446);
  nand n49727(x49727, x68738, x49729);
  nand n49728(x49728, x49727, x49726);
  nand n49730(x49730, x16745, x48505);
  nand n49731(x49731, x68738, x49733);
  nand n49732(x49732, x49731, x49730);
  nand n49734(x49734, x16745, x48564);
  nand n49735(x49735, x68738, x49737);
  nand n49736(x49736, x49735, x49734);
  nand n49738(x49738, x16745, x48623);
  nand n49739(x49739, x68738, x49741);
  nand n49740(x49740, x49739, x49738);
  nand n49742(x49742, x16745, x48682);
  nand n49743(x49743, x68738, x49745);
  nand n49744(x49744, x49743, x49742);
  nand n49746(x49746, x16745, x48741);
  nand n49747(x49747, x68738, x49749);
  nand n49748(x49748, x49747, x49746);
  nand n49750(x49750, x16745, x48800);
  nand n49751(x49751, x68738, x49753);
  nand n49752(x49752, x49751, x49750);
  nand n49754(x49754, x16745, x48859);
  nand n49755(x49755, x68738, x49757);
  nand n49756(x49756, x49755, x49754);
  nand n49758(x49758, x16745, x48918);
  nand n49759(x49759, x68738, x49761);
  nand n49760(x49760, x49759, x49758);
  nand n49762(x49762, x16745, x48977);
  nand n49763(x49763, x68738, x49765);
  nand n49764(x49764, x49763, x49762);
  nand n49766(x49766, x16745, x49036);
  nand n49767(x49767, x68738, x49769);
  nand n49768(x49768, x49767, x49766);
  nand n49770(x49770, x16745, x49095);
  nand n49771(x49771, x68738, x49773);
  nand n49772(x49772, x49771, x49770);
  nand n49774(x49774, x16745, x49154);
  nand n49775(x49775, x68738, x49777);
  nand n49776(x49776, x49775, x49774);
  nand n49778(x49778, x16745, x49213);
  nand n49779(x49779, x68738, x49781);
  nand n49780(x49780, x49779, x49778);
  nand n49782(x49782, x16745, x49272);
  nand n49783(x49783, x68738, x49785);
  nand n49784(x49784, x49783, x49782);
  nand n49786(x49786, x16745, x49331);
  nand n49787(x49787, x68738, x49789);
  nand n49788(x49788, x49787, x49786);
  nand n49790(x49790, x16745, x49390);
  nand n49791(x49791, x68738, x49793);
  nand n49792(x49792, x49791, x49790);
  nand n49794(x49794, x16745, x49449);
  nand n49795(x49795, x68738, x49797);
  nand n49796(x49796, x49795, x49794);
  nand n49798(x49798, x16745, x49508);
  nand n49799(x49799, x68738, x49801);
  nand n49800(x49800, x49799, x49798);
  nand n49802(x49802, x16745, x49567);
  nand n49803(x49803, x68738, x49805);
  nand n49804(x49804, x49803, x49802);
  nand n49806(x49806, x16745, x49626);
  nand n49807(x49807, x68738, x49809);
  nand n49808(x49808, x49807, x49806);
  nand n49810(x49810, x16745, x49685);
  nand n49811(x49811, x68738, x49813);
  nand n49812(x49812, x49811, x49810);
  nand n49814(x49814, x16747, x73677);
  nand n49815(x49815, x49814, x16746);
  nand n49816(x49816, x16747, x73682);
  nand n49817(x49817, x49816, x16750);
  nand n49818(x49818, x16747, x73687);
  nand n49819(x49819, x49818, x16753);
  nand n49820(x49820, x16747, x73692);
  nand n49821(x49821, x49820, x16756);
  nand n49822(x49822, x16747, x73697);
  nand n49823(x49823, x49822, x16759);
  nand n49824(x49824, x16747, x73702);
  nand n49825(x49825, x49824, x16762);
  nand n49826(x49826, x16747, x73707);
  nand n49827(x49827, x49826, x16765);
  nand n49828(x49828, x16747, x73712);
  nand n49829(x49829, x49828, x16768);
  nand n49830(x49830, x16747, x73717);
  nand n49831(x49831, x49830, x16771);
  nand n49832(x49832, x16747, x73722);
  nand n49833(x49833, x49832, x16774);
  nand n49834(x49834, x16747, x73727);
  nand n49835(x49835, x49834, x16777);
  nand n49836(x49836, x16747, x73732);
  nand n49837(x49837, x49836, x16780);
  nand n49838(x49838, x16747, x73737);
  nand n49839(x49839, x49838, x16783);
  nand n49840(x49840, x16747, x73742);
  nand n49841(x49841, x49840, x16786);
  nand n49842(x49842, x16747, x73747);
  nand n49843(x49843, x49842, x16789);
  nand n49844(x49844, x16747, x73752);
  nand n49845(x49845, x49844, x16792);
  nand n49846(x49846, x16747, x73757);
  nand n49847(x49847, x49846, x16795);
  nand n49848(x49848, x16747, x73762);
  nand n49849(x49849, x49848, x16798);
  nand n49850(x49850, x16747, x73767);
  nand n49851(x49851, x49850, x16801);
  nand n49852(x49852, x16747, x73772);
  nand n49853(x49853, x49852, x16804);
  nand n49854(x49854, x16747, x73777);
  nand n49855(x49855, x49854, x16807);
  nand n49856(x49856, x16747, x73782);
  nand n49857(x49857, x49856, x16810);
  nand n49858(x49858, x16747, x73787);
  nand n49859(x49859, x49858, x16813);
  nand n49860(x49860, x16747, x73792);
  nand n49861(x49861, x49860, x16816);
  nand n49862(x49862, x16747, x73797);
  nand n49863(x49863, x49862, x16819);
  nand n49864(x49864, x16747, x73802);
  nand n49865(x49865, x49864, x16822);
  nand n49866(x49866, x16747, x73807);
  nand n49867(x49867, x49866, x16825);
  nand n49868(x49868, x16747, x73812);
  nand n49869(x49869, x49868, x16828);
  nand n49870(x49870, x16747, x73817);
  nand n49871(x49871, x49870, x16831);
  nand n49872(x49872, x16747, x73822);
  nand n49873(x49873, x49872, x16834);
  nand n49874(x49874, x16747, x73827);
  nand n49875(x49875, x49874, x16837);
  nand n49876(x49876, x16747, x73832);
  nand n49877(x49877, x49876, x16840);
  nand n49910(x49910, x71977, x49878);
  nand n49911(x49911, x16876, x49815);
  nand n49912(x49912, x49911, x49910);
  nand n49913(x49913, x71977, x49879);
  nand n49914(x49914, x16876, x49817);
  nand n49915(x49915, x49914, x49913);
  nand n49916(x49916, x71977, x49880);
  nand n49917(x49917, x16876, x49819);
  nand n49918(x49918, x49917, x49916);
  nand n49919(x49919, x71977, x49881);
  nand n49920(x49920, x16876, x49821);
  nand n49921(x49921, x49920, x49919);
  nand n49922(x49922, x71977, x49882);
  nand n49923(x49923, x16876, x49823);
  nand n49924(x49924, x49923, x49922);
  nand n49925(x49925, x71977, x49883);
  nand n49926(x49926, x16876, x49825);
  nand n49927(x49927, x49926, x49925);
  nand n49928(x49928, x71977, x49884);
  nand n49929(x49929, x16876, x49827);
  nand n49930(x49930, x49929, x49928);
  nand n49931(x49931, x71977, x49885);
  nand n49932(x49932, x16876, x49829);
  nand n49933(x49933, x49932, x49931);
  nand n49934(x49934, x71977, x49886);
  nand n49935(x49935, x16876, x49831);
  nand n49936(x49936, x49935, x49934);
  nand n49937(x49937, x71977, x49887);
  nand n49938(x49938, x16876, x49833);
  nand n49939(x49939, x49938, x49937);
  nand n49940(x49940, x71977, x49888);
  nand n49941(x49941, x16876, x49835);
  nand n49942(x49942, x49941, x49940);
  nand n49943(x49943, x71977, x49889);
  nand n49944(x49944, x16876, x49837);
  nand n49945(x49945, x49944, x49943);
  nand n49946(x49946, x71977, x49890);
  nand n49947(x49947, x16876, x49839);
  nand n49948(x49948, x49947, x49946);
  nand n49949(x49949, x71977, x49891);
  nand n49950(x49950, x16876, x49841);
  nand n49951(x49951, x49950, x49949);
  nand n49952(x49952, x71977, x49892);
  nand n49953(x49953, x16876, x49843);
  nand n49954(x49954, x49953, x49952);
  nand n49955(x49955, x71977, x49893);
  nand n49956(x49956, x16876, x49845);
  nand n49957(x49957, x49956, x49955);
  nand n49958(x49958, x71977, x49894);
  nand n49959(x49959, x16876, x49847);
  nand n49960(x49960, x49959, x49958);
  nand n49961(x49961, x71977, x49895);
  nand n49962(x49962, x16876, x49849);
  nand n49963(x49963, x49962, x49961);
  nand n49964(x49964, x71977, x49896);
  nand n49965(x49965, x16876, x49851);
  nand n49966(x49966, x49965, x49964);
  nand n49967(x49967, x71977, x49897);
  nand n49968(x49968, x16876, x49853);
  nand n49969(x49969, x49968, x49967);
  nand n49970(x49970, x71977, x49898);
  nand n49971(x49971, x16876, x49855);
  nand n49972(x49972, x49971, x49970);
  nand n49973(x49973, x71977, x49899);
  nand n49974(x49974, x16876, x49857);
  nand n49975(x49975, x49974, x49973);
  nand n49976(x49976, x71977, x49900);
  nand n49977(x49977, x16876, x49859);
  nand n49978(x49978, x49977, x49976);
  nand n49979(x49979, x71977, x49901);
  nand n49980(x49980, x16876, x49861);
  nand n49981(x49981, x49980, x49979);
  nand n49982(x49982, x71977, x49902);
  nand n49983(x49983, x16876, x49863);
  nand n49984(x49984, x49983, x49982);
  nand n49985(x49985, x71977, x49903);
  nand n49986(x49986, x16876, x49865);
  nand n49987(x49987, x49986, x49985);
  nand n49988(x49988, x71977, x49904);
  nand n49989(x49989, x16876, x49867);
  nand n49990(x49990, x49989, x49988);
  nand n49991(x49991, x71977, x49905);
  nand n49992(x49992, x16876, x49869);
  nand n49993(x49993, x49992, x49991);
  nand n49994(x49994, x71977, x49906);
  nand n49995(x49995, x16876, x49871);
  nand n49996(x49996, x49995, x49994);
  nand n49997(x49997, x71977, x49907);
  nand n49998(x49998, x16876, x49873);
  nand n49999(x49999, x49998, x49997);
  nand n50000(x50000, x71977, x49908);
  nand n50001(x50001, x16876, x49875);
  nand n50002(x50002, x50001, x50000);
  nand n50003(x50003, x71977, x49909);
  nand n50004(x50004, x16876, x49877);
  nand n50005(x50005, x50004, x50003);
  nand n50006(x50006, x73517, x49912);
  nand n50009(x50009, x50008, x50007);
  nand n50010(x50010, x50009, x50006);
  nand n50012(x50012, x73522, x49915);
  nand n50015(x50015, x50014, x50013);
  nand n50016(x50016, x50015, x50012);
  nand n50018(x50018, x73527, x49918);
  nand n50021(x50021, x50020, x50019);
  nand n50022(x50022, x50021, x50018);
  nand n50024(x50024, x73532, x49921);
  nand n50027(x50027, x50026, x50025);
  nand n50028(x50028, x50027, x50024);
  nand n50030(x50030, x73537, x49924);
  nand n50033(x50033, x50032, x50031);
  nand n50034(x50034, x50033, x50030);
  nand n50036(x50036, x73542, x49927);
  nand n50039(x50039, x50038, x50037);
  nand n50040(x50040, x50039, x50036);
  nand n50042(x50042, x73547, x49930);
  nand n50045(x50045, x50044, x50043);
  nand n50046(x50046, x50045, x50042);
  nand n50048(x50048, x73552, x49933);
  nand n50051(x50051, x50050, x50049);
  nand n50052(x50052, x50051, x50048);
  nand n50054(x50054, x73557, x49936);
  nand n50057(x50057, x50056, x50055);
  nand n50058(x50058, x50057, x50054);
  nand n50060(x50060, x73562, x49939);
  nand n50063(x50063, x50062, x50061);
  nand n50064(x50064, x50063, x50060);
  nand n50066(x50066, x73567, x49942);
  nand n50069(x50069, x50068, x50067);
  nand n50070(x50070, x50069, x50066);
  nand n50072(x50072, x73572, x49945);
  nand n50075(x50075, x50074, x50073);
  nand n50076(x50076, x50075, x50072);
  nand n50078(x50078, x73577, x49948);
  nand n50081(x50081, x50080, x50079);
  nand n50082(x50082, x50081, x50078);
  nand n50084(x50084, x73582, x49951);
  nand n50087(x50087, x50086, x50085);
  nand n50088(x50088, x50087, x50084);
  nand n50090(x50090, x73587, x49954);
  nand n50093(x50093, x50092, x50091);
  nand n50094(x50094, x50093, x50090);
  nand n50096(x50096, x73592, x49957);
  nand n50099(x50099, x50098, x50097);
  nand n50100(x50100, x50099, x50096);
  nand n50102(x50102, x73597, x49960);
  nand n50105(x50105, x50104, x50103);
  nand n50106(x50106, x50105, x50102);
  nand n50108(x50108, x73602, x49963);
  nand n50111(x50111, x50110, x50109);
  nand n50112(x50112, x50111, x50108);
  nand n50114(x50114, x73607, x49966);
  nand n50117(x50117, x50116, x50115);
  nand n50118(x50118, x50117, x50114);
  nand n50120(x50120, x73612, x49969);
  nand n50123(x50123, x50122, x50121);
  nand n50124(x50124, x50123, x50120);
  nand n50126(x50126, x73617, x49972);
  nand n50129(x50129, x50128, x50127);
  nand n50130(x50130, x50129, x50126);
  nand n50132(x50132, x73622, x49975);
  nand n50135(x50135, x50134, x50133);
  nand n50136(x50136, x50135, x50132);
  nand n50138(x50138, x73627, x49978);
  nand n50141(x50141, x50140, x50139);
  nand n50142(x50142, x50141, x50138);
  nand n50144(x50144, x73632, x49981);
  nand n50147(x50147, x50146, x50145);
  nand n50148(x50148, x50147, x50144);
  nand n50150(x50150, x73637, x49984);
  nand n50153(x50153, x50152, x50151);
  nand n50154(x50154, x50153, x50150);
  nand n50156(x50156, x73642, x49987);
  nand n50159(x50159, x50158, x50157);
  nand n50160(x50160, x50159, x50156);
  nand n50162(x50162, x73647, x49990);
  nand n50165(x50165, x50164, x50163);
  nand n50166(x50166, x50165, x50162);
  nand n50168(x50168, x73652, x49993);
  nand n50171(x50171, x50170, x50169);
  nand n50172(x50172, x50171, x50168);
  nand n50174(x50174, x73657, x49996);
  nand n50177(x50177, x50176, x50175);
  nand n50178(x50178, x50177, x50174);
  nand n50180(x50180, x73662, x49999);
  nand n50183(x50183, x50182, x50181);
  nand n50184(x50184, x50183, x50180);
  nand n50186(x50186, x73667, x50002);
  nand n50189(x50189, x50188, x50187);
  nand n50190(x50190, x50189, x50186);
  nand n50192(x50192, x73672, x50005);
  nand n50195(x50195, x50194, x50193);
  nand n50196(x50196, x50195, x50192);
  nand n50228(x50228, x50011, x71977);
  nand n50229(x50229, x50228, x50006);
  nand n50230(x50230, x50017, x50198);
  nand n50231(x50231, x50230, x50012);
  nand n50232(x50232, x50017, x50011);
  nand n50234(x50234, x50023, x50199);
  nand n50235(x50235, x50234, x50018);
  nand n50236(x50236, x50023, x50017);
  nand n50238(x50238, x50029, x50200);
  nand n50239(x50239, x50238, x50024);
  nand n50240(x50240, x50029, x50023);
  nand n50242(x50242, x50035, x50201);
  nand n50243(x50243, x50242, x50030);
  nand n50244(x50244, x50035, x50029);
  nand n50246(x50246, x50041, x50202);
  nand n50247(x50247, x50246, x50036);
  nand n50248(x50248, x50041, x50035);
  nand n50250(x50250, x50047, x50203);
  nand n50251(x50251, x50250, x50042);
  nand n50252(x50252, x50047, x50041);
  nand n50254(x50254, x50053, x50204);
  nand n50255(x50255, x50254, x50048);
  nand n50256(x50256, x50053, x50047);
  nand n50258(x50258, x50059, x50205);
  nand n50259(x50259, x50258, x50054);
  nand n50260(x50260, x50059, x50053);
  nand n50262(x50262, x50065, x50206);
  nand n50263(x50263, x50262, x50060);
  nand n50264(x50264, x50065, x50059);
  nand n50266(x50266, x50071, x50207);
  nand n50267(x50267, x50266, x50066);
  nand n50268(x50268, x50071, x50065);
  nand n50270(x50270, x50077, x50208);
  nand n50271(x50271, x50270, x50072);
  nand n50272(x50272, x50077, x50071);
  nand n50274(x50274, x50083, x50209);
  nand n50275(x50275, x50274, x50078);
  nand n50276(x50276, x50083, x50077);
  nand n50278(x50278, x50089, x50210);
  nand n50279(x50279, x50278, x50084);
  nand n50280(x50280, x50089, x50083);
  nand n50282(x50282, x50095, x50211);
  nand n50283(x50283, x50282, x50090);
  nand n50284(x50284, x50095, x50089);
  nand n50286(x50286, x50101, x50212);
  nand n50287(x50287, x50286, x50096);
  nand n50288(x50288, x50101, x50095);
  nand n50290(x50290, x50107, x50213);
  nand n50291(x50291, x50290, x50102);
  nand n50292(x50292, x50107, x50101);
  nand n50294(x50294, x50113, x50214);
  nand n50295(x50295, x50294, x50108);
  nand n50296(x50296, x50113, x50107);
  nand n50298(x50298, x50119, x50215);
  nand n50299(x50299, x50298, x50114);
  nand n50300(x50300, x50119, x50113);
  nand n50302(x50302, x50125, x50216);
  nand n50303(x50303, x50302, x50120);
  nand n50304(x50304, x50125, x50119);
  nand n50306(x50306, x50131, x50217);
  nand n50307(x50307, x50306, x50126);
  nand n50308(x50308, x50131, x50125);
  nand n50310(x50310, x50137, x50218);
  nand n50311(x50311, x50310, x50132);
  nand n50312(x50312, x50137, x50131);
  nand n50314(x50314, x50143, x50219);
  nand n50315(x50315, x50314, x50138);
  nand n50316(x50316, x50143, x50137);
  nand n50318(x50318, x50149, x50220);
  nand n50319(x50319, x50318, x50144);
  nand n50320(x50320, x50149, x50143);
  nand n50322(x50322, x50155, x50221);
  nand n50323(x50323, x50322, x50150);
  nand n50324(x50324, x50155, x50149);
  nand n50326(x50326, x50161, x50222);
  nand n50327(x50327, x50326, x50156);
  nand n50328(x50328, x50161, x50155);
  nand n50330(x50330, x50167, x50223);
  nand n50331(x50331, x50330, x50162);
  nand n50332(x50332, x50167, x50161);
  nand n50334(x50334, x50173, x50224);
  nand n50335(x50335, x50334, x50168);
  nand n50336(x50336, x50173, x50167);
  nand n50338(x50338, x50179, x50225);
  nand n50339(x50339, x50338, x50174);
  nand n50340(x50340, x50179, x50173);
  nand n50342(x50342, x50185, x50226);
  nand n50343(x50343, x50342, x50180);
  nand n50344(x50344, x50185, x50179);
  nand n50346(x50346, x50191, x50227);
  nand n50347(x50347, x50346, x50186);
  nand n50348(x50348, x50191, x50185);
  nand n50350(x50350, x50233, x71977);
  nand n50352(x50352, x50350, x50351);
  nand n50353(x50353, x50237, x50229);
  nand n50355(x50355, x50353, x50354);
  nand n50356(x50356, x50241, x50231);
  nand n50358(x50358, x50356, x50357);
  nand n50359(x50359, x50241, x50233);
  nand n50361(x50361, x50245, x50235);
  nand n50363(x50363, x50361, x50362);
  nand n50364(x50364, x50245, x50237);
  nand n50366(x50366, x50249, x50239);
  nand n50368(x50368, x50366, x50367);
  nand n50369(x50369, x50249, x50241);
  nand n50371(x50371, x50253, x50243);
  nand n50373(x50373, x50371, x50372);
  nand n50374(x50374, x50253, x50245);
  nand n50376(x50376, x50257, x50247);
  nand n50378(x50378, x50376, x50377);
  nand n50379(x50379, x50257, x50249);
  nand n50381(x50381, x50261, x50251);
  nand n50383(x50383, x50381, x50382);
  nand n50384(x50384, x50261, x50253);
  nand n50386(x50386, x50265, x50255);
  nand n50388(x50388, x50386, x50387);
  nand n50389(x50389, x50265, x50257);
  nand n50391(x50391, x50269, x50259);
  nand n50393(x50393, x50391, x50392);
  nand n50394(x50394, x50269, x50261);
  nand n50396(x50396, x50273, x50263);
  nand n50398(x50398, x50396, x50397);
  nand n50399(x50399, x50273, x50265);
  nand n50401(x50401, x50277, x50267);
  nand n50403(x50403, x50401, x50402);
  nand n50404(x50404, x50277, x50269);
  nand n50406(x50406, x50281, x50271);
  nand n50408(x50408, x50406, x50407);
  nand n50409(x50409, x50281, x50273);
  nand n50411(x50411, x50285, x50275);
  nand n50413(x50413, x50411, x50412);
  nand n50414(x50414, x50285, x50277);
  nand n50416(x50416, x50289, x50279);
  nand n50418(x50418, x50416, x50417);
  nand n50419(x50419, x50289, x50281);
  nand n50421(x50421, x50293, x50283);
  nand n50423(x50423, x50421, x50422);
  nand n50424(x50424, x50293, x50285);
  nand n50426(x50426, x50297, x50287);
  nand n50428(x50428, x50426, x50427);
  nand n50429(x50429, x50297, x50289);
  nand n50431(x50431, x50301, x50291);
  nand n50433(x50433, x50431, x50432);
  nand n50434(x50434, x50301, x50293);
  nand n50436(x50436, x50305, x50295);
  nand n50438(x50438, x50436, x50437);
  nand n50439(x50439, x50305, x50297);
  nand n50441(x50441, x50309, x50299);
  nand n50443(x50443, x50441, x50442);
  nand n50444(x50444, x50309, x50301);
  nand n50446(x50446, x50313, x50303);
  nand n50448(x50448, x50446, x50447);
  nand n50449(x50449, x50313, x50305);
  nand n50451(x50451, x50317, x50307);
  nand n50453(x50453, x50451, x50452);
  nand n50454(x50454, x50317, x50309);
  nand n50456(x50456, x50321, x50311);
  nand n50458(x50458, x50456, x50457);
  nand n50459(x50459, x50321, x50313);
  nand n50461(x50461, x50325, x50315);
  nand n50463(x50463, x50461, x50462);
  nand n50464(x50464, x50325, x50317);
  nand n50466(x50466, x50329, x50319);
  nand n50468(x50468, x50466, x50467);
  nand n50469(x50469, x50329, x50321);
  nand n50471(x50471, x50333, x50323);
  nand n50473(x50473, x50471, x50472);
  nand n50474(x50474, x50333, x50325);
  nand n50476(x50476, x50337, x50327);
  nand n50478(x50478, x50476, x50477);
  nand n50479(x50479, x50337, x50329);
  nand n50481(x50481, x50341, x50331);
  nand n50483(x50483, x50481, x50482);
  nand n50484(x50484, x50341, x50333);
  nand n50486(x50486, x50345, x50335);
  nand n50488(x50488, x50486, x50487);
  nand n50489(x50489, x50345, x50337);
  nand n50491(x50491, x50349, x50339);
  nand n50493(x50493, x50491, x50492);
  nand n50494(x50494, x50349, x50341);
  nand n50496(x50496, x50360, x71977);
  nand n50498(x50498, x50496, x50497);
  nand n50499(x50499, x50365, x50229);
  nand n50501(x50501, x50499, x50500);
  nand n50502(x50502, x50370, x50352);
  nand n50504(x50504, x50502, x50503);
  nand n50505(x50505, x50375, x50355);
  nand n50507(x50507, x50505, x50506);
  nand n50508(x50508, x50380, x50358);
  nand n50510(x50510, x50508, x50509);
  nand n50511(x50511, x50380, x50360);
  nand n50513(x50513, x50385, x50363);
  nand n50515(x50515, x50513, x50514);
  nand n50516(x50516, x50385, x50365);
  nand n50518(x50518, x50390, x50368);
  nand n50520(x50520, x50518, x50519);
  nand n50521(x50521, x50390, x50370);
  nand n50523(x50523, x50395, x50373);
  nand n50525(x50525, x50523, x50524);
  nand n50526(x50526, x50395, x50375);
  nand n50528(x50528, x50400, x50378);
  nand n50530(x50530, x50528, x50529);
  nand n50531(x50531, x50400, x50380);
  nand n50533(x50533, x50405, x50383);
  nand n50535(x50535, x50533, x50534);
  nand n50536(x50536, x50405, x50385);
  nand n50538(x50538, x50410, x50388);
  nand n50540(x50540, x50538, x50539);
  nand n50541(x50541, x50410, x50390);
  nand n50543(x50543, x50415, x50393);
  nand n50545(x50545, x50543, x50544);
  nand n50546(x50546, x50415, x50395);
  nand n50548(x50548, x50420, x50398);
  nand n50550(x50550, x50548, x50549);
  nand n50551(x50551, x50420, x50400);
  nand n50553(x50553, x50425, x50403);
  nand n50555(x50555, x50553, x50554);
  nand n50556(x50556, x50425, x50405);
  nand n50558(x50558, x50430, x50408);
  nand n50560(x50560, x50558, x50559);
  nand n50561(x50561, x50430, x50410);
  nand n50563(x50563, x50435, x50413);
  nand n50565(x50565, x50563, x50564);
  nand n50566(x50566, x50435, x50415);
  nand n50568(x50568, x50440, x50418);
  nand n50570(x50570, x50568, x50569);
  nand n50571(x50571, x50440, x50420);
  nand n50573(x50573, x50445, x50423);
  nand n50575(x50575, x50573, x50574);
  nand n50576(x50576, x50445, x50425);
  nand n50578(x50578, x50450, x50428);
  nand n50580(x50580, x50578, x50579);
  nand n50581(x50581, x50450, x50430);
  nand n50583(x50583, x50455, x50433);
  nand n50585(x50585, x50583, x50584);
  nand n50586(x50586, x50455, x50435);
  nand n50588(x50588, x50460, x50438);
  nand n50590(x50590, x50588, x50589);
  nand n50591(x50591, x50460, x50440);
  nand n50593(x50593, x50465, x50443);
  nand n50595(x50595, x50593, x50594);
  nand n50596(x50596, x50465, x50445);
  nand n50598(x50598, x50470, x50448);
  nand n50600(x50600, x50598, x50599);
  nand n50601(x50601, x50470, x50450);
  nand n50603(x50603, x50475, x50453);
  nand n50605(x50605, x50603, x50604);
  nand n50606(x50606, x50475, x50455);
  nand n50608(x50608, x50480, x50458);
  nand n50610(x50610, x50608, x50609);
  nand n50611(x50611, x50480, x50460);
  nand n50613(x50613, x50485, x50463);
  nand n50615(x50615, x50613, x50614);
  nand n50616(x50616, x50485, x50465);
  nand n50618(x50618, x50490, x50468);
  nand n50620(x50620, x50618, x50619);
  nand n50621(x50621, x50490, x50470);
  nand n50623(x50623, x50495, x50473);
  nand n50625(x50625, x50623, x50624);
  nand n50626(x50626, x50495, x50475);
  nand n50628(x50628, x50512, x71977);
  nand n50630(x50630, x50628, x50629);
  nand n50631(x50631, x50517, x50229);
  nand n50633(x50633, x50631, x50632);
  nand n50634(x50634, x50522, x50352);
  nand n50636(x50636, x50634, x50635);
  nand n50637(x50637, x50527, x50355);
  nand n50639(x50639, x50637, x50638);
  nand n50640(x50640, x50532, x50498);
  nand n50642(x50642, x50640, x50641);
  nand n50643(x50643, x50537, x50501);
  nand n50645(x50645, x50643, x50644);
  nand n50646(x50646, x50542, x50504);
  nand n50648(x50648, x50646, x50647);
  nand n50649(x50649, x50547, x50507);
  nand n50651(x50651, x50649, x50650);
  nand n50652(x50652, x50552, x50510);
  nand n50654(x50654, x50652, x50653);
  nand n50655(x50655, x50552, x50512);
  nand n50657(x50657, x50557, x50515);
  nand n50659(x50659, x50657, x50658);
  nand n50660(x50660, x50557, x50517);
  nand n50662(x50662, x50562, x50520);
  nand n50664(x50664, x50662, x50663);
  nand n50665(x50665, x50562, x50522);
  nand n50667(x50667, x50567, x50525);
  nand n50669(x50669, x50667, x50668);
  nand n50670(x50670, x50567, x50527);
  nand n50672(x50672, x50572, x50530);
  nand n50674(x50674, x50672, x50673);
  nand n50675(x50675, x50572, x50532);
  nand n50677(x50677, x50577, x50535);
  nand n50679(x50679, x50677, x50678);
  nand n50680(x50680, x50577, x50537);
  nand n50682(x50682, x50582, x50540);
  nand n50684(x50684, x50682, x50683);
  nand n50685(x50685, x50582, x50542);
  nand n50687(x50687, x50587, x50545);
  nand n50689(x50689, x50687, x50688);
  nand n50690(x50690, x50587, x50547);
  nand n50692(x50692, x50592, x50550);
  nand n50694(x50694, x50692, x50693);
  nand n50695(x50695, x50592, x50552);
  nand n50697(x50697, x50597, x50555);
  nand n50699(x50699, x50697, x50698);
  nand n50700(x50700, x50597, x50557);
  nand n50702(x50702, x50602, x50560);
  nand n50704(x50704, x50702, x50703);
  nand n50705(x50705, x50602, x50562);
  nand n50707(x50707, x50607, x50565);
  nand n50709(x50709, x50707, x50708);
  nand n50710(x50710, x50607, x50567);
  nand n50712(x50712, x50612, x50570);
  nand n50714(x50714, x50712, x50713);
  nand n50715(x50715, x50612, x50572);
  nand n50717(x50717, x50617, x50575);
  nand n50719(x50719, x50717, x50718);
  nand n50720(x50720, x50617, x50577);
  nand n50722(x50722, x50622, x50580);
  nand n50724(x50724, x50722, x50723);
  nand n50725(x50725, x50622, x50582);
  nand n50727(x50727, x50627, x50585);
  nand n50729(x50729, x50727, x50728);
  nand n50730(x50730, x50627, x50587);
  nand n50732(x50732, x50656, x71977);
  nand n50734(x50734, x50732, x50733);
  nand n50735(x50735, x50661, x50229);
  nand n50737(x50737, x50735, x50736);
  nand n50738(x50738, x50666, x50352);
  nand n50740(x50740, x50738, x50739);
  nand n50741(x50741, x50671, x50355);
  nand n50743(x50743, x50741, x50742);
  nand n50744(x50744, x50676, x50498);
  nand n50746(x50746, x50744, x50745);
  nand n50747(x50747, x50681, x50501);
  nand n50749(x50749, x50747, x50748);
  nand n50750(x50750, x50686, x50504);
  nand n50752(x50752, x50750, x50751);
  nand n50753(x50753, x50691, x50507);
  nand n50755(x50755, x50753, x50754);
  nand n50756(x50756, x50696, x50630);
  nand n50758(x50758, x50756, x50757);
  nand n50759(x50759, x50701, x50633);
  nand n50761(x50761, x50759, x50760);
  nand n50762(x50762, x50706, x50636);
  nand n50764(x50764, x50762, x50763);
  nand n50765(x50765, x50711, x50639);
  nand n50767(x50767, x50765, x50766);
  nand n50768(x50768, x50716, x50642);
  nand n50770(x50770, x50768, x50769);
  nand n50771(x50771, x50721, x50645);
  nand n50773(x50773, x50771, x50772);
  nand n50774(x50774, x50726, x50648);
  nand n50776(x50776, x50774, x50775);
  nand n50777(x50777, x50731, x50651);
  nand n50779(x50779, x50777, x50778);
  nand n50780(x50780, x50010, x16876);
  nand n50781(x50781, x50780, x50228);
  nand n50783(x50783, x50017, x50229);
  nand n50785(x50785, x50016, x50784);
  nand n50786(x50786, x50785, x50783);
  nand n50788(x50788, x50023, x50352);
  nand n50790(x50790, x50022, x50789);
  nand n50791(x50791, x50790, x50788);
  nand n50793(x50793, x50029, x50355);
  nand n50795(x50795, x50028, x50794);
  nand n50796(x50796, x50795, x50793);
  nand n50798(x50798, x50035, x50498);
  nand n50800(x50800, x50034, x50799);
  nand n50801(x50801, x50800, x50798);
  nand n50803(x50803, x50041, x50501);
  nand n50805(x50805, x50040, x50804);
  nand n50806(x50806, x50805, x50803);
  nand n50808(x50808, x50047, x50504);
  nand n50810(x50810, x50046, x50809);
  nand n50811(x50811, x50810, x50808);
  nand n50813(x50813, x50053, x50507);
  nand n50815(x50815, x50052, x50814);
  nand n50816(x50816, x50815, x50813);
  nand n50818(x50818, x50059, x50630);
  nand n50820(x50820, x50058, x50819);
  nand n50821(x50821, x50820, x50818);
  nand n50823(x50823, x50065, x50633);
  nand n50825(x50825, x50064, x50824);
  nand n50826(x50826, x50825, x50823);
  nand n50828(x50828, x50071, x50636);
  nand n50830(x50830, x50070, x50829);
  nand n50831(x50831, x50830, x50828);
  nand n50833(x50833, x50077, x50639);
  nand n50835(x50835, x50076, x50834);
  nand n50836(x50836, x50835, x50833);
  nand n50838(x50838, x50083, x50642);
  nand n50840(x50840, x50082, x50839);
  nand n50841(x50841, x50840, x50838);
  nand n50843(x50843, x50089, x50645);
  nand n50845(x50845, x50088, x50844);
  nand n50846(x50846, x50845, x50843);
  nand n50848(x50848, x50095, x50648);
  nand n50850(x50850, x50094, x50849);
  nand n50851(x50851, x50850, x50848);
  nand n50853(x50853, x50101, x50651);
  nand n50855(x50855, x50100, x50854);
  nand n50856(x50856, x50855, x50853);
  nand n50858(x50858, x50107, x50734);
  nand n50860(x50860, x50106, x50859);
  nand n50861(x50861, x50860, x50858);
  nand n50863(x50863, x50113, x50737);
  nand n50865(x50865, x50112, x50864);
  nand n50866(x50866, x50865, x50863);
  nand n50868(x50868, x50119, x50740);
  nand n50870(x50870, x50118, x50869);
  nand n50871(x50871, x50870, x50868);
  nand n50873(x50873, x50125, x50743);
  nand n50875(x50875, x50124, x50874);
  nand n50876(x50876, x50875, x50873);
  nand n50878(x50878, x50131, x50746);
  nand n50880(x50880, x50130, x50879);
  nand n50881(x50881, x50880, x50878);
  nand n50883(x50883, x50137, x50749);
  nand n50885(x50885, x50136, x50884);
  nand n50886(x50886, x50885, x50883);
  nand n50888(x50888, x50143, x50752);
  nand n50890(x50890, x50142, x50889);
  nand n50891(x50891, x50890, x50888);
  nand n50893(x50893, x50149, x50755);
  nand n50895(x50895, x50148, x50894);
  nand n50896(x50896, x50895, x50893);
  nand n50898(x50898, x50155, x50758);
  nand n50900(x50900, x50154, x50899);
  nand n50901(x50901, x50900, x50898);
  nand n50903(x50903, x50161, x50761);
  nand n50905(x50905, x50160, x50904);
  nand n50906(x50906, x50905, x50903);
  nand n50908(x50908, x50167, x50764);
  nand n50910(x50910, x50166, x50909);
  nand n50911(x50911, x50910, x50908);
  nand n50913(x50913, x50173, x50767);
  nand n50915(x50915, x50172, x50914);
  nand n50916(x50916, x50915, x50913);
  nand n50918(x50918, x50179, x50770);
  nand n50920(x50920, x50178, x50919);
  nand n50921(x50921, x50920, x50918);
  nand n50923(x50923, x50185, x50773);
  nand n50925(x50925, x50184, x50924);
  nand n50926(x50926, x50925, x50923);
  nand n50928(x50928, x50191, x50776);
  nand n50930(x50930, x50190, x50929);
  nand n50931(x50931, x50930, x50928);
  nand n50933(x50933, x50197, x50779);
  nand n50935(x50935, x50196, x50934);
  nand n50936(x50936, x50935, x50933);
  nand n50938(x50938, x73517, x49815);
  nand n50939(x50939, x73522, x49815);
  nand n50941(x50941, x73517, x49817);
  nand n50943(x50943, x73527, x49815);
  nand n50945(x50945, x73522, x49817);
  nand n50947(x50947, x73517, x49819);
  nand n50949(x50949, x73532, x49815);
  nand n50951(x50951, x73527, x49817);
  nand n50953(x50953, x73522, x49819);
  nand n50955(x50955, x73517, x49821);
  nand n50956(x50956, x73537, x49815);
  nand n50958(x50958, x73532, x49817);
  nand n50960(x50960, x73527, x49819);
  nand n50962(x50962, x73522, x49821);
  nand n50964(x50964, x73517, x49823);
  nand n50966(x50966, x73542, x49815);
  nand n50968(x50968, x73537, x49817);
  nand n50970(x50970, x73532, x49819);
  nand n50972(x50972, x73527, x49821);
  nand n50974(x50974, x73522, x49823);
  nand n50976(x50976, x73517, x49825);
  nand n50978(x50978, x73547, x49815);
  nand n50980(x50980, x73542, x49817);
  nand n50982(x50982, x73537, x49819);
  nand n50984(x50984, x73532, x49821);
  nand n50986(x50986, x73527, x49823);
  nand n50988(x50988, x73522, x49825);
  nand n50990(x50990, x73517, x49827);
  nand n50991(x50991, x73552, x49815);
  nand n50993(x50993, x73547, x49817);
  nand n50995(x50995, x73542, x49819);
  nand n50997(x50997, x73537, x49821);
  nand n50999(x50999, x73532, x49823);
  nand n51001(x51001, x73527, x49825);
  nand n51003(x51003, x73522, x49827);
  nand n51005(x51005, x73517, x49829);
  nand n51007(x51007, x73557, x49815);
  nand n51009(x51009, x73552, x49817);
  nand n51011(x51011, x73547, x49819);
  nand n51013(x51013, x73542, x49821);
  nand n51015(x51015, x73537, x49823);
  nand n51017(x51017, x73532, x49825);
  nand n51019(x51019, x73527, x49827);
  nand n51021(x51021, x73522, x49829);
  nand n51023(x51023, x73517, x49831);
  nand n51025(x51025, x73562, x49815);
  nand n51027(x51027, x73557, x49817);
  nand n51029(x51029, x73552, x49819);
  nand n51031(x51031, x73547, x49821);
  nand n51033(x51033, x73542, x49823);
  nand n51035(x51035, x73537, x49825);
  nand n51037(x51037, x73532, x49827);
  nand n51039(x51039, x73527, x49829);
  nand n51041(x51041, x73522, x49831);
  nand n51043(x51043, x73517, x49833);
  nand n51044(x51044, x73567, x49815);
  nand n51046(x51046, x73562, x49817);
  nand n51048(x51048, x73557, x49819);
  nand n51050(x51050, x73552, x49821);
  nand n51052(x51052, x73547, x49823);
  nand n51054(x51054, x73542, x49825);
  nand n51056(x51056, x73537, x49827);
  nand n51058(x51058, x73532, x49829);
  nand n51060(x51060, x73527, x49831);
  nand n51062(x51062, x73522, x49833);
  nand n51064(x51064, x73517, x49835);
  nand n51066(x51066, x73572, x49815);
  nand n51068(x51068, x73567, x49817);
  nand n51070(x51070, x73562, x49819);
  nand n51072(x51072, x73557, x49821);
  nand n51074(x51074, x73552, x49823);
  nand n51076(x51076, x73547, x49825);
  nand n51078(x51078, x73542, x49827);
  nand n51080(x51080, x73537, x49829);
  nand n51082(x51082, x73532, x49831);
  nand n51084(x51084, x73527, x49833);
  nand n51086(x51086, x73522, x49835);
  nand n51088(x51088, x73517, x49837);
  nand n51090(x51090, x73577, x49815);
  nand n51092(x51092, x73572, x49817);
  nand n51094(x51094, x73567, x49819);
  nand n51096(x51096, x73562, x49821);
  nand n51098(x51098, x73557, x49823);
  nand n51100(x51100, x73552, x49825);
  nand n51102(x51102, x73547, x49827);
  nand n51104(x51104, x73542, x49829);
  nand n51106(x51106, x73537, x49831);
  nand n51108(x51108, x73532, x49833);
  nand n51110(x51110, x73527, x49835);
  nand n51112(x51112, x73522, x49837);
  nand n51114(x51114, x73517, x49839);
  nand n51115(x51115, x73582, x49815);
  nand n51117(x51117, x73577, x49817);
  nand n51119(x51119, x73572, x49819);
  nand n51121(x51121, x73567, x49821);
  nand n51123(x51123, x73562, x49823);
  nand n51125(x51125, x73557, x49825);
  nand n51127(x51127, x73552, x49827);
  nand n51129(x51129, x73547, x49829);
  nand n51131(x51131, x73542, x49831);
  nand n51133(x51133, x73537, x49833);
  nand n51135(x51135, x73532, x49835);
  nand n51137(x51137, x73527, x49837);
  nand n51139(x51139, x73522, x49839);
  nand n51141(x51141, x73517, x49841);
  nand n51143(x51143, x73587, x49815);
  nand n51145(x51145, x73582, x49817);
  nand n51147(x51147, x73577, x49819);
  nand n51149(x51149, x73572, x49821);
  nand n51151(x51151, x73567, x49823);
  nand n51153(x51153, x73562, x49825);
  nand n51155(x51155, x73557, x49827);
  nand n51157(x51157, x73552, x49829);
  nand n51159(x51159, x73547, x49831);
  nand n51161(x51161, x73542, x49833);
  nand n51163(x51163, x73537, x49835);
  nand n51165(x51165, x73532, x49837);
  nand n51167(x51167, x73527, x49839);
  nand n51169(x51169, x73522, x49841);
  nand n51171(x51171, x73517, x49843);
  nand n51173(x51173, x73592, x49815);
  nand n51175(x51175, x73587, x49817);
  nand n51177(x51177, x73582, x49819);
  nand n51179(x51179, x73577, x49821);
  nand n51181(x51181, x73572, x49823);
  nand n51183(x51183, x73567, x49825);
  nand n51185(x51185, x73562, x49827);
  nand n51187(x51187, x73557, x49829);
  nand n51189(x51189, x73552, x49831);
  nand n51191(x51191, x73547, x49833);
  nand n51193(x51193, x73542, x49835);
  nand n51195(x51195, x73537, x49837);
  nand n51197(x51197, x73532, x49839);
  nand n51199(x51199, x73527, x49841);
  nand n51201(x51201, x73522, x49843);
  nand n51203(x51203, x73517, x49845);
  nand n51204(x51204, x73597, x49815);
  nand n51206(x51206, x73592, x49817);
  nand n51208(x51208, x73587, x49819);
  nand n51210(x51210, x73582, x49821);
  nand n51212(x51212, x73577, x49823);
  nand n51214(x51214, x73572, x49825);
  nand n51216(x51216, x73567, x49827);
  nand n51218(x51218, x73562, x49829);
  nand n51220(x51220, x73557, x49831);
  nand n51222(x51222, x73552, x49833);
  nand n51224(x51224, x73547, x49835);
  nand n51226(x51226, x73542, x49837);
  nand n51228(x51228, x73537, x49839);
  nand n51230(x51230, x73532, x49841);
  nand n51232(x51232, x73527, x49843);
  nand n51234(x51234, x73522, x49845);
  nand n51236(x51236, x73517, x49847);
  nand n51238(x51238, x73602, x49815);
  nand n51240(x51240, x73597, x49817);
  nand n51242(x51242, x73592, x49819);
  nand n51244(x51244, x73587, x49821);
  nand n51246(x51246, x73582, x49823);
  nand n51248(x51248, x73577, x49825);
  nand n51250(x51250, x73572, x49827);
  nand n51252(x51252, x73567, x49829);
  nand n51254(x51254, x73562, x49831);
  nand n51256(x51256, x73557, x49833);
  nand n51258(x51258, x73552, x49835);
  nand n51260(x51260, x73547, x49837);
  nand n51262(x51262, x73542, x49839);
  nand n51264(x51264, x73537, x49841);
  nand n51266(x51266, x73532, x49843);
  nand n51268(x51268, x73527, x49845);
  nand n51270(x51270, x73522, x49847);
  nand n51272(x51272, x73517, x49849);
  nand n51274(x51274, x73607, x49815);
  nand n51276(x51276, x73602, x49817);
  nand n51278(x51278, x73597, x49819);
  nand n51280(x51280, x73592, x49821);
  nand n51282(x51282, x73587, x49823);
  nand n51284(x51284, x73582, x49825);
  nand n51286(x51286, x73577, x49827);
  nand n51288(x51288, x73572, x49829);
  nand n51290(x51290, x73567, x49831);
  nand n51292(x51292, x73562, x49833);
  nand n51294(x51294, x73557, x49835);
  nand n51296(x51296, x73552, x49837);
  nand n51298(x51298, x73547, x49839);
  nand n51300(x51300, x73542, x49841);
  nand n51302(x51302, x73537, x49843);
  nand n51304(x51304, x73532, x49845);
  nand n51306(x51306, x73527, x49847);
  nand n51308(x51308, x73522, x49849);
  nand n51310(x51310, x73517, x49851);
  nand n51311(x51311, x73612, x49815);
  nand n51313(x51313, x73607, x49817);
  nand n51315(x51315, x73602, x49819);
  nand n51317(x51317, x73597, x49821);
  nand n51319(x51319, x73592, x49823);
  nand n51321(x51321, x73587, x49825);
  nand n51323(x51323, x73582, x49827);
  nand n51325(x51325, x73577, x49829);
  nand n51327(x51327, x73572, x49831);
  nand n51329(x51329, x73567, x49833);
  nand n51331(x51331, x73562, x49835);
  nand n51333(x51333, x73557, x49837);
  nand n51335(x51335, x73552, x49839);
  nand n51337(x51337, x73547, x49841);
  nand n51339(x51339, x73542, x49843);
  nand n51341(x51341, x73537, x49845);
  nand n51343(x51343, x73532, x49847);
  nand n51345(x51345, x73527, x49849);
  nand n51347(x51347, x73522, x49851);
  nand n51349(x51349, x73517, x49853);
  nand n51351(x51351, x73617, x49815);
  nand n51353(x51353, x73612, x49817);
  nand n51355(x51355, x73607, x49819);
  nand n51357(x51357, x73602, x49821);
  nand n51359(x51359, x73597, x49823);
  nand n51361(x51361, x73592, x49825);
  nand n51363(x51363, x73587, x49827);
  nand n51365(x51365, x73582, x49829);
  nand n51367(x51367, x73577, x49831);
  nand n51369(x51369, x73572, x49833);
  nand n51371(x51371, x73567, x49835);
  nand n51373(x51373, x73562, x49837);
  nand n51375(x51375, x73557, x49839);
  nand n51377(x51377, x73552, x49841);
  nand n51379(x51379, x73547, x49843);
  nand n51381(x51381, x73542, x49845);
  nand n51383(x51383, x73537, x49847);
  nand n51385(x51385, x73532, x49849);
  nand n51387(x51387, x73527, x49851);
  nand n51389(x51389, x73522, x49853);
  nand n51391(x51391, x73517, x49855);
  nand n51393(x51393, x73622, x49815);
  nand n51395(x51395, x73617, x49817);
  nand n51397(x51397, x73612, x49819);
  nand n51399(x51399, x73607, x49821);
  nand n51401(x51401, x73602, x49823);
  nand n51403(x51403, x73597, x49825);
  nand n51405(x51405, x73592, x49827);
  nand n51407(x51407, x73587, x49829);
  nand n51409(x51409, x73582, x49831);
  nand n51411(x51411, x73577, x49833);
  nand n51413(x51413, x73572, x49835);
  nand n51415(x51415, x73567, x49837);
  nand n51417(x51417, x73562, x49839);
  nand n51419(x51419, x73557, x49841);
  nand n51421(x51421, x73552, x49843);
  nand n51423(x51423, x73547, x49845);
  nand n51425(x51425, x73542, x49847);
  nand n51427(x51427, x73537, x49849);
  nand n51429(x51429, x73532, x49851);
  nand n51431(x51431, x73527, x49853);
  nand n51433(x51433, x73522, x49855);
  nand n51435(x51435, x73517, x49857);
  nand n51436(x51436, x73627, x49815);
  nand n51438(x51438, x73622, x49817);
  nand n51440(x51440, x73617, x49819);
  nand n51442(x51442, x73612, x49821);
  nand n51444(x51444, x73607, x49823);
  nand n51446(x51446, x73602, x49825);
  nand n51448(x51448, x73597, x49827);
  nand n51450(x51450, x73592, x49829);
  nand n51452(x51452, x73587, x49831);
  nand n51454(x51454, x73582, x49833);
  nand n51456(x51456, x73577, x49835);
  nand n51458(x51458, x73572, x49837);
  nand n51460(x51460, x73567, x49839);
  nand n51462(x51462, x73562, x49841);
  nand n51464(x51464, x73557, x49843);
  nand n51466(x51466, x73552, x49845);
  nand n51468(x51468, x73547, x49847);
  nand n51470(x51470, x73542, x49849);
  nand n51472(x51472, x73537, x49851);
  nand n51474(x51474, x73532, x49853);
  nand n51476(x51476, x73527, x49855);
  nand n51478(x51478, x73522, x49857);
  nand n51480(x51480, x73517, x49859);
  nand n51482(x51482, x73632, x49815);
  nand n51484(x51484, x73627, x49817);
  nand n51486(x51486, x73622, x49819);
  nand n51488(x51488, x73617, x49821);
  nand n51490(x51490, x73612, x49823);
  nand n51492(x51492, x73607, x49825);
  nand n51494(x51494, x73602, x49827);
  nand n51496(x51496, x73597, x49829);
  nand n51498(x51498, x73592, x49831);
  nand n51500(x51500, x73587, x49833);
  nand n51502(x51502, x73582, x49835);
  nand n51504(x51504, x73577, x49837);
  nand n51506(x51506, x73572, x49839);
  nand n51508(x51508, x73567, x49841);
  nand n51510(x51510, x73562, x49843);
  nand n51512(x51512, x73557, x49845);
  nand n51514(x51514, x73552, x49847);
  nand n51516(x51516, x73547, x49849);
  nand n51518(x51518, x73542, x49851);
  nand n51520(x51520, x73537, x49853);
  nand n51522(x51522, x73532, x49855);
  nand n51524(x51524, x73527, x49857);
  nand n51526(x51526, x73522, x49859);
  nand n51528(x51528, x73517, x49861);
  nand n51530(x51530, x73637, x49815);
  nand n51532(x51532, x73632, x49817);
  nand n51534(x51534, x73627, x49819);
  nand n51536(x51536, x73622, x49821);
  nand n51538(x51538, x73617, x49823);
  nand n51540(x51540, x73612, x49825);
  nand n51542(x51542, x73607, x49827);
  nand n51544(x51544, x73602, x49829);
  nand n51546(x51546, x73597, x49831);
  nand n51548(x51548, x73592, x49833);
  nand n51550(x51550, x73587, x49835);
  nand n51552(x51552, x73582, x49837);
  nand n51554(x51554, x73577, x49839);
  nand n51556(x51556, x73572, x49841);
  nand n51558(x51558, x73567, x49843);
  nand n51560(x51560, x73562, x49845);
  nand n51562(x51562, x73557, x49847);
  nand n51564(x51564, x73552, x49849);
  nand n51566(x51566, x73547, x49851);
  nand n51568(x51568, x73542, x49853);
  nand n51570(x51570, x73537, x49855);
  nand n51572(x51572, x73532, x49857);
  nand n51574(x51574, x73527, x49859);
  nand n51576(x51576, x73522, x49861);
  nand n51578(x51578, x73517, x49863);
  nand n51579(x51579, x73642, x49815);
  nand n51581(x51581, x73637, x49817);
  nand n51583(x51583, x73632, x49819);
  nand n51585(x51585, x73627, x49821);
  nand n51587(x51587, x73622, x49823);
  nand n51589(x51589, x73617, x49825);
  nand n51591(x51591, x73612, x49827);
  nand n51593(x51593, x73607, x49829);
  nand n51595(x51595, x73602, x49831);
  nand n51597(x51597, x73597, x49833);
  nand n51599(x51599, x73592, x49835);
  nand n51601(x51601, x73587, x49837);
  nand n51603(x51603, x73582, x49839);
  nand n51605(x51605, x73577, x49841);
  nand n51607(x51607, x73572, x49843);
  nand n51609(x51609, x73567, x49845);
  nand n51611(x51611, x73562, x49847);
  nand n51613(x51613, x73557, x49849);
  nand n51615(x51615, x73552, x49851);
  nand n51617(x51617, x73547, x49853);
  nand n51619(x51619, x73542, x49855);
  nand n51621(x51621, x73537, x49857);
  nand n51623(x51623, x73532, x49859);
  nand n51625(x51625, x73527, x49861);
  nand n51627(x51627, x73522, x49863);
  nand n51629(x51629, x73517, x49865);
  nand n51631(x51631, x73647, x49815);
  nand n51633(x51633, x73642, x49817);
  nand n51635(x51635, x73637, x49819);
  nand n51637(x51637, x73632, x49821);
  nand n51639(x51639, x73627, x49823);
  nand n51641(x51641, x73622, x49825);
  nand n51643(x51643, x73617, x49827);
  nand n51645(x51645, x73612, x49829);
  nand n51647(x51647, x73607, x49831);
  nand n51649(x51649, x73602, x49833);
  nand n51651(x51651, x73597, x49835);
  nand n51653(x51653, x73592, x49837);
  nand n51655(x51655, x73587, x49839);
  nand n51657(x51657, x73582, x49841);
  nand n51659(x51659, x73577, x49843);
  nand n51661(x51661, x73572, x49845);
  nand n51663(x51663, x73567, x49847);
  nand n51665(x51665, x73562, x49849);
  nand n51667(x51667, x73557, x49851);
  nand n51669(x51669, x73552, x49853);
  nand n51671(x51671, x73547, x49855);
  nand n51673(x51673, x73542, x49857);
  nand n51675(x51675, x73537, x49859);
  nand n51677(x51677, x73532, x49861);
  nand n51679(x51679, x73527, x49863);
  nand n51681(x51681, x73522, x49865);
  nand n51683(x51683, x73517, x49867);
  nand n51685(x51685, x73652, x49815);
  nand n51687(x51687, x73647, x49817);
  nand n51689(x51689, x73642, x49819);
  nand n51691(x51691, x73637, x49821);
  nand n51693(x51693, x73632, x49823);
  nand n51695(x51695, x73627, x49825);
  nand n51697(x51697, x73622, x49827);
  nand n51699(x51699, x73617, x49829);
  nand n51701(x51701, x73612, x49831);
  nand n51703(x51703, x73607, x49833);
  nand n51705(x51705, x73602, x49835);
  nand n51707(x51707, x73597, x49837);
  nand n51709(x51709, x73592, x49839);
  nand n51711(x51711, x73587, x49841);
  nand n51713(x51713, x73582, x49843);
  nand n51715(x51715, x73577, x49845);
  nand n51717(x51717, x73572, x49847);
  nand n51719(x51719, x73567, x49849);
  nand n51721(x51721, x73562, x49851);
  nand n51723(x51723, x73557, x49853);
  nand n51725(x51725, x73552, x49855);
  nand n51727(x51727, x73547, x49857);
  nand n51729(x51729, x73542, x49859);
  nand n51731(x51731, x73537, x49861);
  nand n51733(x51733, x73532, x49863);
  nand n51735(x51735, x73527, x49865);
  nand n51737(x51737, x73522, x49867);
  nand n51739(x51739, x73517, x49869);
  nand n51740(x51740, x73657, x49815);
  nand n51742(x51742, x73652, x49817);
  nand n51744(x51744, x73647, x49819);
  nand n51746(x51746, x73642, x49821);
  nand n51748(x51748, x73637, x49823);
  nand n51750(x51750, x73632, x49825);
  nand n51752(x51752, x73627, x49827);
  nand n51754(x51754, x73622, x49829);
  nand n51756(x51756, x73617, x49831);
  nand n51758(x51758, x73612, x49833);
  nand n51760(x51760, x73607, x49835);
  nand n51762(x51762, x73602, x49837);
  nand n51764(x51764, x73597, x49839);
  nand n51766(x51766, x73592, x49841);
  nand n51768(x51768, x73587, x49843);
  nand n51770(x51770, x73582, x49845);
  nand n51772(x51772, x73577, x49847);
  nand n51774(x51774, x73572, x49849);
  nand n51776(x51776, x73567, x49851);
  nand n51778(x51778, x73562, x49853);
  nand n51780(x51780, x73557, x49855);
  nand n51782(x51782, x73552, x49857);
  nand n51784(x51784, x73547, x49859);
  nand n51786(x51786, x73542, x49861);
  nand n51788(x51788, x73537, x49863);
  nand n51790(x51790, x73532, x49865);
  nand n51792(x51792, x73527, x49867);
  nand n51794(x51794, x73522, x49869);
  nand n51796(x51796, x73517, x49871);
  nand n51798(x51798, x73662, x49815);
  nand n51800(x51800, x73657, x49817);
  nand n51802(x51802, x73652, x49819);
  nand n51804(x51804, x73647, x49821);
  nand n51806(x51806, x73642, x49823);
  nand n51808(x51808, x73637, x49825);
  nand n51810(x51810, x73632, x49827);
  nand n51812(x51812, x73627, x49829);
  nand n51814(x51814, x73622, x49831);
  nand n51816(x51816, x73617, x49833);
  nand n51818(x51818, x73612, x49835);
  nand n51820(x51820, x73607, x49837);
  nand n51822(x51822, x73602, x49839);
  nand n51824(x51824, x73597, x49841);
  nand n51826(x51826, x73592, x49843);
  nand n51828(x51828, x73587, x49845);
  nand n51830(x51830, x73582, x49847);
  nand n51832(x51832, x73577, x49849);
  nand n51834(x51834, x73572, x49851);
  nand n51836(x51836, x73567, x49853);
  nand n51838(x51838, x73562, x49855);
  nand n51840(x51840, x73557, x49857);
  nand n51842(x51842, x73552, x49859);
  nand n51844(x51844, x73547, x49861);
  nand n51846(x51846, x73542, x49863);
  nand n51848(x51848, x73537, x49865);
  nand n51850(x51850, x73532, x49867);
  nand n51852(x51852, x73527, x49869);
  nand n51854(x51854, x73522, x49871);
  nand n51856(x51856, x73517, x49873);
  nand n51858(x51858, x73667, x49815);
  nand n51860(x51860, x73662, x49817);
  nand n51862(x51862, x73657, x49819);
  nand n51864(x51864, x73652, x49821);
  nand n51866(x51866, x73647, x49823);
  nand n51868(x51868, x73642, x49825);
  nand n51870(x51870, x73637, x49827);
  nand n51872(x51872, x73632, x49829);
  nand n51874(x51874, x73627, x49831);
  nand n51876(x51876, x73622, x49833);
  nand n51878(x51878, x73617, x49835);
  nand n51880(x51880, x73612, x49837);
  nand n51882(x51882, x73607, x49839);
  nand n51884(x51884, x73602, x49841);
  nand n51886(x51886, x73597, x49843);
  nand n51888(x51888, x73592, x49845);
  nand n51890(x51890, x73587, x49847);
  nand n51892(x51892, x73582, x49849);
  nand n51894(x51894, x73577, x49851);
  nand n51896(x51896, x73572, x49853);
  nand n51898(x51898, x73567, x49855);
  nand n51900(x51900, x73562, x49857);
  nand n51902(x51902, x73557, x49859);
  nand n51904(x51904, x73552, x49861);
  nand n51906(x51906, x73547, x49863);
  nand n51908(x51908, x73542, x49865);
  nand n51910(x51910, x73537, x49867);
  nand n51912(x51912, x73532, x49869);
  nand n51914(x51914, x73527, x49871);
  nand n51916(x51916, x73522, x49873);
  nand n51918(x51918, x73517, x49875);
  nand n51919(x51919, x73672, x49815);
  nand n51921(x51921, x73667, x49817);
  nand n51923(x51923, x73662, x49819);
  nand n51925(x51925, x73657, x49821);
  nand n51927(x51927, x73652, x49823);
  nand n51929(x51929, x73647, x49825);
  nand n51931(x51931, x73642, x49827);
  nand n51933(x51933, x73637, x49829);
  nand n51935(x51935, x73632, x49831);
  nand n51937(x51937, x73627, x49833);
  nand n51939(x51939, x73622, x49835);
  nand n51941(x51941, x73617, x49837);
  nand n51943(x51943, x73612, x49839);
  nand n51945(x51945, x73607, x49841);
  nand n51947(x51947, x73602, x49843);
  nand n51949(x51949, x73597, x49845);
  nand n51951(x51951, x73592, x49847);
  nand n51953(x51953, x73587, x49849);
  nand n51955(x51955, x73582, x49851);
  nand n51957(x51957, x73577, x49853);
  nand n51959(x51959, x73572, x49855);
  nand n51961(x51961, x73567, x49857);
  nand n51963(x51963, x73562, x49859);
  nand n51965(x51965, x73557, x49861);
  nand n51967(x51967, x73552, x49863);
  nand n51969(x51969, x73547, x49865);
  nand n51971(x51971, x73542, x49867);
  nand n51973(x51973, x73537, x49869);
  nand n51975(x51975, x73532, x49871);
  nand n51977(x51977, x73527, x49873);
  nand n51979(x51979, x73522, x49875);
  nand n51981(x51981, x73517, x49877);
  nand n51983(x51983, x50940, x50942);
  nand n51984(x51984, x50939, x50941);
  nand n51985(x51985, x51984, x51983);
  nand n51986(x51986, x50944, x50946);
  nand n51987(x51987, x50943, x50945);
  nand n51988(x51988, x51987, x51986);
  nand n51990(x51990, x50948, x51989);
  nand n51991(x51991, x50947, x51988);
  nand n51992(x51992, x51991, x51990);
  nand n51993(x51993, x51986, x51990);
  nand n51994(x51994, x50950, x50952);
  nand n51995(x51995, x50949, x50951);
  nand n51996(x51996, x51995, x51994);
  nand n51998(x51998, x50954, x51997);
  nand n51999(x51999, x50953, x51996);
  nand n52000(x52000, x51999, x51998);
  nand n52001(x52001, x51994, x51998);
  nand n52002(x52002, x50957, x50959);
  nand n52003(x52003, x50956, x50958);
  nand n52004(x52004, x52003, x52002);
  nand n52006(x52006, x50961, x52005);
  nand n52007(x52007, x50960, x52004);
  nand n52008(x52008, x52007, x52006);
  nand n52009(x52009, x52002, x52006);
  nand n52010(x52010, x50963, x50965);
  nand n52011(x52011, x50962, x50964);
  nand n52012(x52012, x52011, x52010);
  nand n52013(x52013, x50967, x50969);
  nand n52014(x52014, x50966, x50968);
  nand n52015(x52015, x52014, x52013);
  nand n52017(x52017, x50971, x52016);
  nand n52018(x52018, x50970, x52015);
  nand n52019(x52019, x52018, x52017);
  nand n52020(x52020, x52013, x52017);
  nand n52021(x52021, x50973, x50975);
  nand n52022(x52022, x50972, x50974);
  nand n52023(x52023, x52022, x52021);
  nand n52025(x52025, x50977, x52024);
  nand n52026(x52026, x50976, x52023);
  nand n52027(x52027, x52026, x52025);
  nand n52028(x52028, x52021, x52025);
  nand n52029(x52029, x50979, x50981);
  nand n52030(x52030, x50978, x50980);
  nand n52031(x52031, x52030, x52029);
  nand n52033(x52033, x50983, x52032);
  nand n52034(x52034, x50982, x52031);
  nand n52035(x52035, x52034, x52033);
  nand n52036(x52036, x52029, x52033);
  nand n52037(x52037, x50985, x50987);
  nand n52038(x52038, x50984, x50986);
  nand n52039(x52039, x52038, x52037);
  nand n52041(x52041, x50989, x52040);
  nand n52042(x52042, x50988, x52039);
  nand n52043(x52043, x52042, x52041);
  nand n52045(x52045, x52037, x52041);
  nand n52046(x52046, x50992, x50994);
  nand n52047(x52047, x50991, x50993);
  nand n52048(x52048, x52047, x52046);
  nand n52050(x52050, x50996, x52049);
  nand n52051(x52051, x50995, x52048);
  nand n52052(x52052, x52051, x52050);
  nand n52053(x52053, x52046, x52050);
  nand n52054(x52054, x50998, x51000);
  nand n52055(x52055, x50997, x50999);
  nand n52056(x52056, x52055, x52054);
  nand n52058(x52058, x51002, x52057);
  nand n52059(x52059, x51001, x52056);
  nand n52060(x52060, x52059, x52058);
  nand n52062(x52062, x52054, x52058);
  nand n52063(x52063, x51004, x51006);
  nand n52064(x52064, x51003, x51005);
  nand n52065(x52065, x52064, x52063);
  nand n52066(x52066, x51008, x51010);
  nand n52067(x52067, x51007, x51009);
  nand n52068(x52068, x52067, x52066);
  nand n52070(x52070, x51012, x52069);
  nand n52071(x52071, x51011, x52068);
  nand n52072(x52072, x52071, x52070);
  nand n52073(x52073, x52066, x52070);
  nand n52074(x52074, x51014, x51016);
  nand n52075(x52075, x51013, x51015);
  nand n52076(x52076, x52075, x52074);
  nand n52078(x52078, x51018, x52077);
  nand n52079(x52079, x51017, x52076);
  nand n52080(x52080, x52079, x52078);
  nand n52082(x52082, x52074, x52078);
  nand n52083(x52083, x51020, x51022);
  nand n52084(x52084, x51019, x51021);
  nand n52085(x52085, x52084, x52083);
  nand n52087(x52087, x51024, x52086);
  nand n52088(x52088, x51023, x52085);
  nand n52089(x52089, x52088, x52087);
  nand n52091(x52091, x52083, x52087);
  nand n52092(x52092, x51026, x51028);
  nand n52093(x52093, x51025, x51027);
  nand n52094(x52094, x52093, x52092);
  nand n52096(x52096, x51030, x52095);
  nand n52097(x52097, x51029, x52094);
  nand n52098(x52098, x52097, x52096);
  nand n52099(x52099, x52092, x52096);
  nand n52100(x52100, x51032, x51034);
  nand n52101(x52101, x51031, x51033);
  nand n52102(x52102, x52101, x52100);
  nand n52104(x52104, x51036, x52103);
  nand n52105(x52105, x51035, x52102);
  nand n52106(x52106, x52105, x52104);
  nand n52108(x52108, x52100, x52104);
  nand n52109(x52109, x51038, x51040);
  nand n52110(x52110, x51037, x51039);
  nand n52111(x52111, x52110, x52109);
  nand n52113(x52113, x51042, x52112);
  nand n52114(x52114, x51041, x52111);
  nand n52115(x52115, x52114, x52113);
  nand n52117(x52117, x52109, x52113);
  nand n52118(x52118, x51045, x51047);
  nand n52119(x52119, x51044, x51046);
  nand n52120(x52120, x52119, x52118);
  nand n52122(x52122, x51049, x52121);
  nand n52123(x52123, x51048, x52120);
  nand n52124(x52124, x52123, x52122);
  nand n52125(x52125, x52118, x52122);
  nand n52126(x52126, x51051, x51053);
  nand n52127(x52127, x51050, x51052);
  nand n52128(x52128, x52127, x52126);
  nand n52130(x52130, x51055, x52129);
  nand n52131(x52131, x51054, x52128);
  nand n52132(x52132, x52131, x52130);
  nand n52134(x52134, x52126, x52130);
  nand n52135(x52135, x51057, x51059);
  nand n52136(x52136, x51056, x51058);
  nand n52137(x52137, x52136, x52135);
  nand n52139(x52139, x51061, x52138);
  nand n52140(x52140, x51060, x52137);
  nand n52141(x52141, x52140, x52139);
  nand n52143(x52143, x52135, x52139);
  nand n52144(x52144, x51063, x51065);
  nand n52145(x52145, x51062, x51064);
  nand n52146(x52146, x52145, x52144);
  nand n52147(x52147, x51067, x51069);
  nand n52148(x52148, x51066, x51068);
  nand n52149(x52149, x52148, x52147);
  nand n52151(x52151, x51071, x52150);
  nand n52152(x52152, x51070, x52149);
  nand n52153(x52153, x52152, x52151);
  nand n52154(x52154, x52147, x52151);
  nand n52155(x52155, x51073, x51075);
  nand n52156(x52156, x51072, x51074);
  nand n52157(x52157, x52156, x52155);
  nand n52159(x52159, x51077, x52158);
  nand n52160(x52160, x51076, x52157);
  nand n52161(x52161, x52160, x52159);
  nand n52163(x52163, x52155, x52159);
  nand n52164(x52164, x51079, x51081);
  nand n52165(x52165, x51078, x51080);
  nand n52166(x52166, x52165, x52164);
  nand n52168(x52168, x51083, x52167);
  nand n52169(x52169, x51082, x52166);
  nand n52170(x52170, x52169, x52168);
  nand n52172(x52172, x52164, x52168);
  nand n52173(x52173, x51085, x51087);
  nand n52174(x52174, x51084, x51086);
  nand n52175(x52175, x52174, x52173);
  nand n52177(x52177, x51089, x52176);
  nand n52178(x52178, x51088, x52175);
  nand n52179(x52179, x52178, x52177);
  nand n52181(x52181, x52173, x52177);
  nand n52182(x52182, x51091, x51093);
  nand n52183(x52183, x51090, x51092);
  nand n52184(x52184, x52183, x52182);
  nand n52186(x52186, x51095, x52185);
  nand n52187(x52187, x51094, x52184);
  nand n52188(x52188, x52187, x52186);
  nand n52189(x52189, x52182, x52186);
  nand n52190(x52190, x51097, x51099);
  nand n52191(x52191, x51096, x51098);
  nand n52192(x52192, x52191, x52190);
  nand n52194(x52194, x51101, x52193);
  nand n52195(x52195, x51100, x52192);
  nand n52196(x52196, x52195, x52194);
  nand n52198(x52198, x52190, x52194);
  nand n52199(x52199, x51103, x51105);
  nand n52200(x52200, x51102, x51104);
  nand n52201(x52201, x52200, x52199);
  nand n52203(x52203, x51107, x52202);
  nand n52204(x52204, x51106, x52201);
  nand n52205(x52205, x52204, x52203);
  nand n52207(x52207, x52199, x52203);
  nand n52208(x52208, x51109, x51111);
  nand n52209(x52209, x51108, x51110);
  nand n52210(x52210, x52209, x52208);
  nand n52212(x52212, x51113, x52211);
  nand n52213(x52213, x51112, x52210);
  nand n52214(x52214, x52213, x52212);
  nand n52216(x52216, x52208, x52212);
  nand n52217(x52217, x51116, x51118);
  nand n52218(x52218, x51115, x51117);
  nand n52219(x52219, x52218, x52217);
  nand n52221(x52221, x51120, x52220);
  nand n52222(x52222, x51119, x52219);
  nand n52223(x52223, x52222, x52221);
  nand n52224(x52224, x52217, x52221);
  nand n52225(x52225, x51122, x51124);
  nand n52226(x52226, x51121, x51123);
  nand n52227(x52227, x52226, x52225);
  nand n52229(x52229, x51126, x52228);
  nand n52230(x52230, x51125, x52227);
  nand n52231(x52231, x52230, x52229);
  nand n52233(x52233, x52225, x52229);
  nand n52234(x52234, x51128, x51130);
  nand n52235(x52235, x51127, x51129);
  nand n52236(x52236, x52235, x52234);
  nand n52238(x52238, x51132, x52237);
  nand n52239(x52239, x51131, x52236);
  nand n52240(x52240, x52239, x52238);
  nand n52242(x52242, x52234, x52238);
  nand n52243(x52243, x51134, x51136);
  nand n52244(x52244, x51133, x51135);
  nand n52245(x52245, x52244, x52243);
  nand n52247(x52247, x51138, x52246);
  nand n52248(x52248, x51137, x52245);
  nand n52249(x52249, x52248, x52247);
  nand n52251(x52251, x52243, x52247);
  nand n52252(x52252, x51140, x51142);
  nand n52253(x52253, x51139, x51141);
  nand n52254(x52254, x52253, x52252);
  nand n52255(x52255, x51144, x51146);
  nand n52256(x52256, x51143, x51145);
  nand n52257(x52257, x52256, x52255);
  nand n52259(x52259, x51148, x52258);
  nand n52260(x52260, x51147, x52257);
  nand n52261(x52261, x52260, x52259);
  nand n52262(x52262, x52255, x52259);
  nand n52263(x52263, x51150, x51152);
  nand n52264(x52264, x51149, x51151);
  nand n52265(x52265, x52264, x52263);
  nand n52267(x52267, x51154, x52266);
  nand n52268(x52268, x51153, x52265);
  nand n52269(x52269, x52268, x52267);
  nand n52271(x52271, x52263, x52267);
  nand n52272(x52272, x51156, x51158);
  nand n52273(x52273, x51155, x51157);
  nand n52274(x52274, x52273, x52272);
  nand n52276(x52276, x51160, x52275);
  nand n52277(x52277, x51159, x52274);
  nand n52278(x52278, x52277, x52276);
  nand n52280(x52280, x52272, x52276);
  nand n52281(x52281, x51162, x51164);
  nand n52282(x52282, x51161, x51163);
  nand n52283(x52283, x52282, x52281);
  nand n52285(x52285, x51166, x52284);
  nand n52286(x52286, x51165, x52283);
  nand n52287(x52287, x52286, x52285);
  nand n52289(x52289, x52281, x52285);
  nand n52290(x52290, x51168, x51170);
  nand n52291(x52291, x51167, x51169);
  nand n52292(x52292, x52291, x52290);
  nand n52294(x52294, x51172, x52293);
  nand n52295(x52295, x51171, x52292);
  nand n52296(x52296, x52295, x52294);
  nand n52297(x52297, x52290, x52294);
  nand n52298(x52298, x51174, x51176);
  nand n52299(x52299, x51173, x51175);
  nand n52300(x52300, x52299, x52298);
  nand n52302(x52302, x51178, x52301);
  nand n52303(x52303, x51177, x52300);
  nand n52304(x52304, x52303, x52302);
  nand n52305(x52305, x52298, x52302);
  nand n52306(x52306, x51180, x51182);
  nand n52307(x52307, x51179, x51181);
  nand n52308(x52308, x52307, x52306);
  nand n52310(x52310, x51184, x52309);
  nand n52311(x52311, x51183, x52308);
  nand n52312(x52312, x52311, x52310);
  nand n52314(x52314, x52306, x52310);
  nand n52315(x52315, x51186, x51188);
  nand n52316(x52316, x51185, x51187);
  nand n52317(x52317, x52316, x52315);
  nand n52319(x52319, x51190, x52318);
  nand n52320(x52320, x51189, x52317);
  nand n52321(x52321, x52320, x52319);
  nand n52323(x52323, x52315, x52319);
  nand n52324(x52324, x51192, x51194);
  nand n52325(x52325, x51191, x51193);
  nand n52326(x52326, x52325, x52324);
  nand n52328(x52328, x51196, x52327);
  nand n52329(x52329, x51195, x52326);
  nand n52330(x52330, x52329, x52328);
  nand n52332(x52332, x52324, x52328);
  nand n52333(x52333, x51198, x51200);
  nand n52334(x52334, x51197, x51199);
  nand n52335(x52335, x52334, x52333);
  nand n52337(x52337, x51202, x52336);
  nand n52338(x52338, x51201, x52335);
  nand n52339(x52339, x52338, x52337);
  nand n52341(x52341, x52333, x52337);
  nand n52342(x52342, x51205, x51207);
  nand n52343(x52343, x51204, x51206);
  nand n52344(x52344, x52343, x52342);
  nand n52346(x52346, x51209, x52345);
  nand n52347(x52347, x51208, x52344);
  nand n52348(x52348, x52347, x52346);
  nand n52349(x52349, x52342, x52346);
  nand n52350(x52350, x51211, x51213);
  nand n52351(x52351, x51210, x51212);
  nand n52352(x52352, x52351, x52350);
  nand n52354(x52354, x51215, x52353);
  nand n52355(x52355, x51214, x52352);
  nand n52356(x52356, x52355, x52354);
  nand n52358(x52358, x52350, x52354);
  nand n52359(x52359, x51217, x51219);
  nand n52360(x52360, x51216, x51218);
  nand n52361(x52361, x52360, x52359);
  nand n52363(x52363, x51221, x52362);
  nand n52364(x52364, x51220, x52361);
  nand n52365(x52365, x52364, x52363);
  nand n52367(x52367, x52359, x52363);
  nand n52368(x52368, x51223, x51225);
  nand n52369(x52369, x51222, x51224);
  nand n52370(x52370, x52369, x52368);
  nand n52372(x52372, x51227, x52371);
  nand n52373(x52373, x51226, x52370);
  nand n52374(x52374, x52373, x52372);
  nand n52376(x52376, x52368, x52372);
  nand n52377(x52377, x51229, x51231);
  nand n52378(x52378, x51228, x51230);
  nand n52379(x52379, x52378, x52377);
  nand n52381(x52381, x51233, x52380);
  nand n52382(x52382, x51232, x52379);
  nand n52383(x52383, x52382, x52381);
  nand n52385(x52385, x52377, x52381);
  nand n52386(x52386, x51235, x51237);
  nand n52387(x52387, x51234, x51236);
  nand n52388(x52388, x52387, x52386);
  nand n52389(x52389, x51239, x51241);
  nand n52390(x52390, x51238, x51240);
  nand n52391(x52391, x52390, x52389);
  nand n52393(x52393, x51243, x52392);
  nand n52394(x52394, x51242, x52391);
  nand n52395(x52395, x52394, x52393);
  nand n52396(x52396, x52389, x52393);
  nand n52397(x52397, x51245, x51247);
  nand n52398(x52398, x51244, x51246);
  nand n52399(x52399, x52398, x52397);
  nand n52401(x52401, x51249, x52400);
  nand n52402(x52402, x51248, x52399);
  nand n52403(x52403, x52402, x52401);
  nand n52405(x52405, x52397, x52401);
  nand n52406(x52406, x51251, x51253);
  nand n52407(x52407, x51250, x51252);
  nand n52408(x52408, x52407, x52406);
  nand n52410(x52410, x51255, x52409);
  nand n52411(x52411, x51254, x52408);
  nand n52412(x52412, x52411, x52410);
  nand n52414(x52414, x52406, x52410);
  nand n52415(x52415, x51257, x51259);
  nand n52416(x52416, x51256, x51258);
  nand n52417(x52417, x52416, x52415);
  nand n52419(x52419, x51261, x52418);
  nand n52420(x52420, x51260, x52417);
  nand n52421(x52421, x52420, x52419);
  nand n52423(x52423, x52415, x52419);
  nand n52424(x52424, x51263, x51265);
  nand n52425(x52425, x51262, x51264);
  nand n52426(x52426, x52425, x52424);
  nand n52428(x52428, x51267, x52427);
  nand n52429(x52429, x51266, x52426);
  nand n52430(x52430, x52429, x52428);
  nand n52432(x52432, x52424, x52428);
  nand n52433(x52433, x51269, x51271);
  nand n52434(x52434, x51268, x51270);
  nand n52435(x52435, x52434, x52433);
  nand n52437(x52437, x51273, x52436);
  nand n52438(x52438, x51272, x52435);
  nand n52439(x52439, x52438, x52437);
  nand n52441(x52441, x52433, x52437);
  nand n52442(x52442, x51275, x51277);
  nand n52443(x52443, x51274, x51276);
  nand n52444(x52444, x52443, x52442);
  nand n52446(x52446, x51279, x52445);
  nand n52447(x52447, x51278, x52444);
  nand n52448(x52448, x52447, x52446);
  nand n52449(x52449, x52442, x52446);
  nand n52450(x52450, x51281, x51283);
  nand n52451(x52451, x51280, x51282);
  nand n52452(x52452, x52451, x52450);
  nand n52454(x52454, x51285, x52453);
  nand n52455(x52455, x51284, x52452);
  nand n52456(x52456, x52455, x52454);
  nand n52458(x52458, x52450, x52454);
  nand n52459(x52459, x51287, x51289);
  nand n52460(x52460, x51286, x51288);
  nand n52461(x52461, x52460, x52459);
  nand n52463(x52463, x51291, x52462);
  nand n52464(x52464, x51290, x52461);
  nand n52465(x52465, x52464, x52463);
  nand n52467(x52467, x52459, x52463);
  nand n52468(x52468, x51293, x51295);
  nand n52469(x52469, x51292, x51294);
  nand n52470(x52470, x52469, x52468);
  nand n52472(x52472, x51297, x52471);
  nand n52473(x52473, x51296, x52470);
  nand n52474(x52474, x52473, x52472);
  nand n52476(x52476, x52468, x52472);
  nand n52477(x52477, x51299, x51301);
  nand n52478(x52478, x51298, x51300);
  nand n52479(x52479, x52478, x52477);
  nand n52481(x52481, x51303, x52480);
  nand n52482(x52482, x51302, x52479);
  nand n52483(x52483, x52482, x52481);
  nand n52485(x52485, x52477, x52481);
  nand n52486(x52486, x51305, x51307);
  nand n52487(x52487, x51304, x51306);
  nand n52488(x52488, x52487, x52486);
  nand n52490(x52490, x51309, x52489);
  nand n52491(x52491, x51308, x52488);
  nand n52492(x52492, x52491, x52490);
  nand n52494(x52494, x52486, x52490);
  nand n52495(x52495, x51312, x51314);
  nand n52496(x52496, x51311, x51313);
  nand n52497(x52497, x52496, x52495);
  nand n52499(x52499, x51316, x52498);
  nand n52500(x52500, x51315, x52497);
  nand n52501(x52501, x52500, x52499);
  nand n52502(x52502, x52495, x52499);
  nand n52503(x52503, x51318, x51320);
  nand n52504(x52504, x51317, x51319);
  nand n52505(x52505, x52504, x52503);
  nand n52507(x52507, x51322, x52506);
  nand n52508(x52508, x51321, x52505);
  nand n52509(x52509, x52508, x52507);
  nand n52511(x52511, x52503, x52507);
  nand n52512(x52512, x51324, x51326);
  nand n52513(x52513, x51323, x51325);
  nand n52514(x52514, x52513, x52512);
  nand n52516(x52516, x51328, x52515);
  nand n52517(x52517, x51327, x52514);
  nand n52518(x52518, x52517, x52516);
  nand n52520(x52520, x52512, x52516);
  nand n52521(x52521, x51330, x51332);
  nand n52522(x52522, x51329, x51331);
  nand n52523(x52523, x52522, x52521);
  nand n52525(x52525, x51334, x52524);
  nand n52526(x52526, x51333, x52523);
  nand n52527(x52527, x52526, x52525);
  nand n52529(x52529, x52521, x52525);
  nand n52530(x52530, x51336, x51338);
  nand n52531(x52531, x51335, x51337);
  nand n52532(x52532, x52531, x52530);
  nand n52534(x52534, x51340, x52533);
  nand n52535(x52535, x51339, x52532);
  nand n52536(x52536, x52535, x52534);
  nand n52538(x52538, x52530, x52534);
  nand n52539(x52539, x51342, x51344);
  nand n52540(x52540, x51341, x51343);
  nand n52541(x52541, x52540, x52539);
  nand n52543(x52543, x51346, x52542);
  nand n52544(x52544, x51345, x52541);
  nand n52545(x52545, x52544, x52543);
  nand n52547(x52547, x52539, x52543);
  nand n52548(x52548, x51348, x51350);
  nand n52549(x52549, x51347, x51349);
  nand n52550(x52550, x52549, x52548);
  nand n52551(x52551, x51352, x51354);
  nand n52552(x52552, x51351, x51353);
  nand n52553(x52553, x52552, x52551);
  nand n52555(x52555, x51356, x52554);
  nand n52556(x52556, x51355, x52553);
  nand n52557(x52557, x52556, x52555);
  nand n52558(x52558, x52551, x52555);
  nand n52559(x52559, x51358, x51360);
  nand n52560(x52560, x51357, x51359);
  nand n52561(x52561, x52560, x52559);
  nand n52563(x52563, x51362, x52562);
  nand n52564(x52564, x51361, x52561);
  nand n52565(x52565, x52564, x52563);
  nand n52567(x52567, x52559, x52563);
  nand n52568(x52568, x51364, x51366);
  nand n52569(x52569, x51363, x51365);
  nand n52570(x52570, x52569, x52568);
  nand n52572(x52572, x51368, x52571);
  nand n52573(x52573, x51367, x52570);
  nand n52574(x52574, x52573, x52572);
  nand n52576(x52576, x52568, x52572);
  nand n52577(x52577, x51370, x51372);
  nand n52578(x52578, x51369, x51371);
  nand n52579(x52579, x52578, x52577);
  nand n52581(x52581, x51374, x52580);
  nand n52582(x52582, x51373, x52579);
  nand n52583(x52583, x52582, x52581);
  nand n52585(x52585, x52577, x52581);
  nand n52586(x52586, x51376, x51378);
  nand n52587(x52587, x51375, x51377);
  nand n52588(x52588, x52587, x52586);
  nand n52590(x52590, x51380, x52589);
  nand n52591(x52591, x51379, x52588);
  nand n52592(x52592, x52591, x52590);
  nand n52594(x52594, x52586, x52590);
  nand n52595(x52595, x51382, x51384);
  nand n52596(x52596, x51381, x51383);
  nand n52597(x52597, x52596, x52595);
  nand n52599(x52599, x51386, x52598);
  nand n52600(x52600, x51385, x52597);
  nand n52601(x52601, x52600, x52599);
  nand n52603(x52603, x52595, x52599);
  nand n52604(x52604, x51388, x51390);
  nand n52605(x52605, x51387, x51389);
  nand n52606(x52606, x52605, x52604);
  nand n52608(x52608, x51392, x52607);
  nand n52609(x52609, x51391, x52606);
  nand n52610(x52610, x52609, x52608);
  nand n52612(x52612, x52604, x52608);
  nand n52613(x52613, x51394, x51396);
  nand n52614(x52614, x51393, x51395);
  nand n52615(x52615, x52614, x52613);
  nand n52617(x52617, x51398, x52616);
  nand n52618(x52618, x51397, x52615);
  nand n52619(x52619, x52618, x52617);
  nand n52620(x52620, x52613, x52617);
  nand n52621(x52621, x51400, x51402);
  nand n52622(x52622, x51399, x51401);
  nand n52623(x52623, x52622, x52621);
  nand n52625(x52625, x51404, x52624);
  nand n52626(x52626, x51403, x52623);
  nand n52627(x52627, x52626, x52625);
  nand n52629(x52629, x52621, x52625);
  nand n52630(x52630, x51406, x51408);
  nand n52631(x52631, x51405, x51407);
  nand n52632(x52632, x52631, x52630);
  nand n52634(x52634, x51410, x52633);
  nand n52635(x52635, x51409, x52632);
  nand n52636(x52636, x52635, x52634);
  nand n52638(x52638, x52630, x52634);
  nand n52639(x52639, x51412, x51414);
  nand n52640(x52640, x51411, x51413);
  nand n52641(x52641, x52640, x52639);
  nand n52643(x52643, x51416, x52642);
  nand n52644(x52644, x51415, x52641);
  nand n52645(x52645, x52644, x52643);
  nand n52647(x52647, x52639, x52643);
  nand n52648(x52648, x51418, x51420);
  nand n52649(x52649, x51417, x51419);
  nand n52650(x52650, x52649, x52648);
  nand n52652(x52652, x51422, x52651);
  nand n52653(x52653, x51421, x52650);
  nand n52654(x52654, x52653, x52652);
  nand n52656(x52656, x52648, x52652);
  nand n52657(x52657, x51424, x51426);
  nand n52658(x52658, x51423, x51425);
  nand n52659(x52659, x52658, x52657);
  nand n52661(x52661, x51428, x52660);
  nand n52662(x52662, x51427, x52659);
  nand n52663(x52663, x52662, x52661);
  nand n52665(x52665, x52657, x52661);
  nand n52666(x52666, x51430, x51432);
  nand n52667(x52667, x51429, x51431);
  nand n52668(x52668, x52667, x52666);
  nand n52670(x52670, x51434, x52669);
  nand n52671(x52671, x51433, x52668);
  nand n52672(x52672, x52671, x52670);
  nand n52674(x52674, x52666, x52670);
  nand n52675(x52675, x51437, x51439);
  nand n52676(x52676, x51436, x51438);
  nand n52677(x52677, x52676, x52675);
  nand n52679(x52679, x51441, x52678);
  nand n52680(x52680, x51440, x52677);
  nand n52681(x52681, x52680, x52679);
  nand n52682(x52682, x52675, x52679);
  nand n52683(x52683, x51443, x51445);
  nand n52684(x52684, x51442, x51444);
  nand n52685(x52685, x52684, x52683);
  nand n52687(x52687, x51447, x52686);
  nand n52688(x52688, x51446, x52685);
  nand n52689(x52689, x52688, x52687);
  nand n52691(x52691, x52683, x52687);
  nand n52692(x52692, x51449, x51451);
  nand n52693(x52693, x51448, x51450);
  nand n52694(x52694, x52693, x52692);
  nand n52696(x52696, x51453, x52695);
  nand n52697(x52697, x51452, x52694);
  nand n52698(x52698, x52697, x52696);
  nand n52700(x52700, x52692, x52696);
  nand n52701(x52701, x51455, x51457);
  nand n52702(x52702, x51454, x51456);
  nand n52703(x52703, x52702, x52701);
  nand n52705(x52705, x51459, x52704);
  nand n52706(x52706, x51458, x52703);
  nand n52707(x52707, x52706, x52705);
  nand n52709(x52709, x52701, x52705);
  nand n52710(x52710, x51461, x51463);
  nand n52711(x52711, x51460, x51462);
  nand n52712(x52712, x52711, x52710);
  nand n52714(x52714, x51465, x52713);
  nand n52715(x52715, x51464, x52712);
  nand n52716(x52716, x52715, x52714);
  nand n52718(x52718, x52710, x52714);
  nand n52719(x52719, x51467, x51469);
  nand n52720(x52720, x51466, x51468);
  nand n52721(x52721, x52720, x52719);
  nand n52723(x52723, x51471, x52722);
  nand n52724(x52724, x51470, x52721);
  nand n52725(x52725, x52724, x52723);
  nand n52727(x52727, x52719, x52723);
  nand n52728(x52728, x51473, x51475);
  nand n52729(x52729, x51472, x51474);
  nand n52730(x52730, x52729, x52728);
  nand n52732(x52732, x51477, x52731);
  nand n52733(x52733, x51476, x52730);
  nand n52734(x52734, x52733, x52732);
  nand n52736(x52736, x52728, x52732);
  nand n52737(x52737, x51479, x51481);
  nand n52738(x52738, x51478, x51480);
  nand n52739(x52739, x52738, x52737);
  nand n52740(x52740, x51483, x51485);
  nand n52741(x52741, x51482, x51484);
  nand n52742(x52742, x52741, x52740);
  nand n52744(x52744, x51487, x52743);
  nand n52745(x52745, x51486, x52742);
  nand n52746(x52746, x52745, x52744);
  nand n52747(x52747, x52740, x52744);
  nand n52748(x52748, x51489, x51491);
  nand n52749(x52749, x51488, x51490);
  nand n52750(x52750, x52749, x52748);
  nand n52752(x52752, x51493, x52751);
  nand n52753(x52753, x51492, x52750);
  nand n52754(x52754, x52753, x52752);
  nand n52756(x52756, x52748, x52752);
  nand n52757(x52757, x51495, x51497);
  nand n52758(x52758, x51494, x51496);
  nand n52759(x52759, x52758, x52757);
  nand n52761(x52761, x51499, x52760);
  nand n52762(x52762, x51498, x52759);
  nand n52763(x52763, x52762, x52761);
  nand n52765(x52765, x52757, x52761);
  nand n52766(x52766, x51501, x51503);
  nand n52767(x52767, x51500, x51502);
  nand n52768(x52768, x52767, x52766);
  nand n52770(x52770, x51505, x52769);
  nand n52771(x52771, x51504, x52768);
  nand n52772(x52772, x52771, x52770);
  nand n52774(x52774, x52766, x52770);
  nand n52775(x52775, x51507, x51509);
  nand n52776(x52776, x51506, x51508);
  nand n52777(x52777, x52776, x52775);
  nand n52779(x52779, x51511, x52778);
  nand n52780(x52780, x51510, x52777);
  nand n52781(x52781, x52780, x52779);
  nand n52783(x52783, x52775, x52779);
  nand n52784(x52784, x51513, x51515);
  nand n52785(x52785, x51512, x51514);
  nand n52786(x52786, x52785, x52784);
  nand n52788(x52788, x51517, x52787);
  nand n52789(x52789, x51516, x52786);
  nand n52790(x52790, x52789, x52788);
  nand n52792(x52792, x52784, x52788);
  nand n52793(x52793, x51519, x51521);
  nand n52794(x52794, x51518, x51520);
  nand n52795(x52795, x52794, x52793);
  nand n52797(x52797, x51523, x52796);
  nand n52798(x52798, x51522, x52795);
  nand n52799(x52799, x52798, x52797);
  nand n52801(x52801, x52793, x52797);
  nand n52802(x52802, x51525, x51527);
  nand n52803(x52803, x51524, x51526);
  nand n52804(x52804, x52803, x52802);
  nand n52806(x52806, x51529, x52805);
  nand n52807(x52807, x51528, x52804);
  nand n52808(x52808, x52807, x52806);
  nand n52809(x52809, x52802, x52806);
  nand n52810(x52810, x51531, x51533);
  nand n52811(x52811, x51530, x51532);
  nand n52812(x52812, x52811, x52810);
  nand n52814(x52814, x51535, x52813);
  nand n52815(x52815, x51534, x52812);
  nand n52816(x52816, x52815, x52814);
  nand n52817(x52817, x52810, x52814);
  nand n52818(x52818, x51537, x51539);
  nand n52819(x52819, x51536, x51538);
  nand n52820(x52820, x52819, x52818);
  nand n52822(x52822, x51541, x52821);
  nand n52823(x52823, x51540, x52820);
  nand n52824(x52824, x52823, x52822);
  nand n52826(x52826, x52818, x52822);
  nand n52827(x52827, x51543, x51545);
  nand n52828(x52828, x51542, x51544);
  nand n52829(x52829, x52828, x52827);
  nand n52831(x52831, x51547, x52830);
  nand n52832(x52832, x51546, x52829);
  nand n52833(x52833, x52832, x52831);
  nand n52835(x52835, x52827, x52831);
  nand n52836(x52836, x51549, x51551);
  nand n52837(x52837, x51548, x51550);
  nand n52838(x52838, x52837, x52836);
  nand n52840(x52840, x51553, x52839);
  nand n52841(x52841, x51552, x52838);
  nand n52842(x52842, x52841, x52840);
  nand n52844(x52844, x52836, x52840);
  nand n52845(x52845, x51555, x51557);
  nand n52846(x52846, x51554, x51556);
  nand n52847(x52847, x52846, x52845);
  nand n52849(x52849, x51559, x52848);
  nand n52850(x52850, x51558, x52847);
  nand n52851(x52851, x52850, x52849);
  nand n52853(x52853, x52845, x52849);
  nand n52854(x52854, x51561, x51563);
  nand n52855(x52855, x51560, x51562);
  nand n52856(x52856, x52855, x52854);
  nand n52858(x52858, x51565, x52857);
  nand n52859(x52859, x51564, x52856);
  nand n52860(x52860, x52859, x52858);
  nand n52862(x52862, x52854, x52858);
  nand n52863(x52863, x51567, x51569);
  nand n52864(x52864, x51566, x51568);
  nand n52865(x52865, x52864, x52863);
  nand n52867(x52867, x51571, x52866);
  nand n52868(x52868, x51570, x52865);
  nand n52869(x52869, x52868, x52867);
  nand n52871(x52871, x52863, x52867);
  nand n52872(x52872, x51573, x51575);
  nand n52873(x52873, x51572, x51574);
  nand n52874(x52874, x52873, x52872);
  nand n52876(x52876, x51577, x52875);
  nand n52877(x52877, x51576, x52874);
  nand n52878(x52878, x52877, x52876);
  nand n52880(x52880, x52872, x52876);
  nand n52881(x52881, x51580, x51582);
  nand n52882(x52882, x51579, x51581);
  nand n52883(x52883, x52882, x52881);
  nand n52885(x52885, x51584, x52884);
  nand n52886(x52886, x51583, x52883);
  nand n52887(x52887, x52886, x52885);
  nand n52888(x52888, x52881, x52885);
  nand n52889(x52889, x51586, x51588);
  nand n52890(x52890, x51585, x51587);
  nand n52891(x52891, x52890, x52889);
  nand n52893(x52893, x51590, x52892);
  nand n52894(x52894, x51589, x52891);
  nand n52895(x52895, x52894, x52893);
  nand n52897(x52897, x52889, x52893);
  nand n52898(x52898, x51592, x51594);
  nand n52899(x52899, x51591, x51593);
  nand n52900(x52900, x52899, x52898);
  nand n52902(x52902, x51596, x52901);
  nand n52903(x52903, x51595, x52900);
  nand n52904(x52904, x52903, x52902);
  nand n52906(x52906, x52898, x52902);
  nand n52907(x52907, x51598, x51600);
  nand n52908(x52908, x51597, x51599);
  nand n52909(x52909, x52908, x52907);
  nand n52911(x52911, x51602, x52910);
  nand n52912(x52912, x51601, x52909);
  nand n52913(x52913, x52912, x52911);
  nand n52915(x52915, x52907, x52911);
  nand n52916(x52916, x51604, x51606);
  nand n52917(x52917, x51603, x51605);
  nand n52918(x52918, x52917, x52916);
  nand n52920(x52920, x51608, x52919);
  nand n52921(x52921, x51607, x52918);
  nand n52922(x52922, x52921, x52920);
  nand n52924(x52924, x52916, x52920);
  nand n52925(x52925, x51610, x51612);
  nand n52926(x52926, x51609, x51611);
  nand n52927(x52927, x52926, x52925);
  nand n52929(x52929, x51614, x52928);
  nand n52930(x52930, x51613, x52927);
  nand n52931(x52931, x52930, x52929);
  nand n52933(x52933, x52925, x52929);
  nand n52934(x52934, x51616, x51618);
  nand n52935(x52935, x51615, x51617);
  nand n52936(x52936, x52935, x52934);
  nand n52938(x52938, x51620, x52937);
  nand n52939(x52939, x51619, x52936);
  nand n52940(x52940, x52939, x52938);
  nand n52942(x52942, x52934, x52938);
  nand n52943(x52943, x51622, x51624);
  nand n52944(x52944, x51621, x51623);
  nand n52945(x52945, x52944, x52943);
  nand n52947(x52947, x51626, x52946);
  nand n52948(x52948, x51625, x52945);
  nand n52949(x52949, x52948, x52947);
  nand n52951(x52951, x52943, x52947);
  nand n52952(x52952, x51628, x51630);
  nand n52953(x52953, x51627, x51629);
  nand n52954(x52954, x52953, x52952);
  nand n52955(x52955, x51632, x51634);
  nand n52956(x52956, x51631, x51633);
  nand n52957(x52957, x52956, x52955);
  nand n52959(x52959, x51636, x52958);
  nand n52960(x52960, x51635, x52957);
  nand n52961(x52961, x52960, x52959);
  nand n52962(x52962, x52955, x52959);
  nand n52963(x52963, x51638, x51640);
  nand n52964(x52964, x51637, x51639);
  nand n52965(x52965, x52964, x52963);
  nand n52967(x52967, x51642, x52966);
  nand n52968(x52968, x51641, x52965);
  nand n52969(x52969, x52968, x52967);
  nand n52971(x52971, x52963, x52967);
  nand n52972(x52972, x51644, x51646);
  nand n52973(x52973, x51643, x51645);
  nand n52974(x52974, x52973, x52972);
  nand n52976(x52976, x51648, x52975);
  nand n52977(x52977, x51647, x52974);
  nand n52978(x52978, x52977, x52976);
  nand n52980(x52980, x52972, x52976);
  nand n52981(x52981, x51650, x51652);
  nand n52982(x52982, x51649, x51651);
  nand n52983(x52983, x52982, x52981);
  nand n52985(x52985, x51654, x52984);
  nand n52986(x52986, x51653, x52983);
  nand n52987(x52987, x52986, x52985);
  nand n52989(x52989, x52981, x52985);
  nand n52990(x52990, x51656, x51658);
  nand n52991(x52991, x51655, x51657);
  nand n52992(x52992, x52991, x52990);
  nand n52994(x52994, x51660, x52993);
  nand n52995(x52995, x51659, x52992);
  nand n52996(x52996, x52995, x52994);
  nand n52998(x52998, x52990, x52994);
  nand n52999(x52999, x51662, x51664);
  nand n53000(x53000, x51661, x51663);
  nand n53001(x53001, x53000, x52999);
  nand n53003(x53003, x51666, x53002);
  nand n53004(x53004, x51665, x53001);
  nand n53005(x53005, x53004, x53003);
  nand n53007(x53007, x52999, x53003);
  nand n53008(x53008, x51668, x51670);
  nand n53009(x53009, x51667, x51669);
  nand n53010(x53010, x53009, x53008);
  nand n53012(x53012, x51672, x53011);
  nand n53013(x53013, x51671, x53010);
  nand n53014(x53014, x53013, x53012);
  nand n53016(x53016, x53008, x53012);
  nand n53017(x53017, x51674, x51676);
  nand n53018(x53018, x51673, x51675);
  nand n53019(x53019, x53018, x53017);
  nand n53021(x53021, x51678, x53020);
  nand n53022(x53022, x51677, x53019);
  nand n53023(x53023, x53022, x53021);
  nand n53025(x53025, x53017, x53021);
  nand n53026(x53026, x51680, x51682);
  nand n53027(x53027, x51679, x51681);
  nand n53028(x53028, x53027, x53026);
  nand n53030(x53030, x51684, x53029);
  nand n53031(x53031, x51683, x53028);
  nand n53032(x53032, x53031, x53030);
  nand n53034(x53034, x53026, x53030);
  nand n53035(x53035, x51686, x51688);
  nand n53036(x53036, x51685, x51687);
  nand n53037(x53037, x53036, x53035);
  nand n53039(x53039, x51690, x53038);
  nand n53040(x53040, x51689, x53037);
  nand n53041(x53041, x53040, x53039);
  nand n53042(x53042, x53035, x53039);
  nand n53043(x53043, x51692, x51694);
  nand n53044(x53044, x51691, x51693);
  nand n53045(x53045, x53044, x53043);
  nand n53047(x53047, x51696, x53046);
  nand n53048(x53048, x51695, x53045);
  nand n53049(x53049, x53048, x53047);
  nand n53051(x53051, x53043, x53047);
  nand n53052(x53052, x51698, x51700);
  nand n53053(x53053, x51697, x51699);
  nand n53054(x53054, x53053, x53052);
  nand n53056(x53056, x51702, x53055);
  nand n53057(x53057, x51701, x53054);
  nand n53058(x53058, x53057, x53056);
  nand n53060(x53060, x53052, x53056);
  nand n53061(x53061, x51704, x51706);
  nand n53062(x53062, x51703, x51705);
  nand n53063(x53063, x53062, x53061);
  nand n53065(x53065, x51708, x53064);
  nand n53066(x53066, x51707, x53063);
  nand n53067(x53067, x53066, x53065);
  nand n53069(x53069, x53061, x53065);
  nand n53070(x53070, x51710, x51712);
  nand n53071(x53071, x51709, x51711);
  nand n53072(x53072, x53071, x53070);
  nand n53074(x53074, x51714, x53073);
  nand n53075(x53075, x51713, x53072);
  nand n53076(x53076, x53075, x53074);
  nand n53078(x53078, x53070, x53074);
  nand n53079(x53079, x51716, x51718);
  nand n53080(x53080, x51715, x51717);
  nand n53081(x53081, x53080, x53079);
  nand n53083(x53083, x51720, x53082);
  nand n53084(x53084, x51719, x53081);
  nand n53085(x53085, x53084, x53083);
  nand n53087(x53087, x53079, x53083);
  nand n53088(x53088, x51722, x51724);
  nand n53089(x53089, x51721, x51723);
  nand n53090(x53090, x53089, x53088);
  nand n53092(x53092, x51726, x53091);
  nand n53093(x53093, x51725, x53090);
  nand n53094(x53094, x53093, x53092);
  nand n53096(x53096, x53088, x53092);
  nand n53097(x53097, x51728, x51730);
  nand n53098(x53098, x51727, x51729);
  nand n53099(x53099, x53098, x53097);
  nand n53101(x53101, x51732, x53100);
  nand n53102(x53102, x51731, x53099);
  nand n53103(x53103, x53102, x53101);
  nand n53105(x53105, x53097, x53101);
  nand n53106(x53106, x51734, x51736);
  nand n53107(x53107, x51733, x51735);
  nand n53108(x53108, x53107, x53106);
  nand n53110(x53110, x51738, x53109);
  nand n53111(x53111, x51737, x53108);
  nand n53112(x53112, x53111, x53110);
  nand n53114(x53114, x53106, x53110);
  nand n53115(x53115, x51741, x51743);
  nand n53116(x53116, x51740, x51742);
  nand n53117(x53117, x53116, x53115);
  nand n53119(x53119, x51745, x53118);
  nand n53120(x53120, x51744, x53117);
  nand n53121(x53121, x53120, x53119);
  nand n53122(x53122, x53115, x53119);
  nand n53123(x53123, x51747, x51749);
  nand n53124(x53124, x51746, x51748);
  nand n53125(x53125, x53124, x53123);
  nand n53127(x53127, x51751, x53126);
  nand n53128(x53128, x51750, x53125);
  nand n53129(x53129, x53128, x53127);
  nand n53131(x53131, x53123, x53127);
  nand n53132(x53132, x51753, x51755);
  nand n53133(x53133, x51752, x51754);
  nand n53134(x53134, x53133, x53132);
  nand n53136(x53136, x51757, x53135);
  nand n53137(x53137, x51756, x53134);
  nand n53138(x53138, x53137, x53136);
  nand n53140(x53140, x53132, x53136);
  nand n53141(x53141, x51759, x51761);
  nand n53142(x53142, x51758, x51760);
  nand n53143(x53143, x53142, x53141);
  nand n53145(x53145, x51763, x53144);
  nand n53146(x53146, x51762, x53143);
  nand n53147(x53147, x53146, x53145);
  nand n53149(x53149, x53141, x53145);
  nand n53150(x53150, x51765, x51767);
  nand n53151(x53151, x51764, x51766);
  nand n53152(x53152, x53151, x53150);
  nand n53154(x53154, x51769, x53153);
  nand n53155(x53155, x51768, x53152);
  nand n53156(x53156, x53155, x53154);
  nand n53158(x53158, x53150, x53154);
  nand n53159(x53159, x51771, x51773);
  nand n53160(x53160, x51770, x51772);
  nand n53161(x53161, x53160, x53159);
  nand n53163(x53163, x51775, x53162);
  nand n53164(x53164, x51774, x53161);
  nand n53165(x53165, x53164, x53163);
  nand n53167(x53167, x53159, x53163);
  nand n53168(x53168, x51777, x51779);
  nand n53169(x53169, x51776, x51778);
  nand n53170(x53170, x53169, x53168);
  nand n53172(x53172, x51781, x53171);
  nand n53173(x53173, x51780, x53170);
  nand n53174(x53174, x53173, x53172);
  nand n53176(x53176, x53168, x53172);
  nand n53177(x53177, x51783, x51785);
  nand n53178(x53178, x51782, x51784);
  nand n53179(x53179, x53178, x53177);
  nand n53181(x53181, x51787, x53180);
  nand n53182(x53182, x51786, x53179);
  nand n53183(x53183, x53182, x53181);
  nand n53185(x53185, x53177, x53181);
  nand n53186(x53186, x51789, x51791);
  nand n53187(x53187, x51788, x51790);
  nand n53188(x53188, x53187, x53186);
  nand n53190(x53190, x51793, x53189);
  nand n53191(x53191, x51792, x53188);
  nand n53192(x53192, x53191, x53190);
  nand n53194(x53194, x53186, x53190);
  nand n53195(x53195, x51795, x51797);
  nand n53196(x53196, x51794, x51796);
  nand n53197(x53197, x53196, x53195);
  nand n53198(x53198, x51799, x51801);
  nand n53199(x53199, x51798, x51800);
  nand n53200(x53200, x53199, x53198);
  nand n53202(x53202, x51803, x53201);
  nand n53203(x53203, x51802, x53200);
  nand n53204(x53204, x53203, x53202);
  nand n53206(x53206, x53198, x53202);
  nand n53207(x53207, x51805, x51807);
  nand n53208(x53208, x51804, x51806);
  nand n53209(x53209, x53208, x53207);
  nand n53211(x53211, x51809, x53210);
  nand n53212(x53212, x51808, x53209);
  nand n53213(x53213, x53212, x53211);
  nand n53215(x53215, x53207, x53211);
  nand n53216(x53216, x51811, x51813);
  nand n53217(x53217, x51810, x51812);
  nand n53218(x53218, x53217, x53216);
  nand n53220(x53220, x51815, x53219);
  nand n53221(x53221, x51814, x53218);
  nand n53222(x53222, x53221, x53220);
  nand n53224(x53224, x53216, x53220);
  nand n53225(x53225, x51817, x51819);
  nand n53226(x53226, x51816, x51818);
  nand n53227(x53227, x53226, x53225);
  nand n53229(x53229, x51821, x53228);
  nand n53230(x53230, x51820, x53227);
  nand n53231(x53231, x53230, x53229);
  nand n53233(x53233, x53225, x53229);
  nand n53234(x53234, x51823, x51825);
  nand n53235(x53235, x51822, x51824);
  nand n53236(x53236, x53235, x53234);
  nand n53238(x53238, x51827, x53237);
  nand n53239(x53239, x51826, x53236);
  nand n53240(x53240, x53239, x53238);
  nand n53242(x53242, x53234, x53238);
  nand n53243(x53243, x51829, x51831);
  nand n53244(x53244, x51828, x51830);
  nand n53245(x53245, x53244, x53243);
  nand n53247(x53247, x51833, x53246);
  nand n53248(x53248, x51832, x53245);
  nand n53249(x53249, x53248, x53247);
  nand n53251(x53251, x53243, x53247);
  nand n53252(x53252, x51835, x51837);
  nand n53253(x53253, x51834, x51836);
  nand n53254(x53254, x53253, x53252);
  nand n53256(x53256, x51839, x53255);
  nand n53257(x53257, x51838, x53254);
  nand n53258(x53258, x53257, x53256);
  nand n53260(x53260, x53252, x53256);
  nand n53261(x53261, x51841, x51843);
  nand n53262(x53262, x51840, x51842);
  nand n53263(x53263, x53262, x53261);
  nand n53265(x53265, x51845, x53264);
  nand n53266(x53266, x51844, x53263);
  nand n53267(x53267, x53266, x53265);
  nand n53269(x53269, x53261, x53265);
  nand n53270(x53270, x51847, x51849);
  nand n53271(x53271, x51846, x51848);
  nand n53272(x53272, x53271, x53270);
  nand n53274(x53274, x51851, x53273);
  nand n53275(x53275, x51850, x53272);
  nand n53276(x53276, x53275, x53274);
  nand n53278(x53278, x53270, x53274);
  nand n53279(x53279, x51853, x51855);
  nand n53280(x53280, x51852, x51854);
  nand n53281(x53281, x53280, x53279);
  nand n53283(x53283, x51857, x53282);
  nand n53284(x53284, x51856, x53281);
  nand n53285(x53285, x53284, x53283);
  nand n53287(x53287, x53279, x53283);
  nand n53288(x53288, x51859, x51861);
  nand n53289(x53289, x51858, x51860);
  nand n53290(x53290, x53289, x53288);
  nand n53292(x53292, x51863, x53291);
  nand n53293(x53293, x51862, x53290);
  nand n53294(x53294, x53293, x53292);
  nand n53296(x53296, x53288, x53292);
  nand n53297(x53297, x51865, x51867);
  nand n53298(x53298, x51864, x51866);
  nand n53299(x53299, x53298, x53297);
  nand n53301(x53301, x51869, x53300);
  nand n53302(x53302, x51868, x53299);
  nand n53303(x53303, x53302, x53301);
  nand n53305(x53305, x53297, x53301);
  nand n53306(x53306, x51871, x51873);
  nand n53307(x53307, x51870, x51872);
  nand n53308(x53308, x53307, x53306);
  nand n53310(x53310, x51875, x53309);
  nand n53311(x53311, x51874, x53308);
  nand n53312(x53312, x53311, x53310);
  nand n53314(x53314, x53306, x53310);
  nand n53315(x53315, x51877, x51879);
  nand n53316(x53316, x51876, x51878);
  nand n53317(x53317, x53316, x53315);
  nand n53319(x53319, x51881, x53318);
  nand n53320(x53320, x51880, x53317);
  nand n53321(x53321, x53320, x53319);
  nand n53323(x53323, x53315, x53319);
  nand n53324(x53324, x51883, x51885);
  nand n53325(x53325, x51882, x51884);
  nand n53326(x53326, x53325, x53324);
  nand n53328(x53328, x51887, x53327);
  nand n53329(x53329, x51886, x53326);
  nand n53330(x53330, x53329, x53328);
  nand n53332(x53332, x53324, x53328);
  nand n53333(x53333, x51889, x51891);
  nand n53334(x53334, x51888, x51890);
  nand n53335(x53335, x53334, x53333);
  nand n53337(x53337, x51893, x53336);
  nand n53338(x53338, x51892, x53335);
  nand n53339(x53339, x53338, x53337);
  nand n53341(x53341, x53333, x53337);
  nand n53342(x53342, x51895, x51897);
  nand n53343(x53343, x51894, x51896);
  nand n53344(x53344, x53343, x53342);
  nand n53346(x53346, x51899, x53345);
  nand n53347(x53347, x51898, x53344);
  nand n53348(x53348, x53347, x53346);
  nand n53350(x53350, x53342, x53346);
  nand n53351(x53351, x51901, x51903);
  nand n53352(x53352, x51900, x51902);
  nand n53353(x53353, x53352, x53351);
  nand n53355(x53355, x51905, x53354);
  nand n53356(x53356, x51904, x53353);
  nand n53357(x53357, x53356, x53355);
  nand n53359(x53359, x53351, x53355);
  nand n53360(x53360, x51907, x51909);
  nand n53361(x53361, x51906, x51908);
  nand n53362(x53362, x53361, x53360);
  nand n53364(x53364, x51911, x53363);
  nand n53365(x53365, x51910, x53362);
  nand n53366(x53366, x53365, x53364);
  nand n53368(x53368, x53360, x53364);
  nand n53369(x53369, x51913, x51915);
  nand n53370(x53370, x51912, x51914);
  nand n53371(x53371, x53370, x53369);
  nand n53373(x53373, x51917, x53372);
  nand n53374(x53374, x51916, x53371);
  nand n53375(x53375, x53374, x53373);
  nand n53377(x53377, x53369, x53373);
  nand n53378(x53378, x51920, x51922);
  nand n53379(x53379, x51919, x51921);
  nand n53380(x53380, x53379, x53378);
  nand n53382(x53382, x51924, x53381);
  nand n53383(x53383, x51923, x53380);
  nand n53384(x53384, x53383, x53382);
  nand n53386(x53386, x51926, x51928);
  nand n53387(x53387, x51925, x51927);
  nand n53388(x53388, x53387, x53386);
  nand n53390(x53390, x51930, x53389);
  nand n53391(x53391, x51929, x53388);
  nand n53392(x53392, x53391, x53390);
  nand n53394(x53394, x51932, x51934);
  nand n53395(x53395, x51931, x51933);
  nand n53396(x53396, x53395, x53394);
  nand n53398(x53398, x51936, x53397);
  nand n53399(x53399, x51935, x53396);
  nand n53400(x53400, x53399, x53398);
  nand n53402(x53402, x51938, x51940);
  nand n53403(x53403, x51937, x51939);
  nand n53404(x53404, x53403, x53402);
  nand n53406(x53406, x51942, x53405);
  nand n53407(x53407, x51941, x53404);
  nand n53408(x53408, x53407, x53406);
  nand n53410(x53410, x51944, x51946);
  nand n53411(x53411, x51943, x51945);
  nand n53412(x53412, x53411, x53410);
  nand n53414(x53414, x51948, x53413);
  nand n53415(x53415, x51947, x53412);
  nand n53416(x53416, x53415, x53414);
  nand n53418(x53418, x51950, x51952);
  nand n53419(x53419, x51949, x51951);
  nand n53420(x53420, x53419, x53418);
  nand n53422(x53422, x51954, x53421);
  nand n53423(x53423, x51953, x53420);
  nand n53424(x53424, x53423, x53422);
  nand n53426(x53426, x51956, x51958);
  nand n53427(x53427, x51955, x51957);
  nand n53428(x53428, x53427, x53426);
  nand n53430(x53430, x51960, x53429);
  nand n53431(x53431, x51959, x53428);
  nand n53432(x53432, x53431, x53430);
  nand n53434(x53434, x51962, x51964);
  nand n53435(x53435, x51961, x51963);
  nand n53436(x53436, x53435, x53434);
  nand n53438(x53438, x51966, x53437);
  nand n53439(x53439, x51965, x53436);
  nand n53440(x53440, x53439, x53438);
  nand n53442(x53442, x51968, x51970);
  nand n53443(x53443, x51967, x51969);
  nand n53444(x53444, x53443, x53442);
  nand n53446(x53446, x51972, x53445);
  nand n53447(x53447, x51971, x53444);
  nand n53448(x53448, x53447, x53446);
  nand n53450(x53450, x51974, x51976);
  nand n53451(x53451, x51973, x51975);
  nand n53452(x53452, x53451, x53450);
  nand n53454(x53454, x51978, x53453);
  nand n53455(x53455, x51977, x53452);
  nand n53456(x53456, x53455, x53454);
  nand n53458(x53458, x51980, x51982);
  nand n53459(x53459, x51979, x51981);
  nand n53460(x53460, x53459, x53458);
  nand n53464(x53464, x52009, x85589);
  nand n53466(x53466, x53465, x52010);
  nand n53467(x53467, x53466, x53464);
  nand n53468(x53468, x52020, x52028);
  nand n53471(x53471, x53470, x53469);
  nand n53472(x53472, x53471, x53468);
  nand n53473(x53473, x52044, x85590);
  nand n53474(x53474, x52043, x50990);
  nand n53475(x53475, x53474, x53473);
  nand n53476(x53476, x52036, x52045);
  nand n53479(x53479, x53478, x53477);
  nand n53480(x53480, x53479, x53476);
  nand n53481(x53481, x52061, x85591);
  nand n53482(x53482, x52060, x52065);
  nand n53483(x53483, x53482, x53481);
  nand n53484(x53484, x52053, x52062);
  nand n53487(x53487, x53486, x53485);
  nand n53488(x53488, x53487, x53484);
  nand n53490(x53490, x85592, x53489);
  nand n53491(x53491, x52063, x53488);
  nand n53492(x53492, x53491, x53490);
  nand n53493(x53493, x53484, x53490);
  nand n53494(x53494, x52081, x52090);
  nand n53495(x53495, x52080, x52089);
  nand n53496(x53496, x53495, x53494);
  nand n53497(x53497, x52073, x52082);
  nand n53500(x53500, x53499, x53498);
  nand n53501(x53501, x53500, x53497);
  nand n53503(x53503, x52091, x53502);
  nand n53505(x53505, x53504, x53501);
  nand n53506(x53506, x53505, x53503);
  nand n53507(x53507, x53497, x53503);
  nand n53508(x53508, x52107, x52116);
  nand n53509(x53509, x52106, x52115);
  nand n53510(x53510, x53509, x53508);
  nand n53512(x53512, x85593, x53511);
  nand n53513(x53513, x51043, x53510);
  nand n53514(x53514, x53513, x53512);
  nand n53516(x53516, x53508, x53512);
  nand n53517(x53517, x52099, x52108);
  nand n53520(x53520, x53519, x53518);
  nand n53521(x53521, x53520, x53517);
  nand n53523(x53523, x52117, x53522);
  nand n53525(x53525, x53524, x53521);
  nand n53526(x53526, x53525, x53523);
  nand n53527(x53527, x53517, x53523);
  nand n53528(x53528, x52133, x52142);
  nand n53529(x53529, x52132, x52141);
  nand n53530(x53530, x53529, x53528);
  nand n53532(x53532, x85594, x53531);
  nand n53533(x53533, x52146, x53530);
  nand n53534(x53534, x53533, x53532);
  nand n53536(x53536, x53528, x53532);
  nand n53537(x53537, x52125, x52134);
  nand n53540(x53540, x53539, x53538);
  nand n53541(x53541, x53540, x53537);
  nand n53543(x53543, x52143, x53542);
  nand n53545(x53545, x53544, x53541);
  nand n53546(x53546, x53545, x53543);
  nand n53547(x53547, x53537, x53543);
  nand n53548(x53548, x52162, x52171);
  nand n53549(x53549, x52161, x52170);
  nand n53550(x53550, x53549, x53548);
  nand n53552(x53552, x52180, x53551);
  nand n53553(x53553, x52179, x53550);
  nand n53554(x53554, x53553, x53552);
  nand n53556(x53556, x53548, x53552);
  nand n53557(x53557, x52154, x52163);
  nand n53560(x53560, x53559, x53558);
  nand n53561(x53561, x53560, x53557);
  nand n53563(x53563, x52172, x53562);
  nand n53565(x53565, x53564, x53561);
  nand n53566(x53566, x53565, x53563);
  nand n53567(x53567, x53557, x53563);
  nand n53569(x53569, x52197, x52206);
  nand n53570(x53570, x52196, x52205);
  nand n53571(x53571, x53570, x53569);
  nand n53573(x53573, x52215, x53572);
  nand n53574(x53574, x52214, x53571);
  nand n53575(x53575, x53574, x53573);
  nand n53577(x53577, x53569, x53573);
  nand n53578(x53578, x52189, x52198);
  nand n53581(x53581, x53580, x53579);
  nand n53582(x53582, x53581, x53578);
  nand n53584(x53584, x52207, x53583);
  nand n53586(x53586, x53585, x53582);
  nand n53587(x53587, x53586, x53584);
  nand n53588(x53588, x53578, x53584);
  nand n53590(x53590, x52232, x52241);
  nand n53591(x53591, x52231, x52240);
  nand n53592(x53592, x53591, x53590);
  nand n53594(x53594, x52250, x53593);
  nand n53595(x53595, x52249, x53592);
  nand n53596(x53596, x53595, x53594);
  nand n53598(x53598, x53590, x53594);
  nand n53599(x53599, x52224, x52233);
  nand n53602(x53602, x53601, x53600);
  nand n53603(x53603, x53602, x53599);
  nand n53605(x53605, x52242, x53604);
  nand n53607(x53607, x53606, x53603);
  nand n53608(x53608, x53607, x53605);
  nand n53609(x53609, x53599, x53605);
  nand n53610(x53610, x52251, x85595);
  nand n53612(x53612, x53611, x52252);
  nand n53613(x53613, x53612, x53610);
  nand n53614(x53614, x52270, x52279);
  nand n53615(x53615, x52269, x52278);
  nand n53616(x53616, x53615, x53614);
  nand n53618(x53618, x52288, x53617);
  nand n53619(x53619, x52287, x53616);
  nand n53620(x53620, x53619, x53618);
  nand n53622(x53622, x53614, x53618);
  nand n53623(x53623, x52262, x52271);
  nand n53626(x53626, x53625, x53624);
  nand n53627(x53627, x53626, x53623);
  nand n53629(x53629, x52280, x53628);
  nand n53631(x53631, x53630, x53627);
  nand n53632(x53632, x53631, x53629);
  nand n53633(x53633, x53623, x53629);
  nand n53634(x53634, x52289, x52297);
  nand n53637(x53637, x53636, x53635);
  nand n53638(x53638, x53637, x53634);
  nand n53639(x53639, x52313, x52322);
  nand n53640(x53640, x52312, x52321);
  nand n53641(x53641, x53640, x53639);
  nand n53643(x53643, x52331, x53642);
  nand n53644(x53644, x52330, x53641);
  nand n53645(x53645, x53644, x53643);
  nand n53647(x53647, x53639, x53643);
  nand n53648(x53648, x52340, x85596);
  nand n53649(x53649, x52339, x51203);
  nand n53650(x53650, x53649, x53648);
  nand n53651(x53651, x52305, x52314);
  nand n53654(x53654, x53653, x53652);
  nand n53655(x53655, x53654, x53651);
  nand n53657(x53657, x52323, x53656);
  nand n53659(x53659, x53658, x53655);
  nand n53660(x53660, x53659, x53657);
  nand n53661(x53661, x53651, x53657);
  nand n53662(x53662, x52332, x52341);
  nand n53665(x53665, x53664, x53663);
  nand n53666(x53666, x53665, x53662);
  nand n53667(x53667, x52357, x52366);
  nand n53668(x53668, x52356, x52365);
  nand n53669(x53669, x53668, x53667);
  nand n53671(x53671, x52375, x53670);
  nand n53672(x53672, x52374, x53669);
  nand n53673(x53673, x53672, x53671);
  nand n53675(x53675, x53667, x53671);
  nand n53676(x53676, x52384, x85597);
  nand n53677(x53677, x52383, x52388);
  nand n53678(x53678, x53677, x53676);
  nand n53679(x53679, x52349, x52358);
  nand n53682(x53682, x53681, x53680);
  nand n53683(x53683, x53682, x53679);
  nand n53685(x53685, x52367, x53684);
  nand n53687(x53687, x53686, x53683);
  nand n53688(x53688, x53687, x53685);
  nand n53689(x53689, x53679, x53685);
  nand n53690(x53690, x52376, x52385);
  nand n53693(x53693, x53692, x53691);
  nand n53694(x53694, x53693, x53690);
  nand n53696(x53696, x85598, x53695);
  nand n53697(x53697, x52386, x53694);
  nand n53698(x53698, x53697, x53696);
  nand n53700(x53700, x53690, x53696);
  nand n53701(x53701, x52404, x52413);
  nand n53702(x53702, x52403, x52412);
  nand n53703(x53703, x53702, x53701);
  nand n53705(x53705, x52422, x53704);
  nand n53706(x53706, x52421, x53703);
  nand n53707(x53707, x53706, x53705);
  nand n53709(x53709, x53701, x53705);
  nand n53710(x53710, x52431, x52440);
  nand n53711(x53711, x52430, x52439);
  nand n53712(x53712, x53711, x53710);
  nand n53713(x53713, x52396, x52405);
  nand n53716(x53716, x53715, x53714);
  nand n53717(x53717, x53716, x53713);
  nand n53719(x53719, x52414, x53718);
  nand n53721(x53721, x53720, x53717);
  nand n53722(x53722, x53721, x53719);
  nand n53723(x53723, x53713, x53719);
  nand n53724(x53724, x52423, x52432);
  nand n53727(x53727, x53726, x53725);
  nand n53728(x53728, x53727, x53724);
  nand n53730(x53730, x52441, x53729);
  nand n53732(x53732, x53731, x53728);
  nand n53733(x53733, x53732, x53730);
  nand n53735(x53735, x53724, x53730);
  nand n53736(x53736, x52457, x52466);
  nand n53737(x53737, x52456, x52465);
  nand n53738(x53738, x53737, x53736);
  nand n53740(x53740, x52475, x53739);
  nand n53741(x53741, x52474, x53738);
  nand n53742(x53742, x53741, x53740);
  nand n53744(x53744, x53736, x53740);
  nand n53745(x53745, x52484, x52493);
  nand n53746(x53746, x52483, x52492);
  nand n53747(x53747, x53746, x53745);
  nand n53749(x53749, x85599, x53748);
  nand n53750(x53750, x51310, x53747);
  nand n53751(x53751, x53750, x53749);
  nand n53752(x53752, x53745, x53749);
  nand n53753(x53753, x52449, x52458);
  nand n53756(x53756, x53755, x53754);
  nand n53757(x53757, x53756, x53753);
  nand n53759(x53759, x52467, x53758);
  nand n53761(x53761, x53760, x53757);
  nand n53762(x53762, x53761, x53759);
  nand n53763(x53763, x53753, x53759);
  nand n53764(x53764, x52476, x52485);
  nand n53767(x53767, x53766, x53765);
  nand n53768(x53768, x53767, x53764);
  nand n53770(x53770, x52494, x53769);
  nand n53772(x53772, x53771, x53768);
  nand n53773(x53773, x53772, x53770);
  nand n53775(x53775, x53764, x53770);
  nand n53776(x53776, x52510, x52519);
  nand n53777(x53777, x52509, x52518);
  nand n53778(x53778, x53777, x53776);
  nand n53780(x53780, x52528, x53779);
  nand n53781(x53781, x52527, x53778);
  nand n53782(x53782, x53781, x53780);
  nand n53784(x53784, x53776, x53780);
  nand n53785(x53785, x52537, x52546);
  nand n53786(x53786, x52536, x52545);
  nand n53787(x53787, x53786, x53785);
  nand n53789(x53789, x85600, x53788);
  nand n53790(x53790, x52550, x53787);
  nand n53791(x53791, x53790, x53789);
  nand n53792(x53792, x53785, x53789);
  nand n53793(x53793, x52502, x52511);
  nand n53796(x53796, x53795, x53794);
  nand n53797(x53797, x53796, x53793);
  nand n53799(x53799, x52520, x53798);
  nand n53801(x53801, x53800, x53797);
  nand n53802(x53802, x53801, x53799);
  nand n53803(x53803, x53793, x53799);
  nand n53804(x53804, x52529, x52538);
  nand n53807(x53807, x53806, x53805);
  nand n53808(x53808, x53807, x53804);
  nand n53810(x53810, x52547, x53809);
  nand n53812(x53812, x53811, x53808);
  nand n53813(x53813, x53812, x53810);
  nand n53815(x53815, x53804, x53810);
  nand n53816(x53816, x52566, x52575);
  nand n53817(x53817, x52565, x52574);
  nand n53818(x53818, x53817, x53816);
  nand n53820(x53820, x52584, x53819);
  nand n53821(x53821, x52583, x53818);
  nand n53822(x53822, x53821, x53820);
  nand n53824(x53824, x53816, x53820);
  nand n53825(x53825, x52593, x52602);
  nand n53826(x53826, x52592, x52601);
  nand n53827(x53827, x53826, x53825);
  nand n53829(x53829, x52611, x53828);
  nand n53830(x53830, x52610, x53827);
  nand n53831(x53831, x53830, x53829);
  nand n53832(x53832, x53825, x53829);
  nand n53833(x53833, x52558, x52567);
  nand n53836(x53836, x53835, x53834);
  nand n53837(x53837, x53836, x53833);
  nand n53839(x53839, x52576, x53838);
  nand n53841(x53841, x53840, x53837);
  nand n53842(x53842, x53841, x53839);
  nand n53843(x53843, x53833, x53839);
  nand n53844(x53844, x52585, x52594);
  nand n53847(x53847, x53846, x53845);
  nand n53848(x53848, x53847, x53844);
  nand n53850(x53850, x52603, x53849);
  nand n53852(x53852, x53851, x53848);
  nand n53853(x53853, x53852, x53850);
  nand n53855(x53855, x53844, x53850);
  nand n53857(x53857, x52628, x52637);
  nand n53858(x53858, x52627, x52636);
  nand n53859(x53859, x53858, x53857);
  nand n53861(x53861, x52646, x53860);
  nand n53862(x53862, x52645, x53859);
  nand n53863(x53863, x53862, x53861);
  nand n53865(x53865, x53857, x53861);
  nand n53866(x53866, x52655, x52664);
  nand n53867(x53867, x52654, x52663);
  nand n53868(x53868, x53867, x53866);
  nand n53870(x53870, x52673, x53869);
  nand n53871(x53871, x52672, x53868);
  nand n53872(x53872, x53871, x53870);
  nand n53874(x53874, x53866, x53870);
  nand n53875(x53875, x52620, x52629);
  nand n53878(x53878, x53877, x53876);
  nand n53879(x53879, x53878, x53875);
  nand n53881(x53881, x52638, x53880);
  nand n53883(x53883, x53882, x53879);
  nand n53884(x53884, x53883, x53881);
  nand n53885(x53885, x53875, x53881);
  nand n53886(x53886, x52647, x52656);
  nand n53889(x53889, x53888, x53887);
  nand n53890(x53890, x53889, x53886);
  nand n53892(x53892, x52665, x53891);
  nand n53894(x53894, x53893, x53890);
  nand n53895(x53895, x53894, x53892);
  nand n53897(x53897, x53886, x53892);
  nand n53899(x53899, x52690, x52699);
  nand n53900(x53900, x52689, x52698);
  nand n53901(x53901, x53900, x53899);
  nand n53903(x53903, x52708, x53902);
  nand n53904(x53904, x52707, x53901);
  nand n53905(x53905, x53904, x53903);
  nand n53907(x53907, x53899, x53903);
  nand n53908(x53908, x52717, x52726);
  nand n53909(x53909, x52716, x52725);
  nand n53910(x53910, x53909, x53908);
  nand n53912(x53912, x52735, x53911);
  nand n53913(x53913, x52734, x53910);
  nand n53914(x53914, x53913, x53912);
  nand n53916(x53916, x53908, x53912);
  nand n53917(x53917, x52682, x52691);
  nand n53920(x53920, x53919, x53918);
  nand n53921(x53921, x53920, x53917);
  nand n53923(x53923, x52700, x53922);
  nand n53925(x53925, x53924, x53921);
  nand n53926(x53926, x53925, x53923);
  nand n53927(x53927, x53917, x53923);
  nand n53928(x53928, x52709, x52718);
  nand n53931(x53931, x53930, x53929);
  nand n53932(x53932, x53931, x53928);
  nand n53934(x53934, x52727, x53933);
  nand n53936(x53936, x53935, x53932);
  nand n53937(x53937, x53936, x53934);
  nand n53939(x53939, x53928, x53934);
  nand n53940(x53940, x52736, x85601);
  nand n53942(x53942, x53941, x52737);
  nand n53943(x53943, x53942, x53940);
  nand n53944(x53944, x52755, x52764);
  nand n53945(x53945, x52754, x52763);
  nand n53946(x53946, x53945, x53944);
  nand n53948(x53948, x52773, x53947);
  nand n53949(x53949, x52772, x53946);
  nand n53950(x53950, x53949, x53948);
  nand n53952(x53952, x53944, x53948);
  nand n53953(x53953, x52782, x52791);
  nand n53954(x53954, x52781, x52790);
  nand n53955(x53955, x53954, x53953);
  nand n53957(x53957, x52800, x53956);
  nand n53958(x53958, x52799, x53955);
  nand n53959(x53959, x53958, x53957);
  nand n53961(x53961, x53953, x53957);
  nand n53962(x53962, x52747, x52756);
  nand n53965(x53965, x53964, x53963);
  nand n53966(x53966, x53965, x53962);
  nand n53968(x53968, x52765, x53967);
  nand n53970(x53970, x53969, x53966);
  nand n53971(x53971, x53970, x53968);
  nand n53972(x53972, x53962, x53968);
  nand n53973(x53973, x52774, x52783);
  nand n53976(x53976, x53975, x53974);
  nand n53977(x53977, x53976, x53973);
  nand n53979(x53979, x52792, x53978);
  nand n53981(x53981, x53980, x53977);
  nand n53982(x53982, x53981, x53979);
  nand n53984(x53984, x53973, x53979);
  nand n53985(x53985, x52801, x52809);
  nand n53988(x53988, x53987, x53986);
  nand n53989(x53989, x53988, x53985);
  nand n53990(x53990, x52825, x52834);
  nand n53991(x53991, x52824, x52833);
  nand n53992(x53992, x53991, x53990);
  nand n53994(x53994, x52843, x53993);
  nand n53995(x53995, x52842, x53992);
  nand n53996(x53996, x53995, x53994);
  nand n53998(x53998, x53990, x53994);
  nand n53999(x53999, x52852, x52861);
  nand n54000(x54000, x52851, x52860);
  nand n54001(x54001, x54000, x53999);
  nand n54003(x54003, x52870, x54002);
  nand n54004(x54004, x52869, x54001);
  nand n54005(x54005, x54004, x54003);
  nand n54007(x54007, x53999, x54003);
  nand n54008(x54008, x52879, x85602);
  nand n54009(x54009, x52878, x51578);
  nand n54010(x54010, x54009, x54008);
  nand n54011(x54011, x52817, x52826);
  nand n54014(x54014, x54013, x54012);
  nand n54015(x54015, x54014, x54011);
  nand n54017(x54017, x52835, x54016);
  nand n54019(x54019, x54018, x54015);
  nand n54020(x54020, x54019, x54017);
  nand n54022(x54022, x54011, x54017);
  nand n54023(x54023, x52844, x52853);
  nand n54026(x54026, x54025, x54024);
  nand n54027(x54027, x54026, x54023);
  nand n54029(x54029, x52862, x54028);
  nand n54031(x54031, x54030, x54027);
  nand n54032(x54032, x54031, x54029);
  nand n54034(x54034, x54023, x54029);
  nand n54035(x54035, x52871, x52880);
  nand n54038(x54038, x54037, x54036);
  nand n54039(x54039, x54038, x54035);
  nand n54040(x54040, x52896, x52905);
  nand n54041(x54041, x52895, x52904);
  nand n54042(x54042, x54041, x54040);
  nand n54044(x54044, x52914, x54043);
  nand n54045(x54045, x52913, x54042);
  nand n54046(x54046, x54045, x54044);
  nand n54048(x54048, x54040, x54044);
  nand n54049(x54049, x52923, x52932);
  nand n54050(x54050, x52922, x52931);
  nand n54051(x54051, x54050, x54049);
  nand n54053(x54053, x52941, x54052);
  nand n54054(x54054, x52940, x54051);
  nand n54055(x54055, x54054, x54053);
  nand n54057(x54057, x54049, x54053);
  nand n54058(x54058, x52950, x85603);
  nand n54059(x54059, x52949, x52954);
  nand n54060(x54060, x54059, x54058);
  nand n54061(x54061, x52888, x52897);
  nand n54064(x54064, x54063, x54062);
  nand n54065(x54065, x54064, x54061);
  nand n54067(x54067, x52906, x54066);
  nand n54069(x54069, x54068, x54065);
  nand n54070(x54070, x54069, x54067);
  nand n54072(x54072, x54061, x54067);
  nand n54073(x54073, x52915, x52924);
  nand n54076(x54076, x54075, x54074);
  nand n54077(x54077, x54076, x54073);
  nand n54079(x54079, x52933, x54078);
  nand n54081(x54081, x54080, x54077);
  nand n54082(x54082, x54081, x54079);
  nand n54084(x54084, x54073, x54079);
  nand n54085(x54085, x52942, x52951);
  nand n54088(x54088, x54087, x54086);
  nand n54089(x54089, x54088, x54085);
  nand n54091(x54091, x85604, x54090);
  nand n54092(x54092, x52952, x54089);
  nand n54093(x54093, x54092, x54091);
  nand n54095(x54095, x54085, x54091);
  nand n54096(x54096, x52970, x52979);
  nand n54097(x54097, x52969, x52978);
  nand n54098(x54098, x54097, x54096);
  nand n54100(x54100, x52988, x54099);
  nand n54101(x54101, x52987, x54098);
  nand n54102(x54102, x54101, x54100);
  nand n54104(x54104, x54096, x54100);
  nand n54105(x54105, x52997, x53006);
  nand n54106(x54106, x52996, x53005);
  nand n54107(x54107, x54106, x54105);
  nand n54109(x54109, x53015, x54108);
  nand n54110(x54110, x53014, x54107);
  nand n54111(x54111, x54110, x54109);
  nand n54113(x54113, x54105, x54109);
  nand n54114(x54114, x53024, x53033);
  nand n54115(x54115, x53023, x53032);
  nand n54116(x54116, x54115, x54114);
  nand n54117(x54117, x52962, x52971);
  nand n54120(x54120, x54119, x54118);
  nand n54121(x54121, x54120, x54117);
  nand n54123(x54123, x52980, x54122);
  nand n54125(x54125, x54124, x54121);
  nand n54126(x54126, x54125, x54123);
  nand n54128(x54128, x54117, x54123);
  nand n54129(x54129, x52989, x52998);
  nand n54132(x54132, x54131, x54130);
  nand n54133(x54133, x54132, x54129);
  nand n54135(x54135, x53007, x54134);
  nand n54137(x54137, x54136, x54133);
  nand n54138(x54138, x54137, x54135);
  nand n54140(x54140, x54129, x54135);
  nand n54141(x54141, x53016, x53025);
  nand n54144(x54144, x54143, x54142);
  nand n54145(x54145, x54144, x54141);
  nand n54147(x54147, x53034, x54146);
  nand n54149(x54149, x54148, x54145);
  nand n54150(x54150, x54149, x54147);
  nand n54152(x54152, x54141, x54147);
  nand n54153(x54153, x53050, x53059);
  nand n54154(x54154, x53049, x53058);
  nand n54155(x54155, x54154, x54153);
  nand n54157(x54157, x53068, x54156);
  nand n54158(x54158, x53067, x54155);
  nand n54159(x54159, x54158, x54157);
  nand n54161(x54161, x54153, x54157);
  nand n54162(x54162, x53077, x53086);
  nand n54163(x54163, x53076, x53085);
  nand n54164(x54164, x54163, x54162);
  nand n54166(x54166, x53095, x54165);
  nand n54167(x54167, x53094, x54164);
  nand n54168(x54168, x54167, x54166);
  nand n54170(x54170, x54162, x54166);
  nand n54171(x54171, x53104, x53113);
  nand n54172(x54172, x53103, x53112);
  nand n54173(x54173, x54172, x54171);
  nand n54175(x54175, x85605, x54174);
  nand n54176(x54176, x51739, x54173);
  nand n54177(x54177, x54176, x54175);
  nand n54179(x54179, x54171, x54175);
  nand n54180(x54180, x53042, x53051);
  nand n54183(x54183, x54182, x54181);
  nand n54184(x54184, x54183, x54180);
  nand n54186(x54186, x53060, x54185);
  nand n54188(x54188, x54187, x54184);
  nand n54189(x54189, x54188, x54186);
  nand n54191(x54191, x54180, x54186);
  nand n54192(x54192, x53069, x53078);
  nand n54195(x54195, x54194, x54193);
  nand n54196(x54196, x54195, x54192);
  nand n54198(x54198, x53087, x54197);
  nand n54200(x54200, x54199, x54196);
  nand n54201(x54201, x54200, x54198);
  nand n54203(x54203, x54192, x54198);
  nand n54204(x54204, x53096, x53105);
  nand n54207(x54207, x54206, x54205);
  nand n54208(x54208, x54207, x54204);
  nand n54210(x54210, x53114, x54209);
  nand n54212(x54212, x54211, x54208);
  nand n54213(x54213, x54212, x54210);
  nand n54215(x54215, x54204, x54210);
  nand n54216(x54216, x53130, x53139);
  nand n54217(x54217, x53129, x53138);
  nand n54218(x54218, x54217, x54216);
  nand n54220(x54220, x53148, x54219);
  nand n54221(x54221, x53147, x54218);
  nand n54222(x54222, x54221, x54220);
  nand n54224(x54224, x54216, x54220);
  nand n54225(x54225, x53157, x53166);
  nand n54226(x54226, x53156, x53165);
  nand n54227(x54227, x54226, x54225);
  nand n54229(x54229, x53175, x54228);
  nand n54230(x54230, x53174, x54227);
  nand n54231(x54231, x54230, x54229);
  nand n54233(x54233, x54225, x54229);
  nand n54234(x54234, x53184, x53193);
  nand n54235(x54235, x53183, x53192);
  nand n54236(x54236, x54235, x54234);
  nand n54238(x54238, x85606, x54237);
  nand n54239(x54239, x53197, x54236);
  nand n54240(x54240, x54239, x54238);
  nand n54242(x54242, x54234, x54238);
  nand n54243(x54243, x53122, x53131);
  nand n54246(x54246, x54245, x54244);
  nand n54247(x54247, x54246, x54243);
  nand n54249(x54249, x53140, x54248);
  nand n54251(x54251, x54250, x54247);
  nand n54252(x54252, x54251, x54249);
  nand n54254(x54254, x54243, x54249);
  nand n54255(x54255, x53149, x53158);
  nand n54258(x54258, x54257, x54256);
  nand n54259(x54259, x54258, x54255);
  nand n54261(x54261, x53167, x54260);
  nand n54263(x54263, x54262, x54259);
  nand n54264(x54264, x54263, x54261);
  nand n54266(x54266, x54255, x54261);
  nand n54267(x54267, x53176, x53185);
  nand n54270(x54270, x54269, x54268);
  nand n54271(x54271, x54270, x54267);
  nand n54273(x54273, x53194, x54272);
  nand n54275(x54275, x54274, x54271);
  nand n54276(x54276, x54275, x54273);
  nand n54278(x54278, x54267, x54273);
  nand n54279(x54279, x53205, x85649);
  nand n54280(x54280, x53204, x53195);
  nand n54281(x54281, x54280, x54279);
  nand n54283(x54283, x53214, x53223);
  nand n54284(x54284, x53213, x53222);
  nand n54285(x54285, x54284, x54283);
  nand n54287(x54287, x53232, x54286);
  nand n54288(x54288, x53231, x54285);
  nand n54289(x54289, x54288, x54287);
  nand n54291(x54291, x54283, x54287);
  nand n54292(x54292, x53241, x53250);
  nand n54293(x54293, x53240, x53249);
  nand n54294(x54294, x54293, x54292);
  nand n54296(x54296, x53259, x54295);
  nand n54297(x54297, x53258, x54294);
  nand n54298(x54298, x54297, x54296);
  nand n54300(x54300, x54292, x54296);
  nand n54301(x54301, x53268, x53277);
  nand n54302(x54302, x53267, x53276);
  nand n54303(x54303, x54302, x54301);
  nand n54305(x54305, x53286, x54304);
  nand n54306(x54306, x53285, x54303);
  nand n54307(x54307, x54306, x54305);
  nand n54309(x54309, x54301, x54305);
  nand n54310(x54310, x53206, x53215);
  nand n54313(x54313, x54312, x54311);
  nand n54314(x54314, x54313, x54310);
  nand n54316(x54316, x53224, x54315);
  nand n54318(x54318, x54317, x54314);
  nand n54319(x54319, x54318, x54316);
  nand n54321(x54321, x54310, x54316);
  nand n54322(x54322, x53233, x53242);
  nand n54325(x54325, x54324, x54323);
  nand n54326(x54326, x54325, x54322);
  nand n54328(x54328, x53251, x54327);
  nand n54330(x54330, x54329, x54326);
  nand n54331(x54331, x54330, x54328);
  nand n54333(x54333, x54322, x54328);
  nand n54334(x54334, x53260, x53269);
  nand n54337(x54337, x54336, x54335);
  nand n54338(x54338, x54337, x54334);
  nand n54340(x54340, x53278, x54339);
  nand n54342(x54342, x54341, x54338);
  nand n54343(x54343, x54342, x54340);
  nand n54345(x54345, x54334, x54340);
  nand n54347(x54347, x53295, x53287);
  nand n54348(x54348, x53294, x54346);
  nand n54349(x54349, x54348, x54347);
  nand n54351(x54351, x53304, x53313);
  nand n54352(x54352, x53303, x53312);
  nand n54353(x54353, x54352, x54351);
  nand n54355(x54355, x53322, x54354);
  nand n54356(x54356, x53321, x54353);
  nand n54357(x54357, x54356, x54355);
  nand n54359(x54359, x54351, x54355);
  nand n54360(x54360, x53331, x53340);
  nand n54361(x54361, x53330, x53339);
  nand n54362(x54362, x54361, x54360);
  nand n54364(x54364, x53349, x54363);
  nand n54365(x54365, x53348, x54362);
  nand n54366(x54366, x54365, x54364);
  nand n54368(x54368, x54360, x54364);
  nand n54369(x54369, x53358, x53367);
  nand n54370(x54370, x53357, x53366);
  nand n54371(x54371, x54370, x54369);
  nand n54373(x54373, x53376, x54372);
  nand n54374(x54374, x53375, x54371);
  nand n54375(x54375, x54374, x54373);
  nand n54377(x54377, x54369, x54373);
  nand n54378(x54378, x53296, x53305);
  nand n54381(x54381, x54380, x54379);
  nand n54382(x54382, x54381, x54378);
  nand n54384(x54384, x53314, x54383);
  nand n54386(x54386, x54385, x54382);
  nand n54387(x54387, x54386, x54384);
  nand n54389(x54389, x53323, x53332);
  nand n54392(x54392, x54391, x54390);
  nand n54393(x54393, x54392, x54389);
  nand n54395(x54395, x53341, x54394);
  nand n54397(x54397, x54396, x54393);
  nand n54398(x54398, x54397, x54395);
  nand n54400(x54400, x53350, x53359);
  nand n54403(x54403, x54402, x54401);
  nand n54404(x54404, x54403, x54400);
  nand n54406(x54406, x53368, x54405);
  nand n54408(x54408, x54407, x54404);
  nand n54409(x54409, x54408, x54406);
  nand n54412(x54412, x53385, x53377);
  nand n54413(x54413, x53384, x54411);
  nand n54414(x54414, x54413, x54412);
  nand n54416(x54416, x53393, x53401);
  nand n54417(x54417, x53392, x53400);
  nand n54418(x54418, x54417, x54416);
  nand n54420(x54420, x53409, x54419);
  nand n54421(x54421, x53408, x54418);
  nand n54422(x54422, x54421, x54420);
  nand n54424(x54424, x53417, x53425);
  nand n54425(x54425, x53416, x53424);
  nand n54426(x54426, x54425, x54424);
  nand n54428(x54428, x53433, x54427);
  nand n54429(x54429, x53432, x54426);
  nand n54430(x54430, x54429, x54428);
  nand n54432(x54432, x53441, x53449);
  nand n54433(x54433, x53440, x53448);
  nand n54434(x54434, x54433, x54432);
  nand n54436(x54436, x53457, x54435);
  nand n54437(x54437, x53456, x54434);
  nand n54438(x54438, x54437, x54436);
  nand n54440(x54440, x85608, x85654);
  nand n54441(x54441, x50955, x52000);
  nand n54442(x54442, x54441, x54440);
  nand n54444(x54444, x85609, x85655);
  nand n54445(x54445, x52012, x52008);
  nand n54446(x54446, x54445, x54444);
  nand n54448(x54448, x85610, x85656);
  nand n54449(x54449, x52027, x52019);
  nand n54450(x54450, x54449, x54448);
  nand n54452(x54452, x85611, x85658);
  nand n54453(x54453, x53475, x52035);
  nand n54454(x54454, x54453, x54452);
  nand n54456(x54456, x85612, x85662);
  nand n54457(x54457, x53483, x52052);
  nand n54458(x54458, x54457, x54456);
  nand n54460(x54460, x85613, x85666);
  nand n54461(x54461, x53496, x52072);
  nand n54462(x54462, x54461, x54460);
  nand n54465(x54465, x53515, x85669);
  nand n54466(x54466, x53514, x52098);
  nand n54467(x54467, x54466, x54465);
  nand n54471(x54471, x53535, x85671);
  nand n54472(x54472, x53534, x52124);
  nand n54473(x54473, x54472, x54471);
  nand n54477(x54477, x85614, x85672);
  nand n54478(x54478, x52144, x53546);
  nand n54479(x54479, x54478, x54477);
  nand n54481(x54481, x53555, x85673);
  nand n54482(x54482, x53554, x52153);
  nand n54483(x54483, x54482, x54481);
  nand n54487(x54487, x52181, x85674);
  nand n54488(x54488, x53568, x53566);
  nand n54489(x54489, x54488, x54487);
  nand n54491(x54491, x53576, x85675);
  nand n54492(x54492, x53575, x52188);
  nand n54493(x54493, x54492, x54491);
  nand n54497(x54497, x52216, x85677);
  nand n54498(x54498, x53589, x53587);
  nand n54499(x54499, x54498, x54497);
  nand n54501(x54501, x53597, x85678);
  nand n54502(x54502, x53596, x52223);
  nand n54503(x54503, x54502, x54501);
  nand n54507(x54507, x85615, x85680);
  nand n54508(x54508, x53613, x53608);
  nand n54509(x54509, x54508, x54507);
  nand n54511(x54511, x53621, x85681);
  nand n54512(x54512, x53620, x52261);
  nand n54513(x54513, x54512, x54511);
  nand n54515(x54515, x53609, x85616);
  nand n54517(x54517, x54516, x53610);
  nand n54518(x54518, x54517, x54515);
  nand n54520(x54520, x85617, x85684);
  nand n54521(x54521, x53638, x53632);
  nand n54522(x54522, x54521, x54520);
  nand n54524(x54524, x53646, x85686);
  nand n54525(x54525, x53645, x52304);
  nand n54526(x54526, x54525, x54524);
  nand n54528(x54528, x53633, x85618);
  nand n54530(x54530, x54529, x53634);
  nand n54531(x54531, x54530, x54528);
  nand n54533(x54533, x85619, x53647);
  nand n54534(x54534, x53648, x54532);
  nand n54535(x54535, x54534, x54533);
  nand n54537(x54537, x85620, x85691);
  nand n54538(x54538, x53666, x53660);
  nand n54539(x54539, x54538, x54537);
  nand n54541(x54541, x53674, x85693);
  nand n54542(x54542, x53673, x52348);
  nand n54543(x54543, x54542, x54541);
  nand n54545(x54545, x53661, x85621);
  nand n54547(x54547, x54546, x53662);
  nand n54548(x54548, x54547, x54545);
  nand n54550(x54550, x85622, x53675);
  nand n54551(x54551, x53676, x54549);
  nand n54552(x54552, x54551, x54550);
  nand n54554(x54554, x53699, x85698);
  nand n54555(x54555, x53698, x53688);
  nand n54556(x54556, x54555, x54554);
  nand n54558(x54558, x53708, x85700);
  nand n54559(x54559, x53707, x52395);
  nand n54560(x54560, x54559, x54558);
  nand n54562(x54562, x53689, x53700);
  nand n54565(x54565, x54564, x54563);
  nand n54566(x54566, x54565, x54562);
  nand n54568(x54568, x85623, x53709);
  nand n54569(x54569, x53710, x54567);
  nand n54570(x54570, x54569, x54568);
  nand n54572(x54572, x53734, x85705);
  nand n54573(x54573, x53733, x53722);
  nand n54574(x54574, x54573, x54572);
  nand n54576(x54576, x53743, x85707);
  nand n54577(x54577, x53742, x52448);
  nand n54578(x54578, x54577, x54576);
  nand n54580(x54580, x53723, x53735);
  nand n54583(x54583, x54582, x54581);
  nand n54584(x54584, x54583, x54580);
  nand n54586(x54586, x53752, x53744);
  nand n54588(x54588, x54587, x54585);
  nand n54589(x54589, x54588, x54586);
  nand n54591(x54591, x53774, x85712);
  nand n54592(x54592, x53773, x53762);
  nand n54593(x54593, x54592, x54591);
  nand n54595(x54595, x53783, x85714);
  nand n54596(x54596, x53782, x52501);
  nand n54597(x54597, x54596, x54595);
  nand n54599(x54599, x53763, x53775);
  nand n54602(x54602, x54601, x54600);
  nand n54603(x54603, x54602, x54599);
  nand n54605(x54605, x53792, x53784);
  nand n54607(x54607, x54606, x54604);
  nand n54608(x54608, x54607, x54605);
  nand n54610(x54610, x53814, x85719);
  nand n54611(x54611, x53813, x53802);
  nand n54612(x54612, x54611, x54610);
  nand n54614(x54614, x85624, x85625);
  nand n54615(x54615, x52548, x52557);
  nand n54616(x54616, x54615, x54614);
  nand n54618(x54618, x53823, x54617);
  nand n54619(x54619, x53822, x54616);
  nand n54620(x54620, x54619, x54618);
  nand n54622(x54622, x54614, x54618);
  nand n54623(x54623, x53803, x53815);
  nand n54626(x54626, x54625, x54624);
  nand n54627(x54627, x54626, x54623);
  nand n54629(x54629, x53832, x53824);
  nand n54631(x54631, x54630, x54628);
  nand n54632(x54632, x54631, x54629);
  nand n54634(x54634, x53854, x85725);
  nand n54635(x54635, x53853, x53842);
  nand n54636(x54636, x54635, x54634);
  nand n54638(x54638, x52612, x85626);
  nand n54639(x54639, x53856, x52619);
  nand n54640(x54640, x54639, x54638);
  nand n54642(x54642, x53864, x54641);
  nand n54643(x54643, x53863, x54640);
  nand n54644(x54644, x54643, x54642);
  nand n54646(x54646, x54638, x54642);
  nand n54647(x54647, x53873, x85627);
  nand n54648(x54648, x53872, x51435);
  nand n54649(x54649, x54648, x54647);
  nand n54650(x54650, x53843, x53855);
  nand n54653(x54653, x54652, x54651);
  nand n54654(x54654, x54653, x54650);
  nand n54656(x54656, x53874, x53865);
  nand n54658(x54658, x54657, x54655);
  nand n54659(x54659, x54658, x54656);
  nand n54661(x54661, x53896, x85732);
  nand n54662(x54662, x53895, x53884);
  nand n54663(x54663, x54662, x54661);
  nand n54665(x54665, x52674, x85628);
  nand n54666(x54666, x53898, x52681);
  nand n54667(x54667, x54666, x54665);
  nand n54669(x54669, x53906, x54668);
  nand n54670(x54670, x53905, x54667);
  nand n54671(x54671, x54670, x54669);
  nand n54673(x54673, x54665, x54669);
  nand n54674(x54674, x53915, x85629);
  nand n54675(x54675, x53914, x52739);
  nand n54676(x54676, x54675, x54674);
  nand n54677(x54677, x53885, x53897);
  nand n54680(x54680, x54679, x54678);
  nand n54681(x54681, x54680, x54677);
  nand n54683(x54683, x53916, x53907);
  nand n54685(x54685, x54684, x54682);
  nand n54686(x54686, x54685, x54683);
  nand n54688(x54688, x53938, x85739);
  nand n54689(x54689, x53937, x53926);
  nand n54690(x54690, x54689, x54688);
  nand n54692(x54692, x85630, x85632);
  nand n54693(x54693, x53943, x52746);
  nand n54694(x54694, x54693, x54692);
  nand n54696(x54696, x53951, x54695);
  nand n54697(x54697, x53950, x54694);
  nand n54698(x54698, x54697, x54696);
  nand n54700(x54700, x54692, x54696);
  nand n54701(x54701, x53960, x85633);
  nand n54702(x54702, x53959, x52808);
  nand n54703(x54703, x54702, x54701);
  nand n54704(x54704, x53927, x53939);
  nand n54707(x54707, x54706, x54705);
  nand n54708(x54708, x54707, x54704);
  nand n54710(x54710, x85631, x54709);
  nand n54711(x54711, x53940, x54708);
  nand n54712(x54712, x54711, x54710);
  nand n54714(x54714, x54704, x54710);
  nand n54716(x54716, x53961, x53952);
  nand n54718(x54718, x54717, x54715);
  nand n54719(x54719, x54718, x54716);
  nand n54721(x54721, x53983, x85744);
  nand n54722(x54722, x53982, x53971);
  nand n54723(x54723, x54722, x54721);
  nand n54725(x54725, x85634, x85636);
  nand n54726(x54726, x53989, x52816);
  nand n54727(x54727, x54726, x54725);
  nand n54729(x54729, x53997, x54728);
  nand n54730(x54730, x53996, x54727);
  nand n54731(x54731, x54730, x54729);
  nand n54733(x54733, x54725, x54729);
  nand n54734(x54734, x54006, x85637);
  nand n54735(x54735, x54005, x54010);
  nand n54736(x54736, x54735, x54734);
  nand n54737(x54737, x53972, x53984);
  nand n54740(x54740, x54739, x54738);
  nand n54741(x54741, x54740, x54737);
  nand n54743(x54743, x85635, x54742);
  nand n54744(x54744, x53985, x54741);
  nand n54745(x54745, x54744, x54743);
  nand n54747(x54747, x54737, x54743);
  nand n54749(x54749, x54007, x53998);
  nand n54751(x54751, x54750, x54748);
  nand n54752(x54752, x54751, x54749);
  nand n54754(x54754, x85638, x54021);
  nand n54755(x54755, x54008, x54020);
  nand n54756(x54756, x54755, x54754);
  nand n54758(x54758, x54033, x54757);
  nand n54759(x54759, x54032, x54756);
  nand n54760(x54760, x54759, x54758);
  nand n54762(x54762, x54754, x54758);
  nand n54763(x54763, x85639, x85641);
  nand n54764(x54764, x54039, x52887);
  nand n54765(x54765, x54764, x54763);
  nand n54767(x54767, x54047, x54766);
  nand n54768(x54768, x54046, x54765);
  nand n54769(x54769, x54768, x54767);
  nand n54771(x54771, x54763, x54767);
  nand n54772(x54772, x54056, x85642);
  nand n54773(x54773, x54055, x54060);
  nand n54774(x54774, x54773, x54772);
  nand n54775(x54775, x54022, x54034);
  nand n54778(x54778, x54777, x54776);
  nand n54779(x54779, x54778, x54775);
  nand n54781(x54781, x85640, x54780);
  nand n54782(x54782, x54035, x54779);
  nand n54783(x54783, x54782, x54781);
  nand n54785(x54785, x54775, x54781);
  nand n54787(x54787, x54057, x54048);
  nand n54789(x54789, x54788, x54786);
  nand n54790(x54790, x54789, x54787);
  nand n54792(x54792, x85643, x54071);
  nand n54793(x54793, x54058, x54070);
  nand n54794(x54794, x54793, x54792);
  nand n54796(x54796, x54083, x54795);
  nand n54797(x54797, x54082, x54794);
  nand n54798(x54798, x54797, x54796);
  nand n54800(x54800, x54792, x54796);
  nand n54801(x54801, x54094, x85644);
  nand n54802(x54802, x54093, x52961);
  nand n54803(x54803, x54802, x54801);
  nand n54805(x54805, x54103, x54804);
  nand n54806(x54806, x54102, x54803);
  nand n54807(x54807, x54806, x54805);
  nand n54809(x54809, x54801, x54805);
  nand n54810(x54810, x54112, x85645);
  nand n54811(x54811, x54111, x54116);
  nand n54812(x54812, x54811, x54810);
  nand n54813(x54813, x54072, x54084);
  nand n54816(x54816, x54815, x54814);
  nand n54817(x54817, x54816, x54813);
  nand n54819(x54819, x54095, x54818);
  nand n54821(x54821, x54820, x54817);
  nand n54822(x54822, x54821, x54819);
  nand n54824(x54824, x54813, x54819);
  nand n54826(x54826, x54113, x54104);
  nand n54828(x54828, x54827, x54825);
  nand n54829(x54829, x54828, x54826);
  nand n54831(x54831, x85646, x54127);
  nand n54832(x54832, x54114, x54126);
  nand n54833(x54833, x54832, x54831);
  nand n54835(x54835, x54139, x54834);
  nand n54836(x54836, x54138, x54833);
  nand n54837(x54837, x54836, x54835);
  nand n54839(x54839, x54831, x54835);
  nand n54840(x54840, x54151, x85647);
  nand n54841(x54841, x54150, x53041);
  nand n54842(x54842, x54841, x54840);
  nand n54844(x54844, x54160, x54843);
  nand n54845(x54845, x54159, x54842);
  nand n54846(x54846, x54845, x54844);
  nand n54848(x54848, x54840, x54844);
  nand n54849(x54849, x54169, x54178);
  nand n54850(x54850, x54168, x54177);
  nand n54851(x54851, x54850, x54849);
  nand n54852(x54852, x54128, x54140);
  nand n54855(x54855, x54854, x54853);
  nand n54856(x54856, x54855, x54852);
  nand n54858(x54858, x54152, x54857);
  nand n54860(x54860, x54859, x54856);
  nand n54861(x54861, x54860, x54858);
  nand n54863(x54863, x54852, x54858);
  nand n54865(x54865, x54170, x54161);
  nand n54867(x54867, x54866, x54864);
  nand n54868(x54868, x54867, x54865);
  nand n54870(x54870, x54179, x54190);
  nand n54872(x54872, x54871, x54189);
  nand n54873(x54873, x54872, x54870);
  nand n54875(x54875, x54202, x54874);
  nand n54876(x54876, x54201, x54873);
  nand n54877(x54877, x54876, x54875);
  nand n54879(x54879, x54870, x54875);
  nand n54880(x54880, x54214, x85648);
  nand n54881(x54881, x54213, x53121);
  nand n54882(x54882, x54881, x54880);
  nand n54884(x54884, x54223, x54883);
  nand n54885(x54885, x54222, x54882);
  nand n54886(x54886, x54885, x54884);
  nand n54888(x54888, x54880, x54884);
  nand n54889(x54889, x54232, x54241);
  nand n54890(x54890, x54231, x54240);
  nand n54891(x54891, x54890, x54889);
  nand n54892(x54892, x54191, x54203);
  nand n54895(x54895, x54894, x54893);
  nand n54896(x54896, x54895, x54892);
  nand n54898(x54898, x54215, x54897);
  nand n54900(x54900, x54899, x54896);
  nand n54901(x54901, x54900, x54898);
  nand n54903(x54903, x54892, x54898);
  nand n54905(x54905, x54233, x54224);
  nand n54907(x54907, x54906, x54904);
  nand n54908(x54908, x54907, x54905);
  nand n54910(x54910, x54242, x54253);
  nand n54912(x54912, x54911, x54252);
  nand n54913(x54913, x54912, x54910);
  nand n54915(x54915, x54265, x54914);
  nand n54916(x54916, x54264, x54913);
  nand n54917(x54917, x54916, x54915);
  nand n54919(x54919, x54910, x54915);
  nand n54920(x54920, x54277, x54282);
  nand n54921(x54921, x54276, x54281);
  nand n54922(x54922, x54921, x54920);
  nand n54924(x54924, x54290, x54923);
  nand n54925(x54925, x54289, x54922);
  nand n54926(x54926, x54925, x54924);
  nand n54928(x54928, x54920, x54924);
  nand n54929(x54929, x54299, x54308);
  nand n54930(x54930, x54298, x54307);
  nand n54931(x54931, x54930, x54929);
  nand n54932(x54932, x54254, x54266);
  nand n54935(x54935, x54934, x54933);
  nand n54936(x54936, x54935, x54932);
  nand n54938(x54938, x54278, x54937);
  nand n54940(x54940, x54939, x54936);
  nand n54941(x54941, x54940, x54938);
  nand n54943(x54943, x54932, x54938);
  nand n54944(x54944, x85650, x54291);
  nand n54946(x54946, x54279, x54945);
  nand n54947(x54947, x54946, x54944);
  nand n54949(x54949, x54300, x54948);
  nand n54951(x54951, x54950, x54947);
  nand n54952(x54952, x54951, x54949);
  nand n54954(x54954, x54944, x54949);
  nand n54955(x54955, x54309, x54320);
  nand n54957(x54957, x54956, x54319);
  nand n54958(x54958, x54957, x54955);
  nand n54960(x54960, x54332, x54959);
  nand n54961(x54961, x54331, x54958);
  nand n54962(x54962, x54961, x54960);
  nand n54964(x54964, x54955, x54960);
  nand n54965(x54965, x54344, x54350);
  nand n54966(x54966, x54343, x54349);
  nand n54967(x54967, x54966, x54965);
  nand n54969(x54969, x54358, x54968);
  nand n54970(x54970, x54357, x54967);
  nand n54971(x54971, x54970, x54969);
  nand n54973(x54973, x54965, x54969);
  nand n54974(x54974, x54367, x54376);
  nand n54975(x54975, x54366, x54375);
  nand n54976(x54976, x54975, x54974);
  nand n54978(x54978, x85607, x54977);
  nand n54979(x54979, x51918, x54976);
  nand n54980(x54980, x54979, x54978);
  nand n54982(x54982, x54974, x54978);
  nand n54983(x54983, x54321, x54333);
  nand n54986(x54986, x54985, x54984);
  nand n54987(x54987, x54986, x54983);
  nand n54989(x54989, x54345, x54988);
  nand n54991(x54991, x54990, x54987);
  nand n54992(x54992, x54991, x54989);
  nand n54994(x54994, x85651, x54359);
  nand n54996(x54996, x54347, x54995);
  nand n54997(x54997, x54996, x54994);
  nand n54999(x54999, x54368, x54998);
  nand n55001(x55001, x55000, x54997);
  nand n55002(x55002, x55001, x54999);
  nand n55004(x55004, x54377, x54388);
  nand n55006(x55006, x55005, x54387);
  nand n55007(x55007, x55006, x55004);
  nand n55009(x55009, x54399, x55008);
  nand n55010(x55010, x54398, x55007);
  nand n55011(x55011, x55010, x55009);
  nand n55013(x55013, x54410, x54415);
  nand n55014(x55014, x54409, x54414);
  nand n55015(x55015, x55014, x55013);
  nand n55017(x55017, x54423, x55016);
  nand n55018(x55018, x54422, x55015);
  nand n55019(x55019, x55018, x55017);
  nand n55021(x55021, x54431, x54439);
  nand n55022(x55022, x54430, x54438);
  nand n55023(x55023, x55022, x55021);
  nand n55025(x55025, x53461, x55024);
  nand n55026(x55026, x53460, x55023);
  nand n55027(x55027, x55026, x55025);
  nand n55029(x55029, x85652, x85653);
  nand n55030(x55030, x51983, x51992);
  nand n55031(x55031, x55030, x55029);
  nand n55032(x55032, x54443, x51993);
  nand n55033(x55033, x54442, x53462);
  nand n55034(x55034, x55033, x55032);
  nand n55035(x55035, x54447, x52001);
  nand n55036(x55036, x54446, x53463);
  nand n55037(x55037, x55036, x55035);
  nand n55039(x55039, x54451, x85763);
  nand n55040(x55040, x54450, x53467);
  nand n55041(x55041, x55040, x55039);
  nand n55043(x55043, x85657, x85764);
  nand n55044(x55044, x53464, x54448);
  nand n55045(x55045, x55044, x55043);
  nand n55046(x55046, x54455, x85765);
  nand n55047(x55047, x54454, x53472);
  nand n55048(x55048, x55047, x55046);
  nand n55050(x55050, x85659, x85767);
  nand n55051(x55051, x53468, x54452);
  nand n55052(x55052, x55051, x55050);
  nand n55053(x55053, x85660, x85661);
  nand n55054(x55054, x53473, x53480);
  nand n55055(x55055, x55054, x55053);
  nand n55057(x55057, x54459, x55056);
  nand n55058(x55058, x54458, x55055);
  nand n55059(x55059, x55058, x55057);
  nand n55061(x55061, x55053, x55057);
  nand n55062(x55062, x85663, x85768);
  nand n55063(x55063, x53476, x54456);
  nand n55064(x55064, x55063, x55062);
  nand n55065(x55065, x85664, x85665);
  nand n55066(x55066, x53481, x53492);
  nand n55067(x55067, x55066, x55065);
  nand n55069(x55069, x54463, x55068);
  nand n55070(x55070, x54462, x55067);
  nand n55071(x55071, x55070, x55069);
  nand n55073(x55073, x55065, x55069);
  nand n55074(x55074, x53493, x85769);
  nand n55075(x55075, x54464, x54460);
  nand n55076(x55076, x55075, x55074);
  nand n55077(x55077, x85667, x85668);
  nand n55078(x55078, x53494, x53506);
  nand n55079(x55079, x55078, x55077);
  nand n55081(x55081, x54468, x55080);
  nand n55082(x55082, x54467, x55079);
  nand n55083(x55083, x55082, x55081);
  nand n55085(x55085, x55077, x55081);
  nand n55086(x55086, x53507, x85770);
  nand n55087(x55087, x54469, x54465);
  nand n55088(x55088, x55087, x55086);
  nand n55089(x55089, x53516, x85670);
  nand n55090(x55090, x54470, x53526);
  nand n55091(x55091, x55090, x55089);
  nand n55093(x55093, x54474, x55092);
  nand n55094(x55094, x54473, x55091);
  nand n55095(x55095, x55094, x55093);
  nand n55097(x55097, x55089, x55093);
  nand n55098(x55098, x53527, x85771);
  nand n55099(x55099, x54475, x54471);
  nand n55100(x55100, x55099, x55098);
  nand n55101(x55101, x53536, x54480);
  nand n55102(x55102, x54476, x54479);
  nand n55103(x55103, x55102, x55101);
  nand n55105(x55105, x54484, x55104);
  nand n55106(x55106, x54483, x55103);
  nand n55107(x55107, x55106, x55105);
  nand n55109(x55109, x55101, x55105);
  nand n55110(x55110, x53547, x85773);
  nand n55111(x55111, x54485, x54481);
  nand n55112(x55112, x55111, x55110);
  nand n55114(x55114, x53556, x54490);
  nand n55115(x55115, x54486, x54489);
  nand n55116(x55116, x55115, x55114);
  nand n55118(x55118, x54494, x55117);
  nand n55119(x55119, x54493, x55116);
  nand n55120(x55120, x55119, x55118);
  nand n55122(x55122, x55114, x55118);
  nand n55123(x55123, x53567, x85775);
  nand n55124(x55124, x54495, x54491);
  nand n55125(x55125, x55124, x55123);
  nand n55127(x55127, x53577, x54500);
  nand n55128(x55128, x54496, x54499);
  nand n55129(x55129, x55128, x55127);
  nand n55131(x55131, x54504, x55130);
  nand n55132(x55132, x54503, x55129);
  nand n55133(x55133, x55132, x55131);
  nand n55135(x55135, x55127, x55131);
  nand n55136(x55136, x53588, x85777);
  nand n55137(x55137, x54505, x54501);
  nand n55138(x55138, x55137, x55136);
  nand n55140(x55140, x53598, x54510);
  nand n55141(x55141, x54506, x54509);
  nand n55142(x55142, x55141, x55140);
  nand n55144(x55144, x54514, x55143);
  nand n55145(x55145, x54513, x55142);
  nand n55146(x55146, x55145, x55144);
  nand n55148(x55148, x55140, x55144);
  nand n55149(x55149, x85683, x85779);
  nand n55150(x55150, x54518, x54511);
  nand n55151(x55151, x55150, x55149);
  nand n55153(x55153, x53622, x54523);
  nand n55154(x55154, x54519, x54522);
  nand n55155(x55155, x55154, x55153);
  nand n55157(x55157, x54527, x55156);
  nand n55158(x55158, x54526, x55155);
  nand n55159(x55159, x55158, x55157);
  nand n55161(x55161, x55153, x55157);
  nand n55162(x55162, x85685, x85780);
  nand n55163(x55163, x54520, x54515);
  nand n55164(x55164, x55163, x55162);
  nand n55166(x55166, x85688, x85782);
  nand n55167(x55167, x54531, x54524);
  nand n55168(x55168, x55167, x55166);
  nand n55170(x55170, x54536, x54540);
  nand n55171(x55171, x54535, x54539);
  nand n55172(x55172, x55171, x55170);
  nand n55174(x55174, x54544, x55173);
  nand n55175(x55175, x54543, x55172);
  nand n55176(x55176, x55175, x55174);
  nand n55178(x55178, x55170, x55174);
  nand n55179(x55179, x85689, x85690);
  nand n55180(x55180, x54528, x54533);
  nand n55181(x55181, x55180, x55179);
  nand n55183(x55183, x85692, x55182);
  nand n55184(x55184, x54537, x55181);
  nand n55185(x55185, x55184, x55183);
  nand n55187(x55187, x55179, x55183);
  nand n55188(x55188, x85695, x85784);
  nand n55189(x55189, x54548, x54541);
  nand n55190(x55190, x55189, x55188);
  nand n55192(x55192, x54553, x54557);
  nand n55193(x55193, x54552, x54556);
  nand n55194(x55194, x55193, x55192);
  nand n55196(x55196, x54561, x55195);
  nand n55197(x55197, x54560, x55194);
  nand n55198(x55198, x55197, x55196);
  nand n55200(x55200, x55192, x55196);
  nand n55201(x55201, x85696, x85697);
  nand n55202(x55202, x54545, x54550);
  nand n55203(x55203, x55202, x55201);
  nand n55205(x55205, x85699, x55204);
  nand n55206(x55206, x54554, x55203);
  nand n55207(x55207, x55206, x55205);
  nand n55209(x55209, x55201, x55205);
  nand n55210(x55210, x85702, x85786);
  nand n55211(x55211, x54566, x54558);
  nand n55212(x55212, x55211, x55210);
  nand n55214(x55214, x54571, x54575);
  nand n55215(x55215, x54570, x54574);
  nand n55216(x55216, x55215, x55214);
  nand n55218(x55218, x54579, x55217);
  nand n55219(x55219, x54578, x55216);
  nand n55220(x55220, x55219, x55218);
  nand n55222(x55222, x55214, x55218);
  nand n55223(x55223, x85703, x85704);
  nand n55224(x55224, x54562, x54568);
  nand n55225(x55225, x55224, x55223);
  nand n55227(x55227, x85706, x55226);
  nand n55228(x55228, x54572, x55225);
  nand n55229(x55229, x55228, x55227);
  nand n55231(x55231, x55223, x55227);
  nand n55232(x55232, x85709, x85788);
  nand n55233(x55233, x54584, x54576);
  nand n55234(x55234, x55233, x55232);
  nand n55236(x55236, x54590, x54594);
  nand n55237(x55237, x54589, x54593);
  nand n55238(x55238, x55237, x55236);
  nand n55240(x55240, x54598, x55239);
  nand n55241(x55241, x54597, x55238);
  nand n55242(x55242, x55241, x55240);
  nand n55244(x55244, x55236, x55240);
  nand n55245(x55245, x85710, x85711);
  nand n55246(x55246, x54580, x54586);
  nand n55247(x55247, x55246, x55245);
  nand n55249(x55249, x85713, x55248);
  nand n55250(x55250, x54591, x55247);
  nand n55251(x55251, x55250, x55249);
  nand n55253(x55253, x55245, x55249);
  nand n55254(x55254, x85716, x85790);
  nand n55255(x55255, x54603, x54595);
  nand n55256(x55256, x55255, x55254);
  nand n55258(x55258, x54609, x54613);
  nand n55259(x55259, x54608, x54612);
  nand n55260(x55260, x55259, x55258);
  nand n55262(x55262, x54621, x55261);
  nand n55263(x55263, x54620, x55260);
  nand n55264(x55264, x55263, x55262);
  nand n55266(x55266, x55258, x55262);
  nand n55267(x55267, x85717, x85718);
  nand n55268(x55268, x54599, x54605);
  nand n55269(x55269, x55268, x55267);
  nand n55271(x55271, x85720, x55270);
  nand n55272(x55272, x54610, x55269);
  nand n55273(x55273, x55272, x55271);
  nand n55275(x55275, x55267, x55271);
  nand n55277(x55277, x85722, x54622);
  nand n55278(x55278, x54627, x55276);
  nand n55279(x55279, x55278, x55277);
  nand n55281(x55281, x54633, x54637);
  nand n55282(x55282, x54632, x54636);
  nand n55283(x55283, x55282, x55281);
  nand n55285(x55285, x54645, x55284);
  nand n55286(x55286, x54644, x55283);
  nand n55287(x55287, x55286, x55285);
  nand n55289(x55289, x55281, x55285);
  nand n55290(x55290, x85723, x85724);
  nand n55291(x55291, x54623, x54629);
  nand n55292(x55292, x55291, x55290);
  nand n55294(x55294, x85726, x55293);
  nand n55295(x55295, x54634, x55292);
  nand n55296(x55296, x55295, x55294);
  nand n55298(x55298, x55290, x55294);
  nand n55299(x55299, x54646, x85728);
  nand n55301(x55301, x55300, x54647);
  nand n55302(x55302, x55301, x55299);
  nand n55304(x55304, x85729, x55303);
  nand n55305(x55305, x54654, x55302);
  nand n55306(x55306, x55305, x55304);
  nand n55308(x55308, x55299, x55304);
  nand n55309(x55309, x54660, x54664);
  nand n55310(x55310, x54659, x54663);
  nand n55311(x55311, x55310, x55309);
  nand n55313(x55313, x54672, x55312);
  nand n55314(x55314, x54671, x55311);
  nand n55315(x55315, x55314, x55313);
  nand n55317(x55317, x55309, x55313);
  nand n55318(x55318, x85730, x85731);
  nand n55319(x55319, x54650, x54656);
  nand n55320(x55320, x55319, x55318);
  nand n55322(x55322, x85733, x55321);
  nand n55323(x55323, x54661, x55320);
  nand n55324(x55324, x55323, x55322);
  nand n55326(x55326, x55318, x55322);
  nand n55327(x55327, x54673, x85735);
  nand n55329(x55329, x55328, x54674);
  nand n55330(x55330, x55329, x55327);
  nand n55332(x55332, x85736, x55331);
  nand n55333(x55333, x54681, x55330);
  nand n55334(x55334, x55333, x55332);
  nand n55336(x55336, x55327, x55332);
  nand n55337(x55337, x54687, x54691);
  nand n55338(x55338, x54686, x54690);
  nand n55339(x55339, x55338, x55337);
  nand n55341(x55341, x54699, x55340);
  nand n55342(x55342, x54698, x55339);
  nand n55343(x55343, x55342, x55341);
  nand n55345(x55345, x55337, x55341);
  nand n55346(x55346, x85737, x85738);
  nand n55347(x55347, x54677, x54683);
  nand n55348(x55348, x55347, x55346);
  nand n55350(x55350, x85740, x55349);
  nand n55351(x55351, x54688, x55348);
  nand n55352(x55352, x55351, x55350);
  nand n55354(x55354, x55346, x55350);
  nand n55355(x55355, x54700, x85742);
  nand n55357(x55357, x55356, x54701);
  nand n55358(x55358, x55357, x55355);
  nand n55360(x55360, x54713, x55359);
  nand n55361(x55361, x54712, x55358);
  nand n55362(x55362, x55361, x55360);
  nand n55364(x55364, x55355, x55360);
  nand n55365(x55365, x54720, x54724);
  nand n55366(x55366, x54719, x54723);
  nand n55367(x55367, x55366, x55365);
  nand n55369(x55369, x54732, x55368);
  nand n55370(x55370, x54731, x55367);
  nand n55371(x55371, x55370, x55369);
  nand n55373(x55373, x55365, x55369);
  nand n55374(x55374, x54714, x85743);
  nand n55376(x55376, x55375, x54716);
  nand n55377(x55377, x55376, x55374);
  nand n55379(x55379, x85745, x55378);
  nand n55380(x55380, x54721, x55377);
  nand n55381(x55381, x55380, x55379);
  nand n55383(x55383, x55374, x55379);
  nand n55384(x55384, x54733, x85747);
  nand n55386(x55386, x55385, x54734);
  nand n55387(x55387, x55386, x55384);
  nand n55389(x55389, x54746, x55388);
  nand n55390(x55390, x54745, x55387);
  nand n55391(x55391, x55390, x55389);
  nand n55393(x55393, x55384, x55389);
  nand n55394(x55394, x54753, x54761);
  nand n55395(x55395, x54752, x54760);
  nand n55396(x55396, x55395, x55394);
  nand n55398(x55398, x54770, x55397);
  nand n55399(x55399, x54769, x55396);
  nand n55400(x55400, x55399, x55398);
  nand n55402(x55402, x55394, x55398);
  nand n55403(x55403, x54747, x85748);
  nand n55405(x55405, x55404, x54749);
  nand n55406(x55406, x55405, x55403);
  nand n55408(x55408, x54762, x55407);
  nand n55410(x55410, x55409, x55406);
  nand n55411(x55411, x55410, x55408);
  nand n55413(x55413, x55403, x55408);
  nand n55414(x55414, x54771, x85750);
  nand n55416(x55416, x55415, x54772);
  nand n55417(x55417, x55416, x55414);
  nand n55419(x55419, x54784, x55418);
  nand n55420(x55420, x54783, x55417);
  nand n55421(x55421, x55420, x55419);
  nand n55423(x55423, x55414, x55419);
  nand n55424(x55424, x54791, x54799);
  nand n55425(x55425, x54790, x54798);
  nand n55426(x55426, x55425, x55424);
  nand n55428(x55428, x54808, x55427);
  nand n55429(x55429, x54807, x55426);
  nand n55430(x55430, x55429, x55428);
  nand n55432(x55432, x55424, x55428);
  nand n55433(x55433, x54785, x85751);
  nand n55435(x55435, x55434, x54787);
  nand n55436(x55436, x55435, x55433);
  nand n55438(x55438, x54800, x55437);
  nand n55440(x55440, x55439, x55436);
  nand n55441(x55441, x55440, x55438);
  nand n55443(x55443, x55433, x55438);
  nand n55444(x55444, x54809, x85753);
  nand n55446(x55446, x55445, x54810);
  nand n55447(x55447, x55446, x55444);
  nand n55449(x55449, x54823, x55448);
  nand n55450(x55450, x54822, x55447);
  nand n55451(x55451, x55450, x55449);
  nand n55453(x55453, x55444, x55449);
  nand n55454(x55454, x54830, x54838);
  nand n55455(x55455, x54829, x54837);
  nand n55456(x55456, x55455, x55454);
  nand n55458(x55458, x54847, x55457);
  nand n55459(x55459, x54846, x55456);
  nand n55460(x55460, x55459, x55458);
  nand n55462(x55462, x55454, x55458);
  nand n55463(x55463, x54824, x85754);
  nand n55465(x55465, x55464, x54826);
  nand n55466(x55466, x55465, x55463);
  nand n55468(x55468, x54839, x55467);
  nand n55470(x55470, x55469, x55466);
  nand n55471(x55471, x55470, x55468);
  nand n55473(x55473, x55463, x55468);
  nand n55474(x55474, x54848, x85756);
  nand n55476(x55476, x55475, x54849);
  nand n55477(x55477, x55476, x55474);
  nand n55479(x55479, x54862, x55478);
  nand n55480(x55480, x54861, x55477);
  nand n55481(x55481, x55480, x55479);
  nand n55483(x55483, x55474, x55479);
  nand n55484(x55484, x54869, x54878);
  nand n55485(x55485, x54868, x54877);
  nand n55486(x55486, x55485, x55484);
  nand n55488(x55488, x54887, x55487);
  nand n55489(x55489, x54886, x55486);
  nand n55490(x55490, x55489, x55488);
  nand n55492(x55492, x55484, x55488);
  nand n55493(x55493, x54863, x85757);
  nand n55495(x55495, x55494, x54865);
  nand n55496(x55496, x55495, x55493);
  nand n55498(x55498, x54879, x55497);
  nand n55500(x55500, x55499, x55496);
  nand n55501(x55501, x55500, x55498);
  nand n55503(x55503, x55493, x55498);
  nand n55504(x55504, x54888, x85759);
  nand n55506(x55506, x55505, x54889);
  nand n55507(x55507, x55506, x55504);
  nand n55509(x55509, x54902, x55508);
  nand n55510(x55510, x54901, x55507);
  nand n55511(x55511, x55510, x55509);
  nand n55513(x55513, x55504, x55509);
  nand n55514(x55514, x54909, x54918);
  nand n55515(x55515, x54908, x54917);
  nand n55516(x55516, x55515, x55514);
  nand n55518(x55518, x54927, x55517);
  nand n55519(x55519, x54926, x55516);
  nand n55520(x55520, x55519, x55518);
  nand n55522(x55522, x55514, x55518);
  nand n55523(x55523, x54903, x85760);
  nand n55525(x55525, x55524, x54905);
  nand n55526(x55526, x55525, x55523);
  nand n55528(x55528, x54919, x55527);
  nand n55530(x55530, x55529, x55526);
  nand n55531(x55531, x55530, x55528);
  nand n55533(x55533, x55523, x55528);
  nand n55534(x55534, x54928, x85762);
  nand n55536(x55536, x55535, x54929);
  nand n55537(x55537, x55536, x55534);
  nand n55539(x55539, x54942, x55538);
  nand n55540(x55540, x54941, x55537);
  nand n55541(x55541, x55540, x55539);
  nand n55543(x55543, x55534, x55539);
  nand n55544(x55544, x54953, x54963);
  nand n55545(x55545, x54952, x54962);
  nand n55546(x55546, x55545, x55544);
  nand n55548(x55548, x54972, x55547);
  nand n55549(x55549, x54971, x55546);
  nand n55550(x55550, x55549, x55548);
  nand n55552(x55552, x55544, x55548);
  nand n55553(x55553, x54943, x54954);
  nand n55556(x55556, x55555, x55554);
  nand n55557(x55557, x55556, x55553);
  nand n55559(x55559, x54964, x55558);
  nand n55561(x55561, x55560, x55557);
  nand n55562(x55562, x55561, x55559);
  nand n55564(x55564, x54973, x54982);
  nand n55567(x55567, x55566, x55565);
  nand n55568(x55568, x55567, x55564);
  nand n55570(x55570, x54993, x55569);
  nand n55571(x55571, x54992, x55568);
  nand n55572(x55572, x55571, x55570);
  nand n55574(x55574, x55003, x55012);
  nand n55575(x55575, x55002, x55011);
  nand n55576(x55576, x55575, x55574);
  nand n55578(x55578, x55020, x55577);
  nand n55579(x55579, x55019, x55576);
  nand n55580(x55580, x55579, x55578);
  nand n55582(x55582, x55038, x85793);
  nand n55583(x55583, x55037, x54440);
  nand n55584(x55584, x55583, x55582);
  nand n55585(x55585, x55042, x85795);
  nand n55586(x55586, x55041, x54444);
  nand n55587(x55587, x55586, x55585);
  nand n55588(x55588, x55049, x85797);
  nand n55589(x55589, x55048, x55045);
  nand n55590(x55590, x55589, x55588);
  nand n55591(x55591, x85766, x85798);
  nand n55592(x55592, x55046, x55043);
  nand n55593(x55593, x55592, x55591);
  nand n55595(x55595, x55060, x85800);
  nand n55596(x55596, x55059, x55052);
  nand n55597(x55597, x55596, x55595);
  nand n55598(x55598, x55061, x85802);
  nand n55600(x55600, x55599, x55050);
  nand n55601(x55601, x55600, x55598);
  nand n55603(x55603, x55072, x85804);
  nand n55604(x55604, x55071, x55064);
  nand n55605(x55605, x55604, x55603);
  nand n55606(x55606, x55073, x85806);
  nand n55608(x55608, x55607, x55062);
  nand n55609(x55609, x55608, x55606);
  nand n55611(x55611, x55084, x85808);
  nand n55612(x55612, x55083, x55076);
  nand n55613(x55613, x55612, x55611);
  nand n55614(x55614, x55085, x85810);
  nand n55616(x55616, x55615, x55074);
  nand n55617(x55617, x55616, x55614);
  nand n55619(x55619, x55096, x85812);
  nand n55620(x55620, x55095, x55088);
  nand n55621(x55621, x55620, x55619);
  nand n55622(x55622, x55097, x85814);
  nand n55624(x55624, x55623, x55086);
  nand n55625(x55625, x55624, x55622);
  nand n55627(x55627, x55108, x85816);
  nand n55628(x55628, x55107, x55100);
  nand n55629(x55629, x55628, x55627);
  nand n55630(x55630, x55109, x85818);
  nand n55632(x55632, x55631, x55098);
  nand n55633(x55633, x55632, x55630);
  nand n55635(x55635, x85772, x55113);
  nand n55636(x55636, x54477, x55112);
  nand n55637(x55637, x55636, x55635);
  nand n55639(x55639, x55121, x55638);
  nand n55640(x55640, x55120, x55637);
  nand n55641(x55641, x55640, x55639);
  nand n55643(x55643, x55635, x55639);
  nand n55644(x55644, x55122, x85820);
  nand n55646(x55646, x55645, x55110);
  nand n55647(x55647, x55646, x55644);
  nand n55649(x55649, x85774, x55126);
  nand n55650(x55650, x54487, x55125);
  nand n55651(x55651, x55650, x55649);
  nand n55653(x55653, x55134, x55652);
  nand n55654(x55654, x55133, x55651);
  nand n55655(x55655, x55654, x55653);
  nand n55657(x55657, x55649, x55653);
  nand n55658(x55658, x55135, x85822);
  nand n55660(x55660, x55659, x55123);
  nand n55661(x55661, x55660, x55658);
  nand n55663(x55663, x85776, x55139);
  nand n55664(x55664, x54497, x55138);
  nand n55665(x55665, x55664, x55663);
  nand n55667(x55667, x55147, x55666);
  nand n55668(x55668, x55146, x55665);
  nand n55669(x55669, x55668, x55667);
  nand n55671(x55671, x55663, x55667);
  nand n55672(x55672, x55148, x85824);
  nand n55674(x55674, x55673, x55136);
  nand n55675(x55675, x55674, x55672);
  nand n55677(x55677, x85778, x55152);
  nand n55678(x55678, x54507, x55151);
  nand n55679(x55679, x55678, x55677);
  nand n55681(x55681, x55160, x55680);
  nand n55682(x55682, x55159, x55679);
  nand n55683(x55683, x55682, x55681);
  nand n55685(x55685, x55677, x55681);
  nand n55686(x55686, x55161, x85826);
  nand n55688(x55688, x55687, x55149);
  nand n55689(x55689, x55688, x55686);
  nand n55691(x55691, x55165, x55169);
  nand n55692(x55692, x55164, x55168);
  nand n55693(x55693, x55692, x55691);
  nand n55695(x55695, x55177, x55694);
  nand n55696(x55696, x55176, x55693);
  nand n55697(x55697, x55696, x55695);
  nand n55699(x55699, x55691, x55695);
  nand n55700(x55700, x85781, x85783);
  nand n55701(x55701, x55162, x55166);
  nand n55702(x55702, x55701, x55700);
  nand n55704(x55704, x55178, x55703);
  nand n55706(x55706, x55705, x55702);
  nand n55707(x55707, x55706, x55704);
  nand n55709(x55709, x55700, x55704);
  nand n55710(x55710, x55186, x55191);
  nand n55711(x55711, x55185, x55190);
  nand n55712(x55712, x55711, x55710);
  nand n55714(x55714, x55199, x55713);
  nand n55715(x55715, x55198, x55712);
  nand n55716(x55716, x55715, x55714);
  nand n55718(x55718, x55710, x55714);
  nand n55719(x55719, x55187, x85785);
  nand n55721(x55721, x55720, x55188);
  nand n55722(x55722, x55721, x55719);
  nand n55724(x55724, x55200, x55723);
  nand n55726(x55726, x55725, x55722);
  nand n55727(x55727, x55726, x55724);
  nand n55729(x55729, x55719, x55724);
  nand n55730(x55730, x55208, x55213);
  nand n55731(x55731, x55207, x55212);
  nand n55732(x55732, x55731, x55730);
  nand n55734(x55734, x55221, x55733);
  nand n55735(x55735, x55220, x55732);
  nand n55736(x55736, x55735, x55734);
  nand n55738(x55738, x55730, x55734);
  nand n55739(x55739, x55209, x85787);
  nand n55741(x55741, x55740, x55210);
  nand n55742(x55742, x55741, x55739);
  nand n55744(x55744, x55222, x55743);
  nand n55746(x55746, x55745, x55742);
  nand n55747(x55747, x55746, x55744);
  nand n55749(x55749, x55739, x55744);
  nand n55750(x55750, x55230, x55235);
  nand n55751(x55751, x55229, x55234);
  nand n55752(x55752, x55751, x55750);
  nand n55754(x55754, x55243, x55753);
  nand n55755(x55755, x55242, x55752);
  nand n55756(x55756, x55755, x55754);
  nand n55758(x55758, x55750, x55754);
  nand n55759(x55759, x55231, x85789);
  nand n55761(x55761, x55760, x55232);
  nand n55762(x55762, x55761, x55759);
  nand n55764(x55764, x55244, x55763);
  nand n55766(x55766, x55765, x55762);
  nand n55767(x55767, x55766, x55764);
  nand n55769(x55769, x55759, x55764);
  nand n55770(x55770, x55252, x55257);
  nand n55771(x55771, x55251, x55256);
  nand n55772(x55772, x55771, x55770);
  nand n55774(x55774, x55265, x55773);
  nand n55775(x55775, x55264, x55772);
  nand n55776(x55776, x55775, x55774);
  nand n55778(x55778, x55770, x55774);
  nand n55779(x55779, x55253, x85791);
  nand n55781(x55781, x55780, x55254);
  nand n55782(x55782, x55781, x55779);
  nand n55784(x55784, x55266, x55783);
  nand n55786(x55786, x55785, x55782);
  nand n55787(x55787, x55786, x55784);
  nand n55789(x55789, x55779, x55784);
  nand n55790(x55790, x55274, x55280);
  nand n55791(x55791, x55273, x55279);
  nand n55792(x55792, x55791, x55790);
  nand n55794(x55794, x55288, x55793);
  nand n55795(x55795, x55287, x55792);
  nand n55796(x55796, x55795, x55794);
  nand n55798(x55798, x55790, x55794);
  nand n55799(x55799, x55275, x85792);
  nand n55801(x55801, x55800, x55277);
  nand n55802(x55802, x55801, x55799);
  nand n55804(x55804, x55289, x55803);
  nand n55806(x55806, x55805, x55802);
  nand n55807(x55807, x55806, x55804);
  nand n55809(x55809, x55799, x55804);
  nand n55810(x55810, x55297, x55307);
  nand n55811(x55811, x55296, x55306);
  nand n55812(x55812, x55811, x55810);
  nand n55814(x55814, x55316, x55813);
  nand n55815(x55815, x55315, x55812);
  nand n55816(x55816, x55815, x55814);
  nand n55818(x55818, x55810, x55814);
  nand n55819(x55819, x55298, x55308);
  nand n55822(x55822, x55821, x55820);
  nand n55823(x55823, x55822, x55819);
  nand n55825(x55825, x55317, x55824);
  nand n55827(x55827, x55826, x55823);
  nand n55828(x55828, x55827, x55825);
  nand n55830(x55830, x55819, x55825);
  nand n55831(x55831, x55325, x55335);
  nand n55832(x55832, x55324, x55334);
  nand n55833(x55833, x55832, x55831);
  nand n55835(x55835, x55344, x55834);
  nand n55836(x55836, x55343, x55833);
  nand n55837(x55837, x55836, x55835);
  nand n55839(x55839, x55831, x55835);
  nand n55840(x55840, x55326, x55336);
  nand n55843(x55843, x55842, x55841);
  nand n55844(x55844, x55843, x55840);
  nand n55846(x55846, x55345, x55845);
  nand n55848(x55848, x55847, x55844);
  nand n55849(x55849, x55848, x55846);
  nand n55851(x55851, x55840, x55846);
  nand n55852(x55852, x55353, x55363);
  nand n55853(x55853, x55352, x55362);
  nand n55854(x55854, x55853, x55852);
  nand n55856(x55856, x55372, x55855);
  nand n55857(x55857, x55371, x55854);
  nand n55858(x55858, x55857, x55856);
  nand n55860(x55860, x55852, x55856);
  nand n55861(x55861, x55354, x55364);
  nand n55864(x55864, x55863, x55862);
  nand n55865(x55865, x55864, x55861);
  nand n55867(x55867, x55373, x55866);
  nand n55869(x55869, x55868, x55865);
  nand n55870(x55870, x55869, x55867);
  nand n55872(x55872, x55861, x55867);
  nand n55873(x55873, x55382, x55392);
  nand n55874(x55874, x55381, x55391);
  nand n55875(x55875, x55874, x55873);
  nand n55877(x55877, x55401, x55876);
  nand n55878(x55878, x55400, x55875);
  nand n55879(x55879, x55878, x55877);
  nand n55881(x55881, x55873, x55877);
  nand n55882(x55882, x55383, x55393);
  nand n55885(x55885, x55884, x55883);
  nand n55886(x55886, x55885, x55882);
  nand n55888(x55888, x55402, x55887);
  nand n55890(x55890, x55889, x55886);
  nand n55891(x55891, x55890, x55888);
  nand n55893(x55893, x55882, x55888);
  nand n55894(x55894, x55412, x55422);
  nand n55895(x55895, x55411, x55421);
  nand n55896(x55896, x55895, x55894);
  nand n55898(x55898, x55431, x55897);
  nand n55899(x55899, x55430, x55896);
  nand n55900(x55900, x55899, x55898);
  nand n55902(x55902, x55894, x55898);
  nand n55903(x55903, x55413, x55423);
  nand n55906(x55906, x55905, x55904);
  nand n55907(x55907, x55906, x55903);
  nand n55909(x55909, x55432, x55908);
  nand n55911(x55911, x55910, x55907);
  nand n55912(x55912, x55911, x55909);
  nand n55914(x55914, x55903, x55909);
  nand n55915(x55915, x55442, x55452);
  nand n55916(x55916, x55441, x55451);
  nand n55917(x55917, x55916, x55915);
  nand n55919(x55919, x55461, x55918);
  nand n55920(x55920, x55460, x55917);
  nand n55921(x55921, x55920, x55919);
  nand n55923(x55923, x55915, x55919);
  nand n55924(x55924, x55443, x55453);
  nand n55927(x55927, x55926, x55925);
  nand n55928(x55928, x55927, x55924);
  nand n55930(x55930, x55462, x55929);
  nand n55932(x55932, x55931, x55928);
  nand n55933(x55933, x55932, x55930);
  nand n55935(x55935, x55924, x55930);
  nand n55936(x55936, x55472, x55482);
  nand n55937(x55937, x55471, x55481);
  nand n55938(x55938, x55937, x55936);
  nand n55940(x55940, x55491, x55939);
  nand n55941(x55941, x55490, x55938);
  nand n55942(x55942, x55941, x55940);
  nand n55944(x55944, x55936, x55940);
  nand n55945(x55945, x55473, x55483);
  nand n55948(x55948, x55947, x55946);
  nand n55949(x55949, x55948, x55945);
  nand n55951(x55951, x55492, x55950);
  nand n55953(x55953, x55952, x55949);
  nand n55954(x55954, x55953, x55951);
  nand n55956(x55956, x55945, x55951);
  nand n55957(x55957, x55502, x55512);
  nand n55958(x55958, x55501, x55511);
  nand n55959(x55959, x55958, x55957);
  nand n55961(x55961, x55521, x55960);
  nand n55962(x55962, x55520, x55959);
  nand n55963(x55963, x55962, x55961);
  nand n55965(x55965, x55957, x55961);
  nand n55966(x55966, x55503, x55513);
  nand n55969(x55969, x55968, x55967);
  nand n55970(x55970, x55969, x55966);
  nand n55972(x55972, x55522, x55971);
  nand n55974(x55974, x55973, x55970);
  nand n55975(x55975, x55974, x55972);
  nand n55977(x55977, x55966, x55972);
  nand n55978(x55978, x55532, x55542);
  nand n55979(x55979, x55531, x55541);
  nand n55980(x55980, x55979, x55978);
  nand n55982(x55982, x55551, x55981);
  nand n55983(x55983, x55550, x55980);
  nand n55984(x55984, x55983, x55982);
  nand n55986(x55986, x55978, x55982);
  nand n55987(x55987, x55533, x55543);
  nand n55990(x55990, x55989, x55988);
  nand n55991(x55991, x55990, x55987);
  nand n55993(x55993, x55552, x55992);
  nand n55995(x55995, x55994, x55991);
  nand n55996(x55996, x55995, x55993);
  nand n55998(x55998, x55563, x55573);
  nand n55999(x55999, x55562, x55572);
  nand n56000(x56000, x55999, x55998);
  nand n56002(x56002, x55581, x56001);
  nand n56003(x56003, x55580, x56000);
  nand n56004(x56004, x56003, x56002);
  nand n56006(x56006, x85794, x85830);
  nand n56007(x56007, x55035, x55582);
  nand n56008(x56008, x56007, x56006);
  nand n56009(x56009, x85796, x85832);
  nand n56010(x56010, x55039, x55585);
  nand n56011(x56011, x56010, x56009);
  nand n56013(x56013, x55594, x85834);
  nand n56014(x56014, x55593, x55588);
  nand n56015(x56015, x56014, x56013);
  nand n56017(x56017, x85799, x85801);
  nand n56018(x56018, x55591, x55595);
  nand n56019(x56019, x56018, x56017);
  nand n56021(x56021, x55602, x56020);
  nand n56022(x56022, x55601, x56019);
  nand n56023(x56023, x56022, x56021);
  nand n56025(x56025, x56017, x56021);
  nand n56026(x56026, x85803, x85805);
  nand n56027(x56027, x55598, x55603);
  nand n56028(x56028, x56027, x56026);
  nand n56030(x56030, x55610, x56029);
  nand n56031(x56031, x55609, x56028);
  nand n56032(x56032, x56031, x56030);
  nand n56034(x56034, x56026, x56030);
  nand n56035(x56035, x85807, x85809);
  nand n56036(x56036, x55606, x55611);
  nand n56037(x56037, x56036, x56035);
  nand n56039(x56039, x55618, x56038);
  nand n56040(x56040, x55617, x56037);
  nand n56041(x56041, x56040, x56039);
  nand n56043(x56043, x56035, x56039);
  nand n56044(x56044, x85811, x85813);
  nand n56045(x56045, x55614, x55619);
  nand n56046(x56046, x56045, x56044);
  nand n56048(x56048, x55626, x56047);
  nand n56049(x56049, x55625, x56046);
  nand n56050(x56050, x56049, x56048);
  nand n56052(x56052, x56044, x56048);
  nand n56053(x56053, x85815, x85817);
  nand n56054(x56054, x55622, x55627);
  nand n56055(x56055, x56054, x56053);
  nand n56057(x56057, x55634, x56056);
  nand n56058(x56058, x55633, x56055);
  nand n56059(x56059, x56058, x56057);
  nand n56061(x56061, x56053, x56057);
  nand n56062(x56062, x55642, x85676);
  nand n56063(x56063, x55641, x51114);
  nand n56064(x56064, x56063, x56062);
  nand n56067(x56067, x85819, x55643);
  nand n56069(x56069, x55630, x56068);
  nand n56070(x56070, x56069, x56067);
  nand n56072(x56072, x55648, x56071);
  nand n56073(x56073, x55647, x56070);
  nand n56074(x56074, x56073, x56072);
  nand n56076(x56076, x56067, x56072);
  nand n56077(x56077, x55656, x85679);
  nand n56078(x56078, x55655, x52254);
  nand n56079(x56079, x56078, x56077);
  nand n56082(x56082, x85821, x55657);
  nand n56084(x56084, x55644, x56083);
  nand n56085(x56085, x56084, x56082);
  nand n56087(x56087, x55662, x56086);
  nand n56088(x56088, x55661, x56085);
  nand n56089(x56089, x56088, x56087);
  nand n56091(x56091, x56082, x56087);
  nand n56092(x56092, x55670, x85682);
  nand n56093(x56093, x55669, x52296);
  nand n56094(x56094, x56093, x56092);
  nand n56097(x56097, x85823, x55671);
  nand n56099(x56099, x55658, x56098);
  nand n56100(x56100, x56099, x56097);
  nand n56102(x56102, x55676, x56101);
  nand n56103(x56103, x55675, x56100);
  nand n56104(x56104, x56103, x56102);
  nand n56106(x56106, x56097, x56102);
  nand n56107(x56107, x55684, x85687);
  nand n56108(x56108, x55683, x53650);
  nand n56109(x56109, x56108, x56107);
  nand n56112(x56112, x85825, x55685);
  nand n56114(x56114, x55672, x56113);
  nand n56115(x56115, x56114, x56112);
  nand n56117(x56117, x55690, x56116);
  nand n56118(x56118, x55689, x56115);
  nand n56119(x56119, x56118, x56117);
  nand n56121(x56121, x56112, x56117);
  nand n56122(x56122, x55698, x85694);
  nand n56123(x56123, x55697, x53678);
  nand n56124(x56124, x56123, x56122);
  nand n56127(x56127, x85827, x55699);
  nand n56129(x56129, x55686, x56128);
  nand n56130(x56130, x56129, x56127);
  nand n56132(x56132, x55708, x56131);
  nand n56133(x56133, x55707, x56130);
  nand n56134(x56134, x56133, x56132);
  nand n56136(x56136, x56127, x56132);
  nand n56137(x56137, x55717, x85701);
  nand n56138(x56138, x55716, x53712);
  nand n56139(x56139, x56138, x56137);
  nand n56142(x56142, x55709, x55718);
  nand n56145(x56145, x56144, x56143);
  nand n56146(x56146, x56145, x56142);
  nand n56148(x56148, x55728, x56147);
  nand n56149(x56149, x55727, x56146);
  nand n56150(x56150, x56149, x56148);
  nand n56152(x56152, x56142, x56148);
  nand n56153(x56153, x55737, x85708);
  nand n56154(x56154, x55736, x53751);
  nand n56155(x56155, x56154, x56153);
  nand n56158(x56158, x55729, x55738);
  nand n56161(x56161, x56160, x56159);
  nand n56162(x56162, x56161, x56158);
  nand n56164(x56164, x55748, x56163);
  nand n56165(x56165, x55747, x56162);
  nand n56166(x56166, x56165, x56164);
  nand n56168(x56168, x56158, x56164);
  nand n56169(x56169, x55757, x85715);
  nand n56170(x56170, x55756, x53791);
  nand n56171(x56171, x56170, x56169);
  nand n56174(x56174, x55749, x55758);
  nand n56177(x56177, x56176, x56175);
  nand n56178(x56178, x56177, x56174);
  nand n56180(x56180, x55768, x56179);
  nand n56181(x56181, x55767, x56178);
  nand n56182(x56182, x56181, x56180);
  nand n56184(x56184, x56174, x56180);
  nand n56185(x56185, x55777, x85721);
  nand n56186(x56186, x55776, x53831);
  nand n56187(x56187, x56186, x56185);
  nand n56190(x56190, x55769, x55778);
  nand n56193(x56193, x56192, x56191);
  nand n56194(x56194, x56193, x56190);
  nand n56196(x56196, x55788, x56195);
  nand n56197(x56197, x55787, x56194);
  nand n56198(x56198, x56197, x56196);
  nand n56200(x56200, x56190, x56196);
  nand n56201(x56201, x55797, x85727);
  nand n56202(x56202, x55796, x54649);
  nand n56203(x56203, x56202, x56201);
  nand n56206(x56206, x55789, x55798);
  nand n56209(x56209, x56208, x56207);
  nand n56210(x56210, x56209, x56206);
  nand n56212(x56212, x55808, x56211);
  nand n56213(x56213, x55807, x56210);
  nand n56214(x56214, x56213, x56212);
  nand n56216(x56216, x56206, x56212);
  nand n56217(x56217, x55817, x85734);
  nand n56218(x56218, x55816, x54676);
  nand n56219(x56219, x56218, x56217);
  nand n56222(x56222, x55809, x55818);
  nand n56225(x56225, x56224, x56223);
  nand n56226(x56226, x56225, x56222);
  nand n56228(x56228, x55829, x56227);
  nand n56229(x56229, x55828, x56226);
  nand n56230(x56230, x56229, x56228);
  nand n56232(x56232, x56222, x56228);
  nand n56233(x56233, x55838, x85741);
  nand n56234(x56234, x55837, x54703);
  nand n56235(x56235, x56234, x56233);
  nand n56238(x56238, x55830, x55839);
  nand n56241(x56241, x56240, x56239);
  nand n56242(x56242, x56241, x56238);
  nand n56244(x56244, x55850, x56243);
  nand n56245(x56245, x55849, x56242);
  nand n56246(x56246, x56245, x56244);
  nand n56248(x56248, x56238, x56244);
  nand n56249(x56249, x55859, x85746);
  nand n56250(x56250, x55858, x54736);
  nand n56251(x56251, x56250, x56249);
  nand n56254(x56254, x55851, x55860);
  nand n56257(x56257, x56256, x56255);
  nand n56258(x56258, x56257, x56254);
  nand n56260(x56260, x55871, x56259);
  nand n56261(x56261, x55870, x56258);
  nand n56262(x56262, x56261, x56260);
  nand n56264(x56264, x56254, x56260);
  nand n56265(x56265, x55880, x85749);
  nand n56266(x56266, x55879, x54774);
  nand n56267(x56267, x56266, x56265);
  nand n56270(x56270, x55872, x55881);
  nand n56273(x56273, x56272, x56271);
  nand n56274(x56274, x56273, x56270);
  nand n56276(x56276, x55892, x56275);
  nand n56277(x56277, x55891, x56274);
  nand n56278(x56278, x56277, x56276);
  nand n56280(x56280, x56270, x56276);
  nand n56281(x56281, x55901, x85752);
  nand n56282(x56282, x55900, x54812);
  nand n56283(x56283, x56282, x56281);
  nand n56286(x56286, x55893, x55902);
  nand n56289(x56289, x56288, x56287);
  nand n56290(x56290, x56289, x56286);
  nand n56292(x56292, x55913, x56291);
  nand n56293(x56293, x55912, x56290);
  nand n56294(x56294, x56293, x56292);
  nand n56296(x56296, x56286, x56292);
  nand n56297(x56297, x55922, x85755);
  nand n56298(x56298, x55921, x54851);
  nand n56299(x56299, x56298, x56297);
  nand n56302(x56302, x55914, x55923);
  nand n56305(x56305, x56304, x56303);
  nand n56306(x56306, x56305, x56302);
  nand n56308(x56308, x55934, x56307);
  nand n56309(x56309, x55933, x56306);
  nand n56310(x56310, x56309, x56308);
  nand n56312(x56312, x56302, x56308);
  nand n56313(x56313, x55943, x85758);
  nand n56314(x56314, x55942, x54891);
  nand n56315(x56315, x56314, x56313);
  nand n56318(x56318, x55935, x55944);
  nand n56321(x56321, x56320, x56319);
  nand n56322(x56322, x56321, x56318);
  nand n56324(x56324, x55955, x56323);
  nand n56325(x56325, x55954, x56322);
  nand n56326(x56326, x56325, x56324);
  nand n56328(x56328, x56318, x56324);
  nand n56329(x56329, x55964, x85761);
  nand n56330(x56330, x55963, x54931);
  nand n56331(x56331, x56330, x56329);
  nand n56334(x56334, x55956, x55965);
  nand n56337(x56337, x56336, x56335);
  nand n56338(x56338, x56337, x56334);
  nand n56340(x56340, x55976, x56339);
  nand n56341(x56341, x55975, x56338);
  nand n56342(x56342, x56341, x56340);
  nand n56344(x56344, x56334, x56340);
  nand n56345(x56345, x55985, x54981);
  nand n56346(x56346, x55984, x54980);
  nand n56347(x56347, x56346, x56345);
  nand n56350(x56350, x55977, x55986);
  nand n56353(x56353, x56352, x56351);
  nand n56354(x56354, x56353, x56350);
  nand n56356(x56356, x55997, x56355);
  nand n56357(x56357, x55996, x56354);
  nand n56358(x56358, x56357, x56356);
  nand n56360(x56360, x56005, x55028);
  nand n56361(x56361, x56004, x55027);
  nand n56362(x56362, x56361, x56360);
  nand n56364(x56364, x85828, x85840);
  nand n56365(x56365, x55034, x55029);
  nand n56366(x56366, x56365, x56364);
  nand n56367(x56367, x56012, x85843);
  nand n56368(x56368, x56011, x56006);
  nand n56369(x56369, x56368, x56367);
  nand n56370(x56370, x56016, x85845);
  nand n56371(x56371, x56015, x56009);
  nand n56372(x56372, x56371, x56370);
  nand n56374(x56374, x56024, x85847);
  nand n56375(x56375, x56023, x56013);
  nand n56376(x56376, x56375, x56374);
  nand n56379(x56379, x56033, x56025);
  nand n56380(x56380, x56032, x56378);
  nand n56381(x56381, x56380, x56379);
  nand n56384(x56384, x56042, x56034);
  nand n56385(x56385, x56041, x56383);
  nand n56386(x56386, x56385, x56384);
  nand n56389(x56389, x56051, x56043);
  nand n56390(x56390, x56050, x56388);
  nand n56391(x56391, x56390, x56389);
  nand n56394(x56394, x56060, x56052);
  nand n56395(x56395, x56059, x56393);
  nand n56396(x56396, x56395, x56394);
  nand n56398(x56398, x56061, x56066);
  nand n56400(x56400, x56399, x56062);
  nand n56401(x56401, x56400, x56398);
  nand n56403(x56403, x56075, x56402);
  nand n56404(x56404, x56074, x56401);
  nand n56405(x56405, x56404, x56403);
  nand n56407(x56407, x56398, x56403);
  nand n56408(x56408, x56076, x56081);
  nand n56410(x56410, x56409, x56077);
  nand n56411(x56411, x56410, x56408);
  nand n56413(x56413, x56090, x56412);
  nand n56414(x56414, x56089, x56411);
  nand n56415(x56415, x56414, x56413);
  nand n56417(x56417, x56408, x56413);
  nand n56418(x56418, x56091, x56096);
  nand n56420(x56420, x56419, x56092);
  nand n56421(x56421, x56420, x56418);
  nand n56423(x56423, x56105, x56422);
  nand n56424(x56424, x56104, x56421);
  nand n56425(x56425, x56424, x56423);
  nand n56427(x56427, x56418, x56423);
  nand n56428(x56428, x56106, x56111);
  nand n56430(x56430, x56429, x56107);
  nand n56431(x56431, x56430, x56428);
  nand n56433(x56433, x56120, x56432);
  nand n56434(x56434, x56119, x56431);
  nand n56435(x56435, x56434, x56433);
  nand n56437(x56437, x56428, x56433);
  nand n56438(x56438, x56121, x56126);
  nand n56440(x56440, x56439, x56122);
  nand n56441(x56441, x56440, x56438);
  nand n56443(x56443, x56135, x56442);
  nand n56444(x56444, x56134, x56441);
  nand n56445(x56445, x56444, x56443);
  nand n56447(x56447, x56438, x56443);
  nand n56448(x56448, x56136, x56141);
  nand n56450(x56450, x56449, x56137);
  nand n56451(x56451, x56450, x56448);
  nand n56453(x56453, x56151, x56452);
  nand n56454(x56454, x56150, x56451);
  nand n56455(x56455, x56454, x56453);
  nand n56457(x56457, x56448, x56453);
  nand n56458(x56458, x56152, x56157);
  nand n56460(x56460, x56459, x56153);
  nand n56461(x56461, x56460, x56458);
  nand n56463(x56463, x56167, x56462);
  nand n56464(x56464, x56166, x56461);
  nand n56465(x56465, x56464, x56463);
  nand n56467(x56467, x56458, x56463);
  nand n56468(x56468, x56168, x56173);
  nand n56470(x56470, x56469, x56169);
  nand n56471(x56471, x56470, x56468);
  nand n56473(x56473, x56183, x56472);
  nand n56474(x56474, x56182, x56471);
  nand n56475(x56475, x56474, x56473);
  nand n56477(x56477, x56468, x56473);
  nand n56478(x56478, x56184, x56189);
  nand n56480(x56480, x56479, x56185);
  nand n56481(x56481, x56480, x56478);
  nand n56483(x56483, x56199, x56482);
  nand n56484(x56484, x56198, x56481);
  nand n56485(x56485, x56484, x56483);
  nand n56487(x56487, x56478, x56483);
  nand n56488(x56488, x56200, x56205);
  nand n56490(x56490, x56489, x56201);
  nand n56491(x56491, x56490, x56488);
  nand n56493(x56493, x56215, x56492);
  nand n56494(x56494, x56214, x56491);
  nand n56495(x56495, x56494, x56493);
  nand n56497(x56497, x56488, x56493);
  nand n56498(x56498, x56216, x56221);
  nand n56500(x56500, x56499, x56217);
  nand n56501(x56501, x56500, x56498);
  nand n56503(x56503, x56231, x56502);
  nand n56504(x56504, x56230, x56501);
  nand n56505(x56505, x56504, x56503);
  nand n56507(x56507, x56498, x56503);
  nand n56508(x56508, x56232, x56237);
  nand n56510(x56510, x56509, x56233);
  nand n56511(x56511, x56510, x56508);
  nand n56513(x56513, x56247, x56512);
  nand n56514(x56514, x56246, x56511);
  nand n56515(x56515, x56514, x56513);
  nand n56517(x56517, x56508, x56513);
  nand n56518(x56518, x56248, x56253);
  nand n56520(x56520, x56519, x56249);
  nand n56521(x56521, x56520, x56518);
  nand n56523(x56523, x56263, x56522);
  nand n56524(x56524, x56262, x56521);
  nand n56525(x56525, x56524, x56523);
  nand n56527(x56527, x56518, x56523);
  nand n56528(x56528, x56264, x56269);
  nand n56530(x56530, x56529, x56265);
  nand n56531(x56531, x56530, x56528);
  nand n56533(x56533, x56279, x56532);
  nand n56534(x56534, x56278, x56531);
  nand n56535(x56535, x56534, x56533);
  nand n56537(x56537, x56528, x56533);
  nand n56538(x56538, x56280, x56285);
  nand n56540(x56540, x56539, x56281);
  nand n56541(x56541, x56540, x56538);
  nand n56543(x56543, x56295, x56542);
  nand n56544(x56544, x56294, x56541);
  nand n56545(x56545, x56544, x56543);
  nand n56547(x56547, x56538, x56543);
  nand n56548(x56548, x56296, x56301);
  nand n56550(x56550, x56549, x56297);
  nand n56551(x56551, x56550, x56548);
  nand n56553(x56553, x56311, x56552);
  nand n56554(x56554, x56310, x56551);
  nand n56555(x56555, x56554, x56553);
  nand n56557(x56557, x56548, x56553);
  nand n56558(x56558, x56312, x56317);
  nand n56560(x56560, x56559, x56313);
  nand n56561(x56561, x56560, x56558);
  nand n56563(x56563, x56327, x56562);
  nand n56564(x56564, x56326, x56561);
  nand n56565(x56565, x56564, x56563);
  nand n56567(x56567, x56558, x56563);
  nand n56568(x56568, x56328, x56333);
  nand n56570(x56570, x56569, x56329);
  nand n56571(x56571, x56570, x56568);
  nand n56573(x56573, x56343, x56572);
  nand n56574(x56574, x56342, x56571);
  nand n56575(x56575, x56574, x56573);
  nand n56577(x56577, x56568, x56573);
  nand n56578(x56578, x56344, x56349);
  nand n56580(x56580, x56579, x56345);
  nand n56581(x56581, x56580, x56578);
  nand n56583(x56583, x56359, x56582);
  nand n56584(x56584, x56358, x56581);
  nand n56585(x56585, x56584, x56583);
  nand n56587(x56587, x85841, x85842);
  nand n56588(x56588, x56364, x55032);
  nand n56589(x56589, x56588, x56587);
  nand n56591(x56591, x85829, x56590);
  nand n56592(x56592, x55584, x56589);
  nand n56593(x56593, x56592, x56591);
  nand n56594(x56594, x56587, x56591);
  nand n56595(x56595, x85831, x85853);
  nand n56596(x56596, x55587, x56008);
  nand n56597(x56597, x56596, x56595);
  nand n56599(x56599, x85833, x85855);
  nand n56600(x56600, x55590, x56369);
  nand n56601(x56601, x56600, x56599);
  nand n56603(x56603, x85844, x56373);
  nand n56604(x56604, x56367, x56372);
  nand n56605(x56605, x56604, x56603);
  nand n56607(x56607, x85835, x56606);
  nand n56608(x56608, x55597, x56605);
  nand n56609(x56609, x56608, x56607);
  nand n56611(x56611, x56603, x56607);
  nand n56612(x56612, x85846, x56377);
  nand n56613(x56613, x56370, x56376);
  nand n56614(x56614, x56613, x56612);
  nand n56616(x56616, x85836, x56615);
  nand n56617(x56617, x55605, x56614);
  nand n56618(x56618, x56617, x56616);
  nand n56620(x56620, x56612, x56616);
  nand n56621(x56621, x85848, x56382);
  nand n56622(x56622, x56374, x56381);
  nand n56623(x56623, x56622, x56621);
  nand n56625(x56625, x85837, x56624);
  nand n56626(x56626, x55613, x56623);
  nand n56627(x56627, x56626, x56625);
  nand n56629(x56629, x56621, x56625);
  nand n56630(x56630, x85849, x56387);
  nand n56631(x56631, x56379, x56386);
  nand n56632(x56632, x56631, x56630);
  nand n56634(x56634, x85838, x56633);
  nand n56635(x56635, x55621, x56632);
  nand n56636(x56636, x56635, x56634);
  nand n56638(x56638, x56630, x56634);
  nand n56639(x56639, x85850, x56392);
  nand n56640(x56640, x56384, x56391);
  nand n56641(x56641, x56640, x56639);
  nand n56643(x56643, x85839, x56642);
  nand n56644(x56644, x55629, x56641);
  nand n56645(x56645, x56644, x56643);
  nand n56647(x56647, x56639, x56643);
  nand n56648(x56648, x85851, x56397);
  nand n56649(x56649, x56389, x56396);
  nand n56650(x56650, x56649, x56648);
  nand n56652(x56652, x56065, x56651);
  nand n56653(x56653, x56064, x56650);
  nand n56654(x56654, x56653, x56652);
  nand n56656(x56656, x56648, x56652);
  nand n56657(x56657, x85852, x56406);
  nand n56658(x56658, x56394, x56405);
  nand n56659(x56659, x56658, x56657);
  nand n56661(x56661, x56080, x56660);
  nand n56662(x56662, x56079, x56659);
  nand n56663(x56663, x56662, x56661);
  nand n56665(x56665, x56657, x56661);
  nand n56666(x56666, x56407, x56416);
  nand n56668(x56668, x56667, x56415);
  nand n56669(x56669, x56668, x56666);
  nand n56671(x56671, x56095, x56670);
  nand n56672(x56672, x56094, x56669);
  nand n56673(x56673, x56672, x56671);
  nand n56675(x56675, x56666, x56671);
  nand n56676(x56676, x56417, x56426);
  nand n56678(x56678, x56677, x56425);
  nand n56679(x56679, x56678, x56676);
  nand n56681(x56681, x56110, x56680);
  nand n56682(x56682, x56109, x56679);
  nand n56683(x56683, x56682, x56681);
  nand n56685(x56685, x56676, x56681);
  nand n56686(x56686, x56427, x56436);
  nand n56688(x56688, x56687, x56435);
  nand n56689(x56689, x56688, x56686);
  nand n56691(x56691, x56125, x56690);
  nand n56692(x56692, x56124, x56689);
  nand n56693(x56693, x56692, x56691);
  nand n56695(x56695, x56686, x56691);
  nand n56696(x56696, x56437, x56446);
  nand n56698(x56698, x56697, x56445);
  nand n56699(x56699, x56698, x56696);
  nand n56701(x56701, x56140, x56700);
  nand n56702(x56702, x56139, x56699);
  nand n56703(x56703, x56702, x56701);
  nand n56705(x56705, x56696, x56701);
  nand n56706(x56706, x56447, x56456);
  nand n56708(x56708, x56707, x56455);
  nand n56709(x56709, x56708, x56706);
  nand n56711(x56711, x56156, x56710);
  nand n56712(x56712, x56155, x56709);
  nand n56713(x56713, x56712, x56711);
  nand n56715(x56715, x56706, x56711);
  nand n56716(x56716, x56457, x56466);
  nand n56718(x56718, x56717, x56465);
  nand n56719(x56719, x56718, x56716);
  nand n56721(x56721, x56172, x56720);
  nand n56722(x56722, x56171, x56719);
  nand n56723(x56723, x56722, x56721);
  nand n56725(x56725, x56716, x56721);
  nand n56726(x56726, x56467, x56476);
  nand n56728(x56728, x56727, x56475);
  nand n56729(x56729, x56728, x56726);
  nand n56731(x56731, x56188, x56730);
  nand n56732(x56732, x56187, x56729);
  nand n56733(x56733, x56732, x56731);
  nand n56735(x56735, x56726, x56731);
  nand n56736(x56736, x56477, x56486);
  nand n56738(x56738, x56737, x56485);
  nand n56739(x56739, x56738, x56736);
  nand n56741(x56741, x56204, x56740);
  nand n56742(x56742, x56203, x56739);
  nand n56743(x56743, x56742, x56741);
  nand n56745(x56745, x56736, x56741);
  nand n56746(x56746, x56487, x56496);
  nand n56748(x56748, x56747, x56495);
  nand n56749(x56749, x56748, x56746);
  nand n56751(x56751, x56220, x56750);
  nand n56752(x56752, x56219, x56749);
  nand n56753(x56753, x56752, x56751);
  nand n56755(x56755, x56746, x56751);
  nand n56756(x56756, x56497, x56506);
  nand n56758(x56758, x56757, x56505);
  nand n56759(x56759, x56758, x56756);
  nand n56761(x56761, x56236, x56760);
  nand n56762(x56762, x56235, x56759);
  nand n56763(x56763, x56762, x56761);
  nand n56765(x56765, x56756, x56761);
  nand n56766(x56766, x56507, x56516);
  nand n56768(x56768, x56767, x56515);
  nand n56769(x56769, x56768, x56766);
  nand n56771(x56771, x56252, x56770);
  nand n56772(x56772, x56251, x56769);
  nand n56773(x56773, x56772, x56771);
  nand n56775(x56775, x56766, x56771);
  nand n56776(x56776, x56517, x56526);
  nand n56778(x56778, x56777, x56525);
  nand n56779(x56779, x56778, x56776);
  nand n56781(x56781, x56268, x56780);
  nand n56782(x56782, x56267, x56779);
  nand n56783(x56783, x56782, x56781);
  nand n56785(x56785, x56776, x56781);
  nand n56786(x56786, x56527, x56536);
  nand n56788(x56788, x56787, x56535);
  nand n56789(x56789, x56788, x56786);
  nand n56791(x56791, x56284, x56790);
  nand n56792(x56792, x56283, x56789);
  nand n56793(x56793, x56792, x56791);
  nand n56795(x56795, x56786, x56791);
  nand n56796(x56796, x56537, x56546);
  nand n56798(x56798, x56797, x56545);
  nand n56799(x56799, x56798, x56796);
  nand n56801(x56801, x56300, x56800);
  nand n56802(x56802, x56299, x56799);
  nand n56803(x56803, x56802, x56801);
  nand n56805(x56805, x56796, x56801);
  nand n56806(x56806, x56547, x56556);
  nand n56808(x56808, x56807, x56555);
  nand n56809(x56809, x56808, x56806);
  nand n56811(x56811, x56316, x56810);
  nand n56812(x56812, x56315, x56809);
  nand n56813(x56813, x56812, x56811);
  nand n56815(x56815, x56806, x56811);
  nand n56816(x56816, x56557, x56566);
  nand n56818(x56818, x56817, x56565);
  nand n56819(x56819, x56818, x56816);
  nand n56821(x56821, x56332, x56820);
  nand n56822(x56822, x56331, x56819);
  nand n56823(x56823, x56822, x56821);
  nand n56825(x56825, x56816, x56821);
  nand n56826(x56826, x56567, x56576);
  nand n56828(x56828, x56827, x56575);
  nand n56829(x56829, x56828, x56826);
  nand n56831(x56831, x56348, x56830);
  nand n56832(x56832, x56347, x56829);
  nand n56833(x56833, x56832, x56831);
  nand n56835(x56835, x56826, x56831);
  nand n56836(x56836, x56577, x56586);
  nand n56838(x56838, x56837, x56585);
  nand n56839(x56839, x56838, x56836);
  nand n56841(x56841, x56363, x56840);
  nand n56842(x56842, x56362, x56839);
  nand n56843(x56843, x56842, x56841);
  nand n56845(x56845, x56594, x56598);
  nand n56847(x56847, x56846, x56597);
  nand n56848(x56848, x56847, x56845);
  nand n56849(x56849, x85854, x56602);
  nand n56850(x56850, x56595, x56601);
  nand n56851(x56851, x56850, x56849);
  nand n56853(x56853, x85856, x56610);
  nand n56854(x56854, x56599, x56609);
  nand n56855(x56855, x56854, x56853);
  nand n56857(x56857, x56611, x56619);
  nand n56859(x56859, x56858, x56618);
  nand n56860(x56860, x56859, x56857);
  nand n56862(x56862, x56620, x56628);
  nand n56864(x56864, x56863, x56627);
  nand n56865(x56865, x56864, x56862);
  nand n56867(x56867, x56629, x56637);
  nand n56869(x56869, x56868, x56636);
  nand n56870(x56870, x56869, x56867);
  nand n56872(x56872, x56638, x56646);
  nand n56874(x56874, x56873, x56645);
  nand n56875(x56875, x56874, x56872);
  nand n56877(x56877, x56647, x56655);
  nand n56879(x56879, x56878, x56654);
  nand n56880(x56880, x56879, x56877);
  nand n56882(x56882, x56656, x56664);
  nand n56884(x56884, x56883, x56663);
  nand n56885(x56885, x56884, x56882);
  nand n56887(x56887, x56665, x56674);
  nand n56889(x56889, x56888, x56673);
  nand n56890(x56890, x56889, x56887);
  nand n56892(x56892, x56675, x56684);
  nand n56894(x56894, x56893, x56683);
  nand n56895(x56895, x56894, x56892);
  nand n56897(x56897, x56685, x56694);
  nand n56899(x56899, x56898, x56693);
  nand n56900(x56900, x56899, x56897);
  nand n56902(x56902, x56695, x56704);
  nand n56904(x56904, x56903, x56703);
  nand n56905(x56905, x56904, x56902);
  nand n56907(x56907, x56705, x56714);
  nand n56909(x56909, x56908, x56713);
  nand n56910(x56910, x56909, x56907);
  nand n56912(x56912, x56715, x56724);
  nand n56914(x56914, x56913, x56723);
  nand n56915(x56915, x56914, x56912);
  nand n56917(x56917, x56725, x56734);
  nand n56919(x56919, x56918, x56733);
  nand n56920(x56920, x56919, x56917);
  nand n56922(x56922, x56735, x56744);
  nand n56924(x56924, x56923, x56743);
  nand n56925(x56925, x56924, x56922);
  nand n56927(x56927, x56745, x56754);
  nand n56929(x56929, x56928, x56753);
  nand n56930(x56930, x56929, x56927);
  nand n56932(x56932, x56755, x56764);
  nand n56934(x56934, x56933, x56763);
  nand n56935(x56935, x56934, x56932);
  nand n56937(x56937, x56765, x56774);
  nand n56939(x56939, x56938, x56773);
  nand n56940(x56940, x56939, x56937);
  nand n56942(x56942, x56775, x56784);
  nand n56944(x56944, x56943, x56783);
  nand n56945(x56945, x56944, x56942);
  nand n56947(x56947, x56785, x56794);
  nand n56949(x56949, x56948, x56793);
  nand n56950(x56950, x56949, x56947);
  nand n56952(x56952, x56795, x56804);
  nand n56954(x56954, x56953, x56803);
  nand n56955(x56955, x56954, x56952);
  nand n56957(x56957, x56805, x56814);
  nand n56959(x56959, x56958, x56813);
  nand n56960(x56960, x56959, x56957);
  nand n56962(x56962, x56815, x56824);
  nand n56964(x56964, x56963, x56823);
  nand n56965(x56965, x56964, x56962);
  nand n56967(x56967, x56825, x56834);
  nand n56969(x56969, x56968, x56833);
  nand n56970(x56970, x56969, x56967);
  nand n56972(x56972, x56835, x56844);
  nand n56974(x56974, x56973, x56843);
  nand n56975(x56975, x56974, x56972);
  nand n57002(x57002, x56852, x56977);
  nand n57003(x57003, x57002, x56849);
  nand n57004(x57004, x56856, x56978);
  nand n57005(x57005, x57004, x56853);
  nand n57006(x57006, x56856, x56852);
  nand n57008(x57008, x56861, x56979);
  nand n57009(x57009, x57008, x56857);
  nand n57010(x57010, x56861, x56856);
  nand n57012(x57012, x56866, x56980);
  nand n57013(x57013, x57012, x56862);
  nand n57014(x57014, x56866, x56861);
  nand n57016(x57016, x56871, x56981);
  nand n57017(x57017, x57016, x56867);
  nand n57018(x57018, x56871, x56866);
  nand n57020(x57020, x56876, x56982);
  nand n57021(x57021, x57020, x56872);
  nand n57022(x57022, x56876, x56871);
  nand n57024(x57024, x56881, x56983);
  nand n57025(x57025, x57024, x56877);
  nand n57026(x57026, x56881, x56876);
  nand n57028(x57028, x56886, x56984);
  nand n57029(x57029, x57028, x56882);
  nand n57030(x57030, x56886, x56881);
  nand n57032(x57032, x56891, x56985);
  nand n57033(x57033, x57032, x56887);
  nand n57034(x57034, x56891, x56886);
  nand n57036(x57036, x56896, x56986);
  nand n57037(x57037, x57036, x56892);
  nand n57038(x57038, x56896, x56891);
  nand n57040(x57040, x56901, x56987);
  nand n57041(x57041, x57040, x56897);
  nand n57042(x57042, x56901, x56896);
  nand n57044(x57044, x56906, x56988);
  nand n57045(x57045, x57044, x56902);
  nand n57046(x57046, x56906, x56901);
  nand n57048(x57048, x56911, x56989);
  nand n57049(x57049, x57048, x56907);
  nand n57050(x57050, x56911, x56906);
  nand n57052(x57052, x56916, x56990);
  nand n57053(x57053, x57052, x56912);
  nand n57054(x57054, x56916, x56911);
  nand n57056(x57056, x56921, x56991);
  nand n57057(x57057, x57056, x56917);
  nand n57058(x57058, x56921, x56916);
  nand n57060(x57060, x56926, x56992);
  nand n57061(x57061, x57060, x56922);
  nand n57062(x57062, x56926, x56921);
  nand n57064(x57064, x56931, x56993);
  nand n57065(x57065, x57064, x56927);
  nand n57066(x57066, x56931, x56926);
  nand n57068(x57068, x56936, x56994);
  nand n57069(x57069, x57068, x56932);
  nand n57070(x57070, x56936, x56931);
  nand n57072(x57072, x56941, x56995);
  nand n57073(x57073, x57072, x56937);
  nand n57074(x57074, x56941, x56936);
  nand n57076(x57076, x56946, x56996);
  nand n57077(x57077, x57076, x56942);
  nand n57078(x57078, x56946, x56941);
  nand n57080(x57080, x56951, x56997);
  nand n57081(x57081, x57080, x56947);
  nand n57082(x57082, x56951, x56946);
  nand n57084(x57084, x56956, x56998);
  nand n57085(x57085, x57084, x56952);
  nand n57086(x57086, x56956, x56951);
  nand n57088(x57088, x56961, x56999);
  nand n57089(x57089, x57088, x56957);
  nand n57090(x57090, x56961, x56956);
  nand n57092(x57092, x56966, x57000);
  nand n57093(x57093, x57092, x56962);
  nand n57094(x57094, x56966, x56961);
  nand n57096(x57096, x56971, x57001);
  nand n57097(x57097, x57096, x56967);
  nand n57098(x57098, x56971, x56966);
  nand n57101(x57101, x57007, x56977);
  nand n57103(x57103, x57101, x57102);
  nand n57104(x57104, x57011, x57003);
  nand n57106(x57106, x57104, x57105);
  nand n57107(x57107, x57015, x57005);
  nand n57109(x57109, x57107, x57108);
  nand n57110(x57110, x57015, x57007);
  nand n57112(x57112, x57019, x57009);
  nand n57114(x57114, x57112, x57113);
  nand n57115(x57115, x57019, x57011);
  nand n57117(x57117, x57023, x57013);
  nand n57119(x57119, x57117, x57118);
  nand n57120(x57120, x57023, x57015);
  nand n57122(x57122, x57027, x57017);
  nand n57124(x57124, x57122, x57123);
  nand n57125(x57125, x57027, x57019);
  nand n57127(x57127, x57031, x57021);
  nand n57129(x57129, x57127, x57128);
  nand n57130(x57130, x57031, x57023);
  nand n57132(x57132, x57035, x57025);
  nand n57134(x57134, x57132, x57133);
  nand n57135(x57135, x57035, x57027);
  nand n57137(x57137, x57039, x57029);
  nand n57139(x57139, x57137, x57138);
  nand n57140(x57140, x57039, x57031);
  nand n57142(x57142, x57043, x57033);
  nand n57144(x57144, x57142, x57143);
  nand n57145(x57145, x57043, x57035);
  nand n57147(x57147, x57047, x57037);
  nand n57149(x57149, x57147, x57148);
  nand n57150(x57150, x57047, x57039);
  nand n57152(x57152, x57051, x57041);
  nand n57154(x57154, x57152, x57153);
  nand n57155(x57155, x57051, x57043);
  nand n57157(x57157, x57055, x57045);
  nand n57159(x57159, x57157, x57158);
  nand n57160(x57160, x57055, x57047);
  nand n57162(x57162, x57059, x57049);
  nand n57164(x57164, x57162, x57163);
  nand n57165(x57165, x57059, x57051);
  nand n57167(x57167, x57063, x57053);
  nand n57169(x57169, x57167, x57168);
  nand n57170(x57170, x57063, x57055);
  nand n57172(x57172, x57067, x57057);
  nand n57174(x57174, x57172, x57173);
  nand n57175(x57175, x57067, x57059);
  nand n57177(x57177, x57071, x57061);
  nand n57179(x57179, x57177, x57178);
  nand n57180(x57180, x57071, x57063);
  nand n57182(x57182, x57075, x57065);
  nand n57184(x57184, x57182, x57183);
  nand n57185(x57185, x57075, x57067);
  nand n57187(x57187, x57079, x57069);
  nand n57189(x57189, x57187, x57188);
  nand n57190(x57190, x57079, x57071);
  nand n57192(x57192, x57083, x57073);
  nand n57194(x57194, x57192, x57193);
  nand n57195(x57195, x57083, x57075);
  nand n57197(x57197, x57087, x57077);
  nand n57199(x57199, x57197, x57198);
  nand n57200(x57200, x57087, x57079);
  nand n57202(x57202, x57091, x57081);
  nand n57204(x57204, x57202, x57203);
  nand n57205(x57205, x57091, x57083);
  nand n57207(x57207, x57095, x57085);
  nand n57209(x57209, x57207, x57208);
  nand n57210(x57210, x57095, x57087);
  nand n57212(x57212, x57099, x57089);
  nand n57214(x57214, x57212, x57213);
  nand n57215(x57215, x57099, x57091);
  nand n57219(x57219, x57111, x56977);
  nand n57221(x57221, x57219, x57220);
  nand n57222(x57222, x57116, x57003);
  nand n57224(x57224, x57222, x57223);
  nand n57225(x57225, x57121, x57103);
  nand n57227(x57227, x57225, x57226);
  nand n57228(x57228, x57126, x57106);
  nand n57230(x57230, x57228, x57229);
  nand n57231(x57231, x57131, x57109);
  nand n57233(x57233, x57231, x57232);
  nand n57234(x57234, x57131, x57111);
  nand n57236(x57236, x57136, x57114);
  nand n57238(x57238, x57236, x57237);
  nand n57239(x57239, x57136, x57116);
  nand n57241(x57241, x57141, x57119);
  nand n57243(x57243, x57241, x57242);
  nand n57244(x57244, x57141, x57121);
  nand n57246(x57246, x57146, x57124);
  nand n57248(x57248, x57246, x57247);
  nand n57249(x57249, x57146, x57126);
  nand n57251(x57251, x57151, x57129);
  nand n57253(x57253, x57251, x57252);
  nand n57254(x57254, x57151, x57131);
  nand n57256(x57256, x57156, x57134);
  nand n57258(x57258, x57256, x57257);
  nand n57259(x57259, x57156, x57136);
  nand n57261(x57261, x57161, x57139);
  nand n57263(x57263, x57261, x57262);
  nand n57264(x57264, x57161, x57141);
  nand n57266(x57266, x57166, x57144);
  nand n57268(x57268, x57266, x57267);
  nand n57269(x57269, x57166, x57146);
  nand n57271(x57271, x57171, x57149);
  nand n57273(x57273, x57271, x57272);
  nand n57274(x57274, x57171, x57151);
  nand n57276(x57276, x57176, x57154);
  nand n57278(x57278, x57276, x57277);
  nand n57279(x57279, x57176, x57156);
  nand n57281(x57281, x57181, x57159);
  nand n57283(x57283, x57281, x57282);
  nand n57284(x57284, x57181, x57161);
  nand n57286(x57286, x57186, x57164);
  nand n57288(x57288, x57286, x57287);
  nand n57289(x57289, x57186, x57166);
  nand n57291(x57291, x57191, x57169);
  nand n57293(x57293, x57291, x57292);
  nand n57294(x57294, x57191, x57171);
  nand n57296(x57296, x57196, x57174);
  nand n57298(x57298, x57296, x57297);
  nand n57299(x57299, x57196, x57176);
  nand n57301(x57301, x57201, x57179);
  nand n57303(x57303, x57301, x57302);
  nand n57304(x57304, x57201, x57181);
  nand n57306(x57306, x57206, x57184);
  nand n57308(x57308, x57306, x57307);
  nand n57309(x57309, x57206, x57186);
  nand n57311(x57311, x57211, x57189);
  nand n57313(x57313, x57311, x57312);
  nand n57314(x57314, x57211, x57191);
  nand n57316(x57316, x57216, x57194);
  nand n57318(x57318, x57316, x57317);
  nand n57319(x57319, x57216, x57196);
  nand n57325(x57325, x57235, x56977);
  nand n57327(x57327, x57325, x57326);
  nand n57328(x57328, x57240, x57003);
  nand n57330(x57330, x57328, x57329);
  nand n57331(x57331, x57245, x57103);
  nand n57333(x57333, x57331, x57332);
  nand n57334(x57334, x57250, x57106);
  nand n57336(x57336, x57334, x57335);
  nand n57337(x57337, x57255, x57221);
  nand n57339(x57339, x57337, x57338);
  nand n57340(x57340, x57260, x57224);
  nand n57342(x57342, x57340, x57341);
  nand n57343(x57343, x57265, x57227);
  nand n57345(x57345, x57343, x57344);
  nand n57346(x57346, x57270, x57230);
  nand n57348(x57348, x57346, x57347);
  nand n57349(x57349, x57275, x57233);
  nand n57351(x57351, x57349, x57350);
  nand n57352(x57352, x57275, x57235);
  nand n57354(x57354, x57280, x57238);
  nand n57356(x57356, x57354, x57355);
  nand n57357(x57357, x57280, x57240);
  nand n57359(x57359, x57285, x57243);
  nand n57361(x57361, x57359, x57360);
  nand n57362(x57362, x57285, x57245);
  nand n57364(x57364, x57290, x57248);
  nand n57366(x57366, x57364, x57365);
  nand n57367(x57367, x57290, x57250);
  nand n57369(x57369, x57295, x57253);
  nand n57371(x57371, x57369, x57370);
  nand n57372(x57372, x57295, x57255);
  nand n57374(x57374, x57300, x57258);
  nand n57376(x57376, x57374, x57375);
  nand n57377(x57377, x57300, x57260);
  nand n57379(x57379, x57305, x57263);
  nand n57381(x57381, x57379, x57380);
  nand n57382(x57382, x57305, x57265);
  nand n57384(x57384, x57310, x57268);
  nand n57386(x57386, x57384, x57385);
  nand n57387(x57387, x57310, x57270);
  nand n57389(x57389, x57315, x57273);
  nand n57391(x57391, x57389, x57390);
  nand n57392(x57392, x57315, x57275);
  nand n57394(x57394, x57320, x57278);
  nand n57396(x57396, x57394, x57395);
  nand n57397(x57397, x57320, x57280);
  nand n57405(x57405, x57353, x56977);
  nand n57407(x57407, x57405, x57406);
  nand n57408(x57408, x57358, x57003);
  nand n57410(x57410, x57408, x57409);
  nand n57411(x57411, x57363, x57103);
  nand n57413(x57413, x57411, x57412);
  nand n57414(x57414, x57368, x57106);
  nand n57416(x57416, x57414, x57415);
  nand n57417(x57417, x57373, x57221);
  nand n57419(x57419, x57417, x57418);
  nand n57420(x57420, x57378, x57224);
  nand n57422(x57422, x57420, x57421);
  nand n57423(x57423, x57383, x57227);
  nand n57425(x57425, x57423, x57424);
  nand n57426(x57426, x57388, x57230);
  nand n57428(x57428, x57426, x57427);
  nand n57429(x57429, x57393, x57327);
  nand n57431(x57431, x57429, x57430);
  nand n57432(x57432, x57398, x57330);
  nand n57434(x57434, x57432, x57433);
  nand n57435(x57435, x56851, x56845);
  nand n57436(x57436, x57435, x57002);
  nand n57438(x57438, x56856, x57003);
  nand n57439(x57439, x56855, x57100);
  nand n57440(x57440, x57439, x57438);
  nand n57442(x57442, x56861, x57103);
  nand n57443(x57443, x56860, x57217);
  nand n57444(x57444, x57443, x57442);
  nand n57446(x57446, x56866, x57106);
  nand n57447(x57447, x56865, x57218);
  nand n57448(x57448, x57447, x57446);
  nand n57450(x57450, x56871, x57221);
  nand n57451(x57451, x56870, x57321);
  nand n57452(x57452, x57451, x57450);
  nand n57454(x57454, x56876, x57224);
  nand n57455(x57455, x56875, x57322);
  nand n57456(x57456, x57455, x57454);
  nand n57458(x57458, x56881, x57227);
  nand n57459(x57459, x56880, x57323);
  nand n57460(x57460, x57459, x57458);
  nand n57462(x57462, x56886, x57230);
  nand n57463(x57463, x56885, x57324);
  nand n57464(x57464, x57463, x57462);
  nand n57466(x57466, x56891, x57327);
  nand n57468(x57468, x56890, x57467);
  nand n57469(x57469, x57468, x57466);
  nand n57471(x57471, x56896, x57330);
  nand n57473(x57473, x56895, x57472);
  nand n57474(x57474, x57473, x57471);
  nand n57476(x57476, x56901, x57333);
  nand n57477(x57477, x56900, x57399);
  nand n57478(x57478, x57477, x57476);
  nand n57480(x57480, x56906, x57336);
  nand n57481(x57481, x56905, x57400);
  nand n57482(x57482, x57481, x57480);
  nand n57484(x57484, x56911, x57339);
  nand n57485(x57485, x56910, x57401);
  nand n57486(x57486, x57485, x57484);
  nand n57488(x57488, x56916, x57342);
  nand n57489(x57489, x56915, x57402);
  nand n57490(x57490, x57489, x57488);
  nand n57492(x57492, x56921, x57345);
  nand n57493(x57493, x56920, x57403);
  nand n57494(x57494, x57493, x57492);
  nand n57496(x57496, x56926, x57348);
  nand n57497(x57497, x56925, x57404);
  nand n57498(x57498, x57497, x57496);
  nand n57500(x57500, x56931, x57407);
  nand n57502(x57502, x56930, x57501);
  nand n57503(x57503, x57502, x57500);
  nand n57505(x57505, x56936, x57410);
  nand n57507(x57507, x56935, x57506);
  nand n57508(x57508, x57507, x57505);
  nand n57510(x57510, x56941, x57413);
  nand n57512(x57512, x56940, x57511);
  nand n57513(x57513, x57512, x57510);
  nand n57515(x57515, x56946, x57416);
  nand n57517(x57517, x56945, x57516);
  nand n57518(x57518, x57517, x57515);
  nand n57520(x57520, x56951, x57419);
  nand n57522(x57522, x56950, x57521);
  nand n57523(x57523, x57522, x57520);
  nand n57525(x57525, x56956, x57422);
  nand n57527(x57527, x56955, x57526);
  nand n57528(x57528, x57527, x57525);
  nand n57530(x57530, x56961, x57425);
  nand n57532(x57532, x56960, x57531);
  nand n57533(x57533, x57532, x57530);
  nand n57535(x57535, x56966, x57428);
  nand n57537(x57537, x56965, x57536);
  nand n57538(x57538, x57537, x57535);
  nand n57540(x57540, x56971, x57431);
  nand n57542(x57542, x56970, x57541);
  nand n57543(x57543, x57542, x57540);
  nand n57545(x57545, x56976, x57434);
  nand n57547(x57547, x56975, x57546);
  nand n57548(x57548, x57547, x57545);
  nand n57550(x57550, x50014, x50008);
  nand n57552(x57552, x50020, x50014);
  nand n57554(x57554, x50026, x50020);
  nand n57556(x57556, x50032, x50026);
  nand n57558(x57558, x50038, x50032);
  nand n57560(x57560, x50044, x50038);
  nand n57562(x57562, x50050, x50044);
  nand n57564(x57564, x50056, x50050);
  nand n57566(x57566, x50062, x50056);
  nand n57568(x57568, x50068, x50062);
  nand n57570(x57570, x50074, x50068);
  nand n57572(x57572, x50080, x50074);
  nand n57574(x57574, x50086, x50080);
  nand n57576(x57576, x50092, x50086);
  nand n57578(x57578, x50098, x50092);
  nand n57580(x57580, x50104, x50098);
  nand n57582(x57582, x50110, x50104);
  nand n57584(x57584, x50116, x50110);
  nand n57586(x57586, x50122, x50116);
  nand n57588(x57588, x50128, x50122);
  nand n57590(x57590, x50134, x50128);
  nand n57592(x57592, x50140, x50134);
  nand n57594(x57594, x50146, x50140);
  nand n57596(x57596, x50152, x50146);
  nand n57598(x57598, x50158, x50152);
  nand n57600(x57600, x50164, x50158);
  nand n57602(x57602, x50170, x50164);
  nand n57604(x57604, x50176, x50170);
  nand n57606(x57606, x50182, x50176);
  nand n57608(x57608, x50188, x50182);
  nand n57610(x57610, x57553, x50008);
  nand n57611(x57611, x57555, x57551);
  nand n57613(x57613, x57557, x57553);
  nand n57615(x57615, x57559, x57555);
  nand n57617(x57617, x57561, x57557);
  nand n57619(x57619, x57563, x57559);
  nand n57621(x57621, x57565, x57561);
  nand n57623(x57623, x57567, x57563);
  nand n57625(x57625, x57569, x57565);
  nand n57627(x57627, x57571, x57567);
  nand n57629(x57629, x57573, x57569);
  nand n57631(x57631, x57575, x57571);
  nand n57633(x57633, x57577, x57573);
  nand n57635(x57635, x57579, x57575);
  nand n57637(x57637, x57581, x57577);
  nand n57639(x57639, x57583, x57579);
  nand n57641(x57641, x57585, x57581);
  nand n57643(x57643, x57587, x57583);
  nand n57645(x57645, x57589, x57585);
  nand n57647(x57647, x57591, x57587);
  nand n57649(x57649, x57593, x57589);
  nand n57651(x57651, x57595, x57591);
  nand n57653(x57653, x57597, x57593);
  nand n57655(x57655, x57599, x57595);
  nand n57657(x57657, x57601, x57597);
  nand n57659(x57659, x57603, x57599);
  nand n57661(x57661, x57605, x57601);
  nand n57663(x57663, x57607, x57603);
  nand n57665(x57665, x57609, x57605);
  nand n57667(x57667, x57614, x50008);
  nand n57668(x57668, x57616, x57551);
  nand n57669(x57669, x57618, x85862);
  nand n57670(x57670, x57620, x57612);
  nand n57672(x57672, x57622, x57614);
  nand n57674(x57674, x57624, x57616);
  nand n57676(x57676, x57626, x57618);
  nand n57678(x57678, x57628, x57620);
  nand n57680(x57680, x57630, x57622);
  nand n57682(x57682, x57632, x57624);
  nand n57684(x57684, x57634, x57626);
  nand n57686(x57686, x57636, x57628);
  nand n57688(x57688, x57638, x57630);
  nand n57690(x57690, x57640, x57632);
  nand n57692(x57692, x57642, x57634);
  nand n57694(x57694, x57644, x57636);
  nand n57696(x57696, x57646, x57638);
  nand n57698(x57698, x57648, x57640);
  nand n57700(x57700, x57650, x57642);
  nand n57702(x57702, x57652, x57644);
  nand n57704(x57704, x57654, x57646);
  nand n57706(x57706, x57656, x57648);
  nand n57708(x57708, x57658, x57650);
  nand n57710(x57710, x57660, x57652);
  nand n57712(x57712, x57662, x57654);
  nand n57714(x57714, x57664, x57656);
  nand n57716(x57716, x57666, x57658);
  nand n57718(x57718, x57673, x50008);
  nand n57719(x57719, x57675, x57551);
  nand n57720(x57720, x57677, x85862);
  nand n57721(x57721, x57679, x57612);
  nand n57722(x57722, x57681, x85863);
  nand n57723(x57723, x57683, x85864);
  nand n57724(x57724, x57685, x85865);
  nand n57725(x57725, x57687, x57671);
  nand n57726(x57726, x57689, x57673);
  nand n57728(x57728, x57691, x57675);
  nand n57730(x57730, x57693, x57677);
  nand n57732(x57732, x57695, x57679);
  nand n57734(x57734, x57697, x57681);
  nand n57736(x57736, x57699, x57683);
  nand n57738(x57738, x57701, x57685);
  nand n57740(x57740, x57703, x57687);
  nand n57742(x57742, x57705, x57689);
  nand n57744(x57744, x57707, x57691);
  nand n57746(x57746, x57709, x57693);
  nand n57748(x57748, x57711, x57695);
  nand n57750(x57750, x57713, x57697);
  nand n57752(x57752, x57715, x57699);
  nand n57754(x57754, x57717, x57701);
  nand n57756(x57756, x57727, x50008);
  nand n57757(x57757, x57729, x57551);
  nand n57758(x57758, x57731, x85862);
  nand n57759(x57759, x57733, x57612);
  nand n57760(x57760, x57735, x85863);
  nand n57761(x57761, x57737, x85864);
  nand n57762(x57762, x57739, x85865);
  nand n57763(x57763, x57741, x57671);
  nand n57764(x57764, x57743, x85866);
  nand n57765(x57765, x57745, x85867);
  nand n57766(x57766, x57747, x85868);
  nand n57767(x57767, x57749, x85869);
  nand n57768(x57768, x57751, x85870);
  nand n57769(x57769, x57753, x85871);
  nand n57770(x57770, x57755, x85872);
  nand n57771(x57771, x73522, x73517);
  nand n57772(x57772, x57771, x57550);
  nand n57774(x57774, x50020, x57551);
  nand n57775(x57775, x73527, x57550);
  nand n57776(x57776, x57775, x57774);
  nand n57778(x57778, x50026, x85862);
  nand n57779(x57779, x73532, x57610);
  nand n57780(x57780, x57779, x57778);
  nand n57782(x57782, x50032, x57612);
  nand n57783(x57783, x73537, x57611);
  nand n57784(x57784, x57783, x57782);
  nand n57786(x57786, x50038, x85863);
  nand n57787(x57787, x73542, x57667);
  nand n57788(x57788, x57787, x57786);
  nand n57790(x57790, x50044, x85864);
  nand n57791(x57791, x73547, x57668);
  nand n57792(x57792, x57791, x57790);
  nand n57794(x57794, x50050, x85865);
  nand n57795(x57795, x73552, x57669);
  nand n57796(x57796, x57795, x57794);
  nand n57798(x57798, x50056, x57671);
  nand n57799(x57799, x73557, x57670);
  nand n57800(x57800, x57799, x57798);
  nand n57802(x57802, x50062, x85866);
  nand n57803(x57803, x73562, x57718);
  nand n57804(x57804, x57803, x57802);
  nand n57806(x57806, x50068, x85867);
  nand n57807(x57807, x73567, x57719);
  nand n57808(x57808, x57807, x57806);
  nand n57810(x57810, x50074, x85868);
  nand n57811(x57811, x73572, x57720);
  nand n57812(x57812, x57811, x57810);
  nand n57814(x57814, x50080, x85869);
  nand n57815(x57815, x73577, x57721);
  nand n57816(x57816, x57815, x57814);
  nand n57818(x57818, x50086, x85870);
  nand n57819(x57819, x73582, x57722);
  nand n57820(x57820, x57819, x57818);
  nand n57822(x57822, x50092, x85871);
  nand n57823(x57823, x73587, x57723);
  nand n57824(x57824, x57823, x57822);
  nand n57826(x57826, x50098, x85872);
  nand n57827(x57827, x73592, x57724);
  nand n57828(x57828, x57827, x57826);
  nand n57830(x57830, x50104, x85873);
  nand n57831(x57831, x73597, x57725);
  nand n57832(x57832, x57831, x57830);
  nand n57834(x57834, x50110, x85874);
  nand n57835(x57835, x73602, x57756);
  nand n57836(x57836, x57835, x57834);
  nand n57838(x57838, x50116, x85875);
  nand n57839(x57839, x73607, x57757);
  nand n57840(x57840, x57839, x57838);
  nand n57842(x57842, x50122, x85876);
  nand n57843(x57843, x73612, x57758);
  nand n57844(x57844, x57843, x57842);
  nand n57846(x57846, x50128, x85877);
  nand n57847(x57847, x73617, x57759);
  nand n57848(x57848, x57847, x57846);
  nand n57850(x57850, x50134, x85878);
  nand n57851(x57851, x73622, x57760);
  nand n57852(x57852, x57851, x57850);
  nand n57854(x57854, x50140, x85879);
  nand n57855(x57855, x73627, x57761);
  nand n57856(x57856, x57855, x57854);
  nand n57858(x57858, x50146, x85880);
  nand n57859(x57859, x73632, x57762);
  nand n57860(x57860, x57859, x57858);
  nand n57862(x57862, x50152, x85881);
  nand n57863(x57863, x73637, x57763);
  nand n57864(x57864, x57863, x57862);
  nand n57866(x57866, x50158, x85882);
  nand n57867(x57867, x73642, x57764);
  nand n57868(x57868, x57867, x57866);
  nand n57870(x57870, x50164, x85883);
  nand n57871(x57871, x73647, x57765);
  nand n57872(x57872, x57871, x57870);
  nand n57874(x57874, x50170, x85884);
  nand n57875(x57875, x73652, x57766);
  nand n57876(x57876, x57875, x57874);
  nand n57878(x57878, x50176, x85885);
  nand n57879(x57879, x73657, x57767);
  nand n57880(x57880, x57879, x57878);
  nand n57882(x57882, x50182, x85886);
  nand n57883(x57883, x73662, x57768);
  nand n57884(x57884, x57883, x57882);
  nand n57886(x57886, x50188, x85887);
  nand n57887(x57887, x73667, x57769);
  nand n57888(x57888, x57887, x57886);
  nand n57890(x57890, x50194, x85888);
  nand n57891(x57891, x73672, x57770);
  nand n57892(x57892, x57891, x57890);
  nand n57895(x57895, x73597, x49847);
  nand n57897(x57897, x73602, x49849);
  nand n57899(x57899, x73607, x49851);
  nand n57901(x57901, x73612, x49853);
  nand n57903(x57903, x73617, x49855);
  nand n57905(x57905, x73622, x49857);
  nand n57907(x57907, x73627, x49859);
  nand n57909(x57909, x73632, x49861);
  nand n57911(x57911, x73637, x49863);
  nand n57913(x57913, x73642, x49865);
  nand n57915(x57915, x73647, x49867);
  nand n57917(x57917, x73652, x49869);
  nand n57919(x57919, x73657, x49871);
  nand n57921(x57921, x73662, x49873);
  nand n57923(x57923, x73667, x49875);
  nand n57925(x57925, x73672, x49877);
  nand n57927(x57927, x50008, x49878);
  nand n57928(x57928, x50014, x49879);
  nand n57929(x57929, x50020, x49880);
  nand n57930(x57930, x50026, x49881);
  nand n57931(x57931, x50032, x49882);
  nand n57932(x57932, x50038, x49883);
  nand n57933(x57933, x50044, x49884);
  nand n57934(x57934, x50050, x49885);
  nand n57935(x57935, x50056, x49886);
  nand n57936(x57936, x50062, x49887);
  nand n57937(x57937, x50068, x49888);
  nand n57938(x57938, x50074, x49889);
  nand n57939(x57939, x50080, x49890);
  nand n57940(x57940, x50086, x49891);
  nand n57941(x57941, x50092, x49892);
  nand n57942(x57942, x50098, x49893);
  nand n57943(x57943, x50104, x49894);
  nand n57944(x57944, x50110, x49895);
  nand n57945(x57945, x50116, x49896);
  nand n57946(x57946, x50122, x49897);
  nand n57947(x57947, x50128, x49898);
  nand n57948(x57948, x50134, x49899);
  nand n57949(x57949, x50140, x49900);
  nand n57950(x57950, x50146, x49901);
  nand n57951(x57951, x50152, x49902);
  nand n57952(x57952, x50158, x49903);
  nand n57953(x57953, x50164, x49904);
  nand n57954(x57954, x50170, x49905);
  nand n57955(x57955, x50176, x49906);
  nand n57956(x57956, x50182, x49907);
  nand n57957(x57957, x50188, x49908);
  nand n57958(x57958, x50194, x49909);
  nand n57959(x57959, x57927, x50938);
  nand n57961(x57961, x57928, x50945);
  nand n57963(x57963, x57929, x50960);
  nand n57965(x57965, x57930, x50984);
  nand n57967(x57967, x57931, x51015);
  nand n57969(x57969, x57932, x51054);
  nand n57971(x57971, x57933, x51102);
  nand n57973(x57973, x57934, x51157);
  nand n57975(x57975, x57935, x51220);
  nand n57977(x57977, x57936, x51292);
  nand n57979(x57979, x57937, x51371);
  nand n57981(x57981, x57938, x51458);
  nand n57983(x57983, x57939, x51554);
  nand n57985(x57985, x57940, x51657);
  nand n57987(x57987, x57941, x51768);
  nand n57989(x57989, x57942, x51888);
  nand n57991(x57991, x57943, x57895);
  nand n57993(x57993, x57944, x57897);
  nand n57995(x57995, x57945, x57899);
  nand n57997(x57997, x57946, x57901);
  nand n57999(x57999, x57947, x57903);
  nand n58001(x58001, x57948, x57905);
  nand n58003(x58003, x57949, x57907);
  nand n58005(x58005, x57950, x57909);
  nand n58007(x58007, x57951, x57911);
  nand n58009(x58009, x57952, x57913);
  nand n58011(x58011, x57953, x57915);
  nand n58013(x58013, x57954, x57917);
  nand n58015(x58015, x57955, x57919);
  nand n58017(x58017, x57956, x57921);
  nand n58019(x58019, x57957, x57923);
  nand n58021(x58021, x57958, x57925);
  nand n58023(x58023, x49878, x73517);
  nand n58024(x58024, x49878, x73522);
  nand n58025(x58025, x58024, x50938);
  nand n58026(x58026, x49878, x73527);
  nand n58027(x58027, x58026, x50939);
  nand n58028(x58028, x49878, x73532);
  nand n58029(x58029, x58028, x50943);
  nand n58030(x58030, x49878, x73537);
  nand n58031(x58031, x58030, x50949);
  nand n58032(x58032, x49878, x73542);
  nand n58033(x58033, x58032, x50956);
  nand n58034(x58034, x49878, x73547);
  nand n58035(x58035, x58034, x50966);
  nand n58036(x58036, x49878, x73552);
  nand n58037(x58037, x58036, x50978);
  nand n58038(x58038, x49878, x73557);
  nand n58039(x58039, x58038, x50991);
  nand n58040(x58040, x49878, x73562);
  nand n58041(x58041, x58040, x51007);
  nand n58042(x58042, x49878, x73567);
  nand n58043(x58043, x58042, x51025);
  nand n58044(x58044, x49878, x73572);
  nand n58045(x58045, x58044, x51044);
  nand n58046(x58046, x49878, x73577);
  nand n58047(x58047, x58046, x51066);
  nand n58048(x58048, x49878, x73582);
  nand n58049(x58049, x58048, x51090);
  nand n58050(x58050, x49878, x73587);
  nand n58051(x58051, x58050, x51115);
  nand n58052(x58052, x49878, x73592);
  nand n58053(x58053, x58052, x51143);
  nand n58054(x58054, x49878, x73597);
  nand n58055(x58055, x58054, x51173);
  nand n58056(x58056, x49878, x73602);
  nand n58057(x58057, x58056, x51204);
  nand n58058(x58058, x49878, x73607);
  nand n58059(x58059, x58058, x51238);
  nand n58060(x58060, x49878, x73612);
  nand n58061(x58061, x58060, x51274);
  nand n58062(x58062, x49878, x73617);
  nand n58063(x58063, x58062, x51311);
  nand n58064(x58064, x49878, x73622);
  nand n58065(x58065, x58064, x51351);
  nand n58066(x58066, x49878, x73627);
  nand n58067(x58067, x58066, x51393);
  nand n58068(x58068, x49878, x73632);
  nand n58069(x58069, x58068, x51436);
  nand n58070(x58070, x49878, x73637);
  nand n58071(x58071, x58070, x51482);
  nand n58072(x58072, x49878, x73642);
  nand n58073(x58073, x58072, x51530);
  nand n58074(x58074, x49878, x73647);
  nand n58075(x58075, x58074, x51579);
  nand n58076(x58076, x49878, x73652);
  nand n58077(x58077, x58076, x51631);
  nand n58078(x58078, x49878, x73657);
  nand n58079(x58079, x58078, x51685);
  nand n58080(x58080, x49878, x73662);
  nand n58081(x58081, x58080, x51740);
  nand n58082(x58082, x49878, x73667);
  nand n58083(x58083, x58082, x51798);
  nand n58084(x58084, x49878, x73672);
  nand n58085(x58085, x58084, x51858);
  nand n58086(x58086, x49879, x85889);
  nand n58087(x58087, x49879, x58025);
  nand n58088(x58088, x49817, x85889);
  nand n58089(x58089, x49879, x58027);
  nand n58090(x58090, x58089, x58088);
  nand n58091(x58091, x49817, x58025);
  nand n58092(x58092, x49879, x58029);
  nand n58093(x58093, x58092, x58091);
  nand n58094(x58094, x49817, x58027);
  nand n58095(x58095, x49879, x58031);
  nand n58096(x58096, x58095, x58094);
  nand n58097(x58097, x49817, x58029);
  nand n58098(x58098, x49879, x58033);
  nand n58099(x58099, x58098, x58097);
  nand n58100(x58100, x49817, x58031);
  nand n58101(x58101, x49879, x58035);
  nand n58102(x58102, x58101, x58100);
  nand n58103(x58103, x49817, x58033);
  nand n58104(x58104, x49879, x58037);
  nand n58105(x58105, x58104, x58103);
  nand n58106(x58106, x49817, x58035);
  nand n58107(x58107, x49879, x58039);
  nand n58108(x58108, x58107, x58106);
  nand n58109(x58109, x49817, x58037);
  nand n58110(x58110, x49879, x58041);
  nand n58111(x58111, x58110, x58109);
  nand n58112(x58112, x49817, x58039);
  nand n58113(x58113, x49879, x58043);
  nand n58114(x58114, x58113, x58112);
  nand n58115(x58115, x49817, x58041);
  nand n58116(x58116, x49879, x58045);
  nand n58117(x58117, x58116, x58115);
  nand n58118(x58118, x49817, x58043);
  nand n58119(x58119, x49879, x58047);
  nand n58120(x58120, x58119, x58118);
  nand n58121(x58121, x49817, x58045);
  nand n58122(x58122, x49879, x58049);
  nand n58123(x58123, x58122, x58121);
  nand n58124(x58124, x49817, x58047);
  nand n58125(x58125, x49879, x58051);
  nand n58126(x58126, x58125, x58124);
  nand n58127(x58127, x49817, x58049);
  nand n58128(x58128, x49879, x58053);
  nand n58129(x58129, x58128, x58127);
  nand n58130(x58130, x49817, x58051);
  nand n58131(x58131, x49879, x58055);
  nand n58132(x58132, x58131, x58130);
  nand n58133(x58133, x49817, x58053);
  nand n58134(x58134, x49879, x58057);
  nand n58135(x58135, x58134, x58133);
  nand n58136(x58136, x49817, x58055);
  nand n58137(x58137, x49879, x58059);
  nand n58138(x58138, x58137, x58136);
  nand n58139(x58139, x49817, x58057);
  nand n58140(x58140, x49879, x58061);
  nand n58141(x58141, x58140, x58139);
  nand n58142(x58142, x49817, x58059);
  nand n58143(x58143, x49879, x58063);
  nand n58144(x58144, x58143, x58142);
  nand n58145(x58145, x49817, x58061);
  nand n58146(x58146, x49879, x58065);
  nand n58147(x58147, x58146, x58145);
  nand n58148(x58148, x49817, x58063);
  nand n58149(x58149, x49879, x58067);
  nand n58150(x58150, x58149, x58148);
  nand n58151(x58151, x49817, x58065);
  nand n58152(x58152, x49879, x58069);
  nand n58153(x58153, x58152, x58151);
  nand n58154(x58154, x49817, x58067);
  nand n58155(x58155, x49879, x58071);
  nand n58156(x58156, x58155, x58154);
  nand n58157(x58157, x49817, x58069);
  nand n58158(x58158, x49879, x58073);
  nand n58159(x58159, x58158, x58157);
  nand n58160(x58160, x49817, x58071);
  nand n58161(x58161, x49879, x58075);
  nand n58162(x58162, x58161, x58160);
  nand n58163(x58163, x49817, x58073);
  nand n58164(x58164, x49879, x58077);
  nand n58165(x58165, x58164, x58163);
  nand n58166(x58166, x49817, x58075);
  nand n58167(x58167, x49879, x58079);
  nand n58168(x58168, x58167, x58166);
  nand n58169(x58169, x49817, x58077);
  nand n58170(x58170, x49879, x58081);
  nand n58171(x58171, x58170, x58169);
  nand n58172(x58172, x49817, x58079);
  nand n58173(x58173, x49879, x58083);
  nand n58174(x58174, x58173, x58172);
  nand n58175(x58175, x49817, x58081);
  nand n58176(x58176, x49879, x58085);
  nand n58177(x58177, x58176, x58175);
  nand n58178(x58178, x49880, x85890);
  nand n58179(x58179, x49880, x85891);
  nand n58180(x58180, x49880, x58090);
  nand n58181(x58181, x49880, x58093);
  nand n58182(x58182, x49819, x85890);
  nand n58183(x58183, x49880, x58096);
  nand n58184(x58184, x58183, x58182);
  nand n58185(x58185, x49819, x85891);
  nand n58186(x58186, x49880, x58099);
  nand n58187(x58187, x58186, x58185);
  nand n58188(x58188, x49819, x58090);
  nand n58189(x58189, x49880, x58102);
  nand n58190(x58190, x58189, x58188);
  nand n58191(x58191, x49819, x58093);
  nand n58192(x58192, x49880, x58105);
  nand n58193(x58193, x58192, x58191);
  nand n58194(x58194, x49819, x58096);
  nand n58195(x58195, x49880, x58108);
  nand n58196(x58196, x58195, x58194);
  nand n58197(x58197, x49819, x58099);
  nand n58198(x58198, x49880, x58111);
  nand n58199(x58199, x58198, x58197);
  nand n58200(x58200, x49819, x58102);
  nand n58201(x58201, x49880, x58114);
  nand n58202(x58202, x58201, x58200);
  nand n58203(x58203, x49819, x58105);
  nand n58204(x58204, x49880, x58117);
  nand n58205(x58205, x58204, x58203);
  nand n58206(x58206, x49819, x58108);
  nand n58207(x58207, x49880, x58120);
  nand n58208(x58208, x58207, x58206);
  nand n58209(x58209, x49819, x58111);
  nand n58210(x58210, x49880, x58123);
  nand n58211(x58211, x58210, x58209);
  nand n58212(x58212, x49819, x58114);
  nand n58213(x58213, x49880, x58126);
  nand n58214(x58214, x58213, x58212);
  nand n58215(x58215, x49819, x58117);
  nand n58216(x58216, x49880, x58129);
  nand n58217(x58217, x58216, x58215);
  nand n58218(x58218, x49819, x58120);
  nand n58219(x58219, x49880, x58132);
  nand n58220(x58220, x58219, x58218);
  nand n58221(x58221, x49819, x58123);
  nand n58222(x58222, x49880, x58135);
  nand n58223(x58223, x58222, x58221);
  nand n58224(x58224, x49819, x58126);
  nand n58225(x58225, x49880, x58138);
  nand n58226(x58226, x58225, x58224);
  nand n58227(x58227, x49819, x58129);
  nand n58228(x58228, x49880, x58141);
  nand n58229(x58229, x58228, x58227);
  nand n58230(x58230, x49819, x58132);
  nand n58231(x58231, x49880, x58144);
  nand n58232(x58232, x58231, x58230);
  nand n58233(x58233, x49819, x58135);
  nand n58234(x58234, x49880, x58147);
  nand n58235(x58235, x58234, x58233);
  nand n58236(x58236, x49819, x58138);
  nand n58237(x58237, x49880, x58150);
  nand n58238(x58238, x58237, x58236);
  nand n58239(x58239, x49819, x58141);
  nand n58240(x58240, x49880, x58153);
  nand n58241(x58241, x58240, x58239);
  nand n58242(x58242, x49819, x58144);
  nand n58243(x58243, x49880, x58156);
  nand n58244(x58244, x58243, x58242);
  nand n58245(x58245, x49819, x58147);
  nand n58246(x58246, x49880, x58159);
  nand n58247(x58247, x58246, x58245);
  nand n58248(x58248, x49819, x58150);
  nand n58249(x58249, x49880, x58162);
  nand n58250(x58250, x58249, x58248);
  nand n58251(x58251, x49819, x58153);
  nand n58252(x58252, x49880, x58165);
  nand n58253(x58253, x58252, x58251);
  nand n58254(x58254, x49819, x58156);
  nand n58255(x58255, x49880, x58168);
  nand n58256(x58256, x58255, x58254);
  nand n58257(x58257, x49819, x58159);
  nand n58258(x58258, x49880, x58171);
  nand n58259(x58259, x58258, x58257);
  nand n58260(x58260, x49819, x58162);
  nand n58261(x58261, x49880, x58174);
  nand n58262(x58262, x58261, x58260);
  nand n58263(x58263, x49819, x58165);
  nand n58264(x58264, x49880, x58177);
  nand n58265(x58265, x58264, x58263);
  nand n58266(x58266, x49881, x85892);
  nand n58267(x58267, x49881, x85893);
  nand n58268(x58268, x49881, x85894);
  nand n58269(x58269, x49881, x85895);
  nand n58270(x58270, x49881, x58184);
  nand n58271(x58271, x49881, x58187);
  nand n58272(x58272, x49881, x58190);
  nand n58273(x58273, x49881, x58193);
  nand n58274(x58274, x49821, x85892);
  nand n58275(x58275, x49881, x58196);
  nand n58276(x58276, x58275, x58274);
  nand n58277(x58277, x49821, x85893);
  nand n58278(x58278, x49881, x58199);
  nand n58279(x58279, x58278, x58277);
  nand n58280(x58280, x49821, x85894);
  nand n58281(x58281, x49881, x58202);
  nand n58282(x58282, x58281, x58280);
  nand n58283(x58283, x49821, x85895);
  nand n58284(x58284, x49881, x58205);
  nand n58285(x58285, x58284, x58283);
  nand n58286(x58286, x49821, x58184);
  nand n58287(x58287, x49881, x58208);
  nand n58288(x58288, x58287, x58286);
  nand n58289(x58289, x49821, x58187);
  nand n58290(x58290, x49881, x58211);
  nand n58291(x58291, x58290, x58289);
  nand n58292(x58292, x49821, x58190);
  nand n58293(x58293, x49881, x58214);
  nand n58294(x58294, x58293, x58292);
  nand n58295(x58295, x49821, x58193);
  nand n58296(x58296, x49881, x58217);
  nand n58297(x58297, x58296, x58295);
  nand n58298(x58298, x49821, x58196);
  nand n58299(x58299, x49881, x58220);
  nand n58300(x58300, x58299, x58298);
  nand n58301(x58301, x49821, x58199);
  nand n58302(x58302, x49881, x58223);
  nand n58303(x58303, x58302, x58301);
  nand n58304(x58304, x49821, x58202);
  nand n58305(x58305, x49881, x58226);
  nand n58306(x58306, x58305, x58304);
  nand n58307(x58307, x49821, x58205);
  nand n58308(x58308, x49881, x58229);
  nand n58309(x58309, x58308, x58307);
  nand n58310(x58310, x49821, x58208);
  nand n58311(x58311, x49881, x58232);
  nand n58312(x58312, x58311, x58310);
  nand n58313(x58313, x49821, x58211);
  nand n58314(x58314, x49881, x58235);
  nand n58315(x58315, x58314, x58313);
  nand n58316(x58316, x49821, x58214);
  nand n58317(x58317, x49881, x58238);
  nand n58318(x58318, x58317, x58316);
  nand n58319(x58319, x49821, x58217);
  nand n58320(x58320, x49881, x58241);
  nand n58321(x58321, x58320, x58319);
  nand n58322(x58322, x49821, x58220);
  nand n58323(x58323, x49881, x58244);
  nand n58324(x58324, x58323, x58322);
  nand n58325(x58325, x49821, x58223);
  nand n58326(x58326, x49881, x58247);
  nand n58327(x58327, x58326, x58325);
  nand n58328(x58328, x49821, x58226);
  nand n58329(x58329, x49881, x58250);
  nand n58330(x58330, x58329, x58328);
  nand n58331(x58331, x49821, x58229);
  nand n58332(x58332, x49881, x58253);
  nand n58333(x58333, x58332, x58331);
  nand n58334(x58334, x49821, x58232);
  nand n58335(x58335, x49881, x58256);
  nand n58336(x58336, x58335, x58334);
  nand n58337(x58337, x49821, x58235);
  nand n58338(x58338, x49881, x58259);
  nand n58339(x58339, x58338, x58337);
  nand n58340(x58340, x49821, x58238);
  nand n58341(x58341, x49881, x58262);
  nand n58342(x58342, x58341, x58340);
  nand n58343(x58343, x49821, x58241);
  nand n58344(x58344, x49881, x58265);
  nand n58345(x58345, x58344, x58343);
  nand n58346(x58346, x49882, x85896);
  nand n58347(x58347, x49882, x85897);
  nand n58348(x58348, x49882, x85898);
  nand n58349(x58349, x49882, x85899);
  nand n58350(x58350, x49882, x85900);
  nand n58351(x58351, x49882, x85901);
  nand n58352(x58352, x49882, x85902);
  nand n58353(x58353, x49882, x85903);
  nand n58354(x58354, x49882, x58276);
  nand n58355(x58355, x49882, x58279);
  nand n58356(x58356, x49882, x58282);
  nand n58357(x58357, x49882, x58285);
  nand n58358(x58358, x49882, x58288);
  nand n58359(x58359, x49882, x58291);
  nand n58360(x58360, x49882, x58294);
  nand n58361(x58361, x49882, x58297);
  nand n58362(x58362, x49823, x85896);
  nand n58363(x58363, x49882, x58300);
  nand n58364(x58364, x58363, x58362);
  nand n58365(x58365, x49823, x85897);
  nand n58366(x58366, x49882, x58303);
  nand n58367(x58367, x58366, x58365);
  nand n58368(x58368, x49823, x85898);
  nand n58369(x58369, x49882, x58306);
  nand n58370(x58370, x58369, x58368);
  nand n58371(x58371, x49823, x85899);
  nand n58372(x58372, x49882, x58309);
  nand n58373(x58373, x58372, x58371);
  nand n58374(x58374, x49823, x85900);
  nand n58375(x58375, x49882, x58312);
  nand n58376(x58376, x58375, x58374);
  nand n58377(x58377, x49823, x85901);
  nand n58378(x58378, x49882, x58315);
  nand n58379(x58379, x58378, x58377);
  nand n58380(x58380, x49823, x85902);
  nand n58381(x58381, x49882, x58318);
  nand n58382(x58382, x58381, x58380);
  nand n58383(x58383, x49823, x85903);
  nand n58384(x58384, x49882, x58321);
  nand n58385(x58385, x58384, x58383);
  nand n58386(x58386, x49823, x58276);
  nand n58387(x58387, x49882, x58324);
  nand n58388(x58388, x58387, x58386);
  nand n58389(x58389, x49823, x58279);
  nand n58390(x58390, x49882, x58327);
  nand n58391(x58391, x58390, x58389);
  nand n58392(x58392, x49823, x58282);
  nand n58393(x58393, x49882, x58330);
  nand n58394(x58394, x58393, x58392);
  nand n58395(x58395, x49823, x58285);
  nand n58396(x58396, x49882, x58333);
  nand n58397(x58397, x58396, x58395);
  nand n58398(x58398, x49823, x58288);
  nand n58399(x58399, x49882, x58336);
  nand n58400(x58400, x58399, x58398);
  nand n58401(x58401, x49823, x58291);
  nand n58402(x58402, x49882, x58339);
  nand n58403(x58403, x58402, x58401);
  nand n58404(x58404, x49823, x58294);
  nand n58405(x58405, x49882, x58342);
  nand n58406(x58406, x58405, x58404);
  nand n58407(x58407, x49823, x58297);
  nand n58408(x58408, x49882, x58345);
  nand n58409(x58409, x58408, x58407);
  nand n58410(x58410, x58023, x50939);
  nand n58411(x58411, x58024, x50943);
  nand n58412(x58412, x58026, x50949);
  nand n58413(x58413, x58028, x50956);
  nand n58414(x58414, x58030, x50966);
  nand n58415(x58415, x58032, x50978);
  nand n58416(x58416, x58034, x50991);
  nand n58417(x58417, x58036, x51007);
  nand n58418(x58418, x58038, x51025);
  nand n58419(x58419, x58040, x51044);
  nand n58420(x58420, x58042, x51066);
  nand n58421(x58421, x58044, x51090);
  nand n58422(x58422, x58046, x51115);
  nand n58423(x58423, x58048, x51143);
  nand n58424(x58424, x58050, x51173);
  nand n58425(x58425, x58052, x51204);
  nand n58426(x58426, x58054, x51238);
  nand n58427(x58427, x58056, x51274);
  nand n58428(x58428, x58058, x51311);
  nand n58429(x58429, x58060, x51351);
  nand n58430(x58430, x58062, x51393);
  nand n58431(x58431, x58064, x51436);
  nand n58432(x58432, x58066, x51482);
  nand n58433(x58433, x58068, x51530);
  nand n58434(x58434, x58070, x51579);
  nand n58435(x58435, x58072, x51631);
  nand n58436(x58436, x58074, x51685);
  nand n58437(x58437, x58076, x51740);
  nand n58438(x58438, x58078, x51798);
  nand n58439(x58439, x58080, x51858);
  nand n58440(x58440, x58082, x51919);
  nand n58441(x58441, x49817, x58412);
  nand n58442(x58442, x49879, x58410);
  nand n58443(x58443, x58442, x58441);
  nand n58444(x58444, x49817, x58413);
  nand n58445(x58445, x49879, x58411);
  nand n58446(x58446, x58445, x58444);
  nand n58447(x58447, x49817, x58414);
  nand n58448(x58448, x49879, x58412);
  nand n58449(x58449, x58448, x58447);
  nand n58450(x58450, x49817, x58415);
  nand n58451(x58451, x49879, x58413);
  nand n58452(x58452, x58451, x58450);
  nand n58453(x58453, x49817, x58416);
  nand n58454(x58454, x49879, x58414);
  nand n58455(x58455, x58454, x58453);
  nand n58456(x58456, x49817, x58417);
  nand n58457(x58457, x49879, x58415);
  nand n58458(x58458, x58457, x58456);
  nand n58459(x58459, x49817, x58418);
  nand n58460(x58460, x49879, x58416);
  nand n58461(x58461, x58460, x58459);
  nand n58462(x58462, x49817, x58419);
  nand n58463(x58463, x49879, x58417);
  nand n58464(x58464, x58463, x58462);
  nand n58465(x58465, x49817, x58420);
  nand n58466(x58466, x49879, x58418);
  nand n58467(x58467, x58466, x58465);
  nand n58468(x58468, x49817, x58421);
  nand n58469(x58469, x49879, x58419);
  nand n58470(x58470, x58469, x58468);
  nand n58471(x58471, x49817, x58422);
  nand n58472(x58472, x49879, x58420);
  nand n58473(x58473, x58472, x58471);
  nand n58474(x58474, x49817, x58423);
  nand n58475(x58475, x49879, x58421);
  nand n58476(x58476, x58475, x58474);
  nand n58477(x58477, x49817, x58424);
  nand n58478(x58478, x49879, x58422);
  nand n58479(x58479, x58478, x58477);
  nand n58480(x58480, x49817, x58425);
  nand n58481(x58481, x49879, x58423);
  nand n58482(x58482, x58481, x58480);
  nand n58483(x58483, x49817, x58426);
  nand n58484(x58484, x49879, x58424);
  nand n58485(x58485, x58484, x58483);
  nand n58486(x58486, x49817, x58427);
  nand n58487(x58487, x49879, x58425);
  nand n58488(x58488, x58487, x58486);
  nand n58489(x58489, x49817, x58428);
  nand n58490(x58490, x49879, x58426);
  nand n58491(x58491, x58490, x58489);
  nand n58492(x58492, x49817, x58429);
  nand n58493(x58493, x49879, x58427);
  nand n58494(x58494, x58493, x58492);
  nand n58495(x58495, x49817, x58430);
  nand n58496(x58496, x49879, x58428);
  nand n58497(x58497, x58496, x58495);
  nand n58498(x58498, x49817, x58431);
  nand n58499(x58499, x49879, x58429);
  nand n58500(x58500, x58499, x58498);
  nand n58501(x58501, x49817, x58432);
  nand n58502(x58502, x49879, x58430);
  nand n58503(x58503, x58502, x58501);
  nand n58504(x58504, x49817, x58433);
  nand n58505(x58505, x49879, x58431);
  nand n58506(x58506, x58505, x58504);
  nand n58507(x58507, x49817, x58434);
  nand n58508(x58508, x49879, x58432);
  nand n58509(x58509, x58508, x58507);
  nand n58510(x58510, x49817, x58435);
  nand n58511(x58511, x49879, x58433);
  nand n58512(x58512, x58511, x58510);
  nand n58513(x58513, x49817, x58436);
  nand n58514(x58514, x49879, x58434);
  nand n58515(x58515, x58514, x58513);
  nand n58516(x58516, x49817, x58437);
  nand n58517(x58517, x49879, x58435);
  nand n58518(x58518, x58517, x58516);
  nand n58519(x58519, x49817, x58438);
  nand n58520(x58520, x49879, x58436);
  nand n58521(x58521, x58520, x58519);
  nand n58522(x58522, x49817, x58439);
  nand n58523(x58523, x49879, x58437);
  nand n58524(x58524, x58523, x58522);
  nand n58525(x58525, x49817, x58440);
  nand n58526(x58526, x49879, x58438);
  nand n58527(x58527, x58526, x58525);
  nand n58528(x58528, x49817, x85920);
  nand n58529(x58529, x49879, x58439);
  nand n58530(x58530, x58529, x58528);
  nand n58531(x58531, x49879, x58440);
  nand n58532(x58532, x49879, x85920);
  nand n58533(x58533, x49819, x58455);
  nand n58534(x58534, x49880, x58443);
  nand n58535(x58535, x58534, x58533);
  nand n58536(x58536, x49819, x58458);
  nand n58537(x58537, x49880, x58446);
  nand n58538(x58538, x58537, x58536);
  nand n58539(x58539, x49819, x58461);
  nand n58540(x58540, x49880, x58449);
  nand n58541(x58541, x58540, x58539);
  nand n58542(x58542, x49819, x58464);
  nand n58543(x58543, x49880, x58452);
  nand n58544(x58544, x58543, x58542);
  nand n58545(x58545, x49819, x58467);
  nand n58546(x58546, x49880, x58455);
  nand n58547(x58547, x58546, x58545);
  nand n58548(x58548, x49819, x58470);
  nand n58549(x58549, x49880, x58458);
  nand n58550(x58550, x58549, x58548);
  nand n58551(x58551, x49819, x58473);
  nand n58552(x58552, x49880, x58461);
  nand n58553(x58553, x58552, x58551);
  nand n58554(x58554, x49819, x58476);
  nand n58555(x58555, x49880, x58464);
  nand n58556(x58556, x58555, x58554);
  nand n58557(x58557, x49819, x58479);
  nand n58558(x58558, x49880, x58467);
  nand n58559(x58559, x58558, x58557);
  nand n58560(x58560, x49819, x58482);
  nand n58561(x58561, x49880, x58470);
  nand n58562(x58562, x58561, x58560);
  nand n58563(x58563, x49819, x58485);
  nand n58564(x58564, x49880, x58473);
  nand n58565(x58565, x58564, x58563);
  nand n58566(x58566, x49819, x58488);
  nand n58567(x58567, x49880, x58476);
  nand n58568(x58568, x58567, x58566);
  nand n58569(x58569, x49819, x58491);
  nand n58570(x58570, x49880, x58479);
  nand n58571(x58571, x58570, x58569);
  nand n58572(x58572, x49819, x58494);
  nand n58573(x58573, x49880, x58482);
  nand n58574(x58574, x58573, x58572);
  nand n58575(x58575, x49819, x58497);
  nand n58576(x58576, x49880, x58485);
  nand n58577(x58577, x58576, x58575);
  nand n58578(x58578, x49819, x58500);
  nand n58579(x58579, x49880, x58488);
  nand n58580(x58580, x58579, x58578);
  nand n58581(x58581, x49819, x58503);
  nand n58582(x58582, x49880, x58491);
  nand n58583(x58583, x58582, x58581);
  nand n58584(x58584, x49819, x58506);
  nand n58585(x58585, x49880, x58494);
  nand n58586(x58586, x58585, x58584);
  nand n58587(x58587, x49819, x58509);
  nand n58588(x58588, x49880, x58497);
  nand n58589(x58589, x58588, x58587);
  nand n58590(x58590, x49819, x58512);
  nand n58591(x58591, x49880, x58500);
  nand n58592(x58592, x58591, x58590);
  nand n58593(x58593, x49819, x58515);
  nand n58594(x58594, x49880, x58503);
  nand n58595(x58595, x58594, x58593);
  nand n58596(x58596, x49819, x58518);
  nand n58597(x58597, x49880, x58506);
  nand n58598(x58598, x58597, x58596);
  nand n58599(x58599, x49819, x58521);
  nand n58600(x58600, x49880, x58509);
  nand n58601(x58601, x58600, x58599);
  nand n58602(x58602, x49819, x58524);
  nand n58603(x58603, x49880, x58512);
  nand n58604(x58604, x58603, x58602);
  nand n58605(x58605, x49819, x58527);
  nand n58606(x58606, x49880, x58515);
  nand n58607(x58607, x58606, x58605);
  nand n58608(x58608, x49819, x58530);
  nand n58609(x58609, x49880, x58518);
  nand n58610(x58610, x58609, x58608);
  nand n58611(x58611, x49819, x85921);
  nand n58612(x58612, x49880, x58521);
  nand n58613(x58613, x58612, x58611);
  nand n58614(x58614, x49819, x85922);
  nand n58615(x58615, x49880, x58524);
  nand n58616(x58616, x58615, x58614);
  nand n58617(x58617, x49880, x58527);
  nand n58618(x58618, x49880, x58530);
  nand n58619(x58619, x49880, x85921);
  nand n58620(x58620, x49880, x85922);
  nand n58621(x58621, x49821, x58559);
  nand n58622(x58622, x49881, x58535);
  nand n58623(x58623, x58622, x58621);
  nand n58624(x58624, x49821, x58562);
  nand n58625(x58625, x49881, x58538);
  nand n58626(x58626, x58625, x58624);
  nand n58627(x58627, x49821, x58565);
  nand n58628(x58628, x49881, x58541);
  nand n58629(x58629, x58628, x58627);
  nand n58630(x58630, x49821, x58568);
  nand n58631(x58631, x49881, x58544);
  nand n58632(x58632, x58631, x58630);
  nand n58633(x58633, x49821, x58571);
  nand n58634(x58634, x49881, x58547);
  nand n58635(x58635, x58634, x58633);
  nand n58636(x58636, x49821, x58574);
  nand n58637(x58637, x49881, x58550);
  nand n58638(x58638, x58637, x58636);
  nand n58639(x58639, x49821, x58577);
  nand n58640(x58640, x49881, x58553);
  nand n58641(x58641, x58640, x58639);
  nand n58642(x58642, x49821, x58580);
  nand n58643(x58643, x49881, x58556);
  nand n58644(x58644, x58643, x58642);
  nand n58645(x58645, x49821, x58583);
  nand n58646(x58646, x49881, x58559);
  nand n58647(x58647, x58646, x58645);
  nand n58648(x58648, x49821, x58586);
  nand n58649(x58649, x49881, x58562);
  nand n58650(x58650, x58649, x58648);
  nand n58651(x58651, x49821, x58589);
  nand n58652(x58652, x49881, x58565);
  nand n58653(x58653, x58652, x58651);
  nand n58654(x58654, x49821, x58592);
  nand n58655(x58655, x49881, x58568);
  nand n58656(x58656, x58655, x58654);
  nand n58657(x58657, x49821, x58595);
  nand n58658(x58658, x49881, x58571);
  nand n58659(x58659, x58658, x58657);
  nand n58660(x58660, x49821, x58598);
  nand n58661(x58661, x49881, x58574);
  nand n58662(x58662, x58661, x58660);
  nand n58663(x58663, x49821, x58601);
  nand n58664(x58664, x49881, x58577);
  nand n58665(x58665, x58664, x58663);
  nand n58666(x58666, x49821, x58604);
  nand n58667(x58667, x49881, x58580);
  nand n58668(x58668, x58667, x58666);
  nand n58669(x58669, x49821, x58607);
  nand n58670(x58670, x49881, x58583);
  nand n58671(x58671, x58670, x58669);
  nand n58672(x58672, x49821, x58610);
  nand n58673(x58673, x49881, x58586);
  nand n58674(x58674, x58673, x58672);
  nand n58675(x58675, x49821, x58613);
  nand n58676(x58676, x49881, x58589);
  nand n58677(x58677, x58676, x58675);
  nand n58678(x58678, x49821, x58616);
  nand n58679(x58679, x49881, x58592);
  nand n58680(x58680, x58679, x58678);
  nand n58681(x58681, x49821, x85923);
  nand n58682(x58682, x49881, x58595);
  nand n58683(x58683, x58682, x58681);
  nand n58684(x58684, x49821, x85924);
  nand n58685(x58685, x49881, x58598);
  nand n58686(x58686, x58685, x58684);
  nand n58687(x58687, x49821, x85925);
  nand n58688(x58688, x49881, x58601);
  nand n58689(x58689, x58688, x58687);
  nand n58690(x58690, x49821, x85926);
  nand n58691(x58691, x49881, x58604);
  nand n58692(x58692, x58691, x58690);
  nand n58693(x58693, x49881, x58607);
  nand n58694(x58694, x49881, x58610);
  nand n58695(x58695, x49881, x58613);
  nand n58696(x58696, x49881, x58616);
  nand n58697(x58697, x49881, x85923);
  nand n58698(x58698, x49881, x85924);
  nand n58699(x58699, x49881, x85925);
  nand n58700(x58700, x49881, x85926);
  nand n58701(x58701, x49823, x58671);
  nand n58702(x58702, x49882, x58623);
  nand n58703(x58703, x58702, x58701);
  nand n58704(x58704, x49823, x58674);
  nand n58705(x58705, x49882, x58626);
  nand n58706(x58706, x58705, x58704);
  nand n58707(x58707, x49823, x58677);
  nand n58708(x58708, x49882, x58629);
  nand n58709(x58709, x58708, x58707);
  nand n58710(x58710, x49823, x58680);
  nand n58711(x58711, x49882, x58632);
  nand n58712(x58712, x58711, x58710);
  nand n58713(x58713, x49823, x58683);
  nand n58714(x58714, x49882, x58635);
  nand n58715(x58715, x58714, x58713);
  nand n58716(x58716, x49823, x58686);
  nand n58717(x58717, x49882, x58638);
  nand n58718(x58718, x58717, x58716);
  nand n58719(x58719, x49823, x58689);
  nand n58720(x58720, x49882, x58641);
  nand n58721(x58721, x58720, x58719);
  nand n58722(x58722, x49823, x58692);
  nand n58723(x58723, x49882, x58644);
  nand n58724(x58724, x58723, x58722);
  nand n58725(x58725, x49823, x85927);
  nand n58726(x58726, x49882, x58647);
  nand n58727(x58727, x58726, x58725);
  nand n58728(x58728, x49823, x85928);
  nand n58729(x58729, x49882, x58650);
  nand n58730(x58730, x58729, x58728);
  nand n58731(x58731, x49823, x85929);
  nand n58732(x58732, x49882, x58653);
  nand n58733(x58733, x58732, x58731);
  nand n58734(x58734, x49823, x85930);
  nand n58735(x58735, x49882, x58656);
  nand n58736(x58736, x58735, x58734);
  nand n58737(x58737, x49823, x85931);
  nand n58738(x58738, x49882, x58659);
  nand n58739(x58739, x58738, x58737);
  nand n58740(x58740, x49823, x85932);
  nand n58741(x58741, x49882, x58662);
  nand n58742(x58742, x58741, x58740);
  nand n58743(x58743, x49823, x85933);
  nand n58744(x58744, x49882, x58665);
  nand n58745(x58745, x58744, x58743);
  nand n58746(x58746, x49823, x85934);
  nand n58747(x58747, x49882, x58668);
  nand n58748(x58748, x58747, x58746);
  nand n58749(x58749, x49882, x58671);
  nand n58750(x58750, x49882, x58674);
  nand n58751(x58751, x49882, x58677);
  nand n58752(x58752, x49882, x58680);
  nand n58753(x58753, x49882, x58683);
  nand n58754(x58754, x49882, x58686);
  nand n58755(x58755, x49882, x58689);
  nand n58756(x58756, x49882, x58692);
  nand n58757(x58757, x49882, x85927);
  nand n58758(x58758, x49882, x85928);
  nand n58759(x58759, x49882, x85929);
  nand n58760(x58760, x49882, x85930);
  nand n58761(x58761, x49882, x85931);
  nand n58762(x58762, x49882, x85932);
  nand n58763(x58763, x49882, x85933);
  nand n58764(x58764, x49882, x85934);
  nand n58765(x58765, x71977, x49815);
  nand n58766(x58766, x16876, x58703);
  nand n58767(x58767, x58766, x25733);
  nand n58768(x58768, x71977, x85904);
  nand n58769(x58769, x16876, x57894);
  nand n58770(x58770, x71977, x50782);
  nand n58771(x58771, x16876, x50782);
  nand n58772(x58772, x58771, x58770);
  nand n58773(x58773, x71977, x57960);
  nand n58774(x58774, x16876, x57927);
  nand n58775(x58775, x58774, x58773);
  nand n58776(x58776, x71977, x57894);
  nand n58777(x58777, x58766, x58776);
  nand n58778(x58778, x16876, x50008);
  nand n58779(x58779, x58778, x58776);
  nand n58780(x58780, x71977, x73517);
  nand n58781(x58781, x25749, x85951);
  nand n58782(x58782, x71982, x58767);
  nand n58783(x58783, x25749, x85952);
  nand n58784(x58784, x58783, x58782);
  nand n58785(x58785, x71982, x85953);
  nand n58786(x58786, x25749, x58772);
  nand n58787(x58787, x58786, x58785);
  nand n58788(x58788, x71982, x58775);
  nand n58789(x58789, x25749, x58777);
  nand n58790(x58790, x58789, x58788);
  nand n58791(x58791, x71982, x85952);
  nand n58792(x58792, x25749, x85953);
  nand n58793(x58793, x58792, x58791);
  nand n58794(x58794, x71982, x58772);
  nand n58795(x58795, x25749, x58775);
  nand n58796(x58796, x58795, x58794);
  nand n58797(x58797, x71982, x58779);
  nand n58798(x58798, x25749, x85954);
  nand n58799(x58799, x58798, x58797);
  nand n58800(x58800, x71987, x85955);
  nand n58801(x58801, x25772, x58784);
  nand n58802(x58802, x58801, x25771);
  nand n58803(x58803, x71987, x58787);
  nand n58804(x58804, x25772, x58790);
  nand n58805(x58805, x58804, x58803);
  nand n58806(x58806, x71987, x58793);
  nand n58807(x58807, x25772, x58796);
  nand n58808(x58808, x58807, x58806);
  nand n58809(x58809, x71987, x58799);
  nand n58810(x58810, x25782, x85956);
  nand n58811(x58811, x71992, x58802);
  nand n58812(x58812, x25782, x58805);
  nand n58813(x58813, x58812, x58811);
  nand n58814(x58814, x71992, x58808);
  nand n58815(x58815, x25782, x85957);
  nand n58816(x58816, x58815, x58814);
  nand n58817(x58817, x25790, x85958);
  nand n58818(x58818, x71997, x58813);
  nand n58819(x58819, x25790, x58816);
  nand n58820(x58820, x58819, x58818);
  nand n58821(x58821, x72002, x85959);
  nand n58822(x58822, x25796, x58820);
  nand n58823(x58823, x58822, x58821);
  nand n58824(x58824, x71977, x49817);
  nand n58825(x58825, x16876, x58706);
  nand n58826(x58826, x58825, x25801);
  nand n58827(x58827, x71977, x85905);
  nand n58828(x58828, x16876, x85857);
  nand n58829(x58829, x71977, x50787);
  nand n58830(x58830, x16876, x50787);
  nand n58831(x58831, x58830, x58829);
  nand n58832(x58832, x71977, x57962);
  nand n58833(x58833, x16876, x57928);
  nand n58834(x58834, x58833, x58832);
  nand n58835(x58835, x71977, x50946);
  nand n58836(x58836, x58825, x58835);
  nand n58837(x58837, x16876, x50014);
  nand n58838(x58838, x58837, x58835);
  nand n58839(x58839, x71977, x57773);
  nand n58840(x58840, x25749, x85960);
  nand n58841(x58841, x71982, x58826);
  nand n58842(x58842, x25749, x85961);
  nand n58843(x58843, x58842, x58841);
  nand n58844(x58844, x71982, x85962);
  nand n58845(x58845, x25749, x58831);
  nand n58846(x58846, x58845, x58844);
  nand n58847(x58847, x71982, x58834);
  nand n58848(x58848, x25749, x58836);
  nand n58849(x58849, x58848, x58847);
  nand n58850(x58850, x71982, x85961);
  nand n58851(x58851, x25749, x85962);
  nand n58852(x58852, x58851, x58850);
  nand n58853(x58853, x71982, x58831);
  nand n58854(x58854, x25749, x58834);
  nand n58855(x58855, x58854, x58853);
  nand n58856(x58856, x71982, x58838);
  nand n58857(x58857, x25749, x85963);
  nand n58858(x58858, x58857, x58856);
  nand n58859(x58859, x71987, x85964);
  nand n58860(x58860, x25772, x58843);
  nand n58861(x58861, x58860, x25838);
  nand n58862(x58862, x71987, x58846);
  nand n58863(x58863, x25772, x58849);
  nand n58864(x58864, x58863, x58862);
  nand n58865(x58865, x71987, x58852);
  nand n58866(x58866, x25772, x58855);
  nand n58867(x58867, x58866, x58865);
  nand n58868(x58868, x71987, x58858);
  nand n58869(x58869, x25782, x85965);
  nand n58870(x58870, x71992, x58861);
  nand n58871(x58871, x25782, x58864);
  nand n58872(x58872, x58871, x58870);
  nand n58873(x58873, x71992, x58867);
  nand n58874(x58874, x25782, x85966);
  nand n58875(x58875, x58874, x58873);
  nand n58876(x58876, x25790, x85967);
  nand n58877(x58877, x71997, x58872);
  nand n58878(x58878, x25790, x58875);
  nand n58879(x58879, x58878, x58877);
  nand n58880(x58880, x72002, x85968);
  nand n58881(x58881, x25796, x58879);
  nand n58882(x58882, x58881, x58880);
  nand n58883(x58883, x71977, x49819);
  nand n58884(x58884, x16876, x58709);
  nand n58885(x58885, x58884, x25864);
  nand n58886(x58886, x71977, x85906);
  nand n58887(x58887, x16876, x85858);
  nand n58888(x58888, x71977, x50792);
  nand n58889(x58889, x16876, x50792);
  nand n58890(x58890, x58889, x58888);
  nand n58891(x58891, x71977, x57964);
  nand n58892(x58892, x16876, x57929);
  nand n58893(x58893, x58892, x58891);
  nand n58894(x58894, x71977, x50961);
  nand n58895(x58895, x58884, x58894);
  nand n58896(x58896, x16876, x50020);
  nand n58897(x58897, x58896, x58894);
  nand n58898(x58898, x71977, x57777);
  nand n58899(x58899, x25749, x85969);
  nand n58900(x58900, x71982, x58885);
  nand n58901(x58901, x25749, x85970);
  nand n58902(x58902, x58901, x58900);
  nand n58903(x58903, x71982, x85971);
  nand n58904(x58904, x25749, x58890);
  nand n58905(x58905, x58904, x58903);
  nand n58906(x58906, x71982, x58893);
  nand n58907(x58907, x25749, x58895);
  nand n58908(x58908, x58907, x58906);
  nand n58909(x58909, x71982, x85970);
  nand n58910(x58910, x25749, x85971);
  nand n58911(x58911, x58910, x58909);
  nand n58912(x58912, x71982, x58890);
  nand n58913(x58913, x25749, x58893);
  nand n58914(x58914, x58913, x58912);
  nand n58915(x58915, x71982, x58897);
  nand n58916(x58916, x25749, x85972);
  nand n58917(x58917, x58916, x58915);
  nand n58918(x58918, x71987, x85973);
  nand n58919(x58919, x25772, x58902);
  nand n58920(x58920, x58919, x25901);
  nand n58921(x58921, x71987, x58905);
  nand n58922(x58922, x25772, x58908);
  nand n58923(x58923, x58922, x58921);
  nand n58924(x58924, x71987, x58911);
  nand n58925(x58925, x25772, x58914);
  nand n58926(x58926, x58925, x58924);
  nand n58927(x58927, x71987, x58917);
  nand n58928(x58928, x25782, x85974);
  nand n58929(x58929, x71992, x58920);
  nand n58930(x58930, x25782, x58923);
  nand n58931(x58931, x58930, x58929);
  nand n58932(x58932, x71992, x58926);
  nand n58933(x58933, x25782, x85975);
  nand n58934(x58934, x58933, x58932);
  nand n58935(x58935, x25790, x85976);
  nand n58936(x58936, x71997, x58931);
  nand n58937(x58937, x25790, x58934);
  nand n58938(x58938, x58937, x58936);
  nand n58939(x58939, x72002, x85977);
  nand n58940(x58940, x25796, x58938);
  nand n58941(x58941, x58940, x58939);
  nand n58942(x58942, x71977, x49821);
  nand n58943(x58943, x16876, x58712);
  nand n58944(x58944, x58943, x25927);
  nand n58945(x58945, x71977, x85907);
  nand n58946(x58946, x16876, x85859);
  nand n58947(x58947, x71977, x50797);
  nand n58948(x58948, x16876, x50797);
  nand n58949(x58949, x58948, x58947);
  nand n58950(x58950, x71977, x57966);
  nand n58951(x58951, x16876, x57930);
  nand n58952(x58952, x58951, x58950);
  nand n58953(x58953, x71977, x50985);
  nand n58954(x58954, x58943, x58953);
  nand n58955(x58955, x16876, x50026);
  nand n58956(x58956, x58955, x58953);
  nand n58957(x58957, x71977, x57781);
  nand n58958(x58958, x25749, x85978);
  nand n58959(x58959, x71982, x58944);
  nand n58960(x58960, x25749, x85979);
  nand n58961(x58961, x58960, x58959);
  nand n58962(x58962, x71982, x85980);
  nand n58963(x58963, x25749, x58949);
  nand n58964(x58964, x58963, x58962);
  nand n58965(x58965, x71982, x58952);
  nand n58966(x58966, x25749, x58954);
  nand n58967(x58967, x58966, x58965);
  nand n58968(x58968, x71982, x85979);
  nand n58969(x58969, x25749, x85980);
  nand n58970(x58970, x58969, x58968);
  nand n58971(x58971, x71982, x58949);
  nand n58972(x58972, x25749, x58952);
  nand n58973(x58973, x58972, x58971);
  nand n58974(x58974, x71982, x58956);
  nand n58975(x58975, x25749, x85981);
  nand n58976(x58976, x58975, x58974);
  nand n58977(x58977, x71987, x85982);
  nand n58978(x58978, x25772, x58961);
  nand n58979(x58979, x58978, x25964);
  nand n58980(x58980, x71987, x58964);
  nand n58981(x58981, x25772, x58967);
  nand n58982(x58982, x58981, x58980);
  nand n58983(x58983, x71987, x58970);
  nand n58984(x58984, x25772, x58973);
  nand n58985(x58985, x58984, x58983);
  nand n58986(x58986, x71987, x58976);
  nand n58987(x58987, x25782, x85983);
  nand n58988(x58988, x71992, x58979);
  nand n58989(x58989, x25782, x58982);
  nand n58990(x58990, x58989, x58988);
  nand n58991(x58991, x71992, x58985);
  nand n58992(x58992, x25782, x85984);
  nand n58993(x58993, x58992, x58991);
  nand n58994(x58994, x25790, x85985);
  nand n58995(x58995, x71997, x58990);
  nand n58996(x58996, x25790, x58993);
  nand n58997(x58997, x58996, x58995);
  nand n58998(x58998, x72002, x85986);
  nand n58999(x58999, x25796, x58997);
  nand n59000(x59000, x58999, x58998);
  nand n59001(x59001, x71977, x49823);
  nand n59002(x59002, x16876, x58715);
  nand n59003(x59003, x59002, x25990);
  nand n59004(x59004, x71977, x85908);
  nand n59005(x59005, x16876, x85860);
  nand n59006(x59006, x71977, x50802);
  nand n59007(x59007, x16876, x50802);
  nand n59008(x59008, x59007, x59006);
  nand n59009(x59009, x71977, x57968);
  nand n59010(x59010, x16876, x57931);
  nand n59011(x59011, x59010, x59009);
  nand n59012(x59012, x71977, x51016);
  nand n59013(x59013, x59002, x59012);
  nand n59014(x59014, x16876, x50032);
  nand n59015(x59015, x59014, x59012);
  nand n59016(x59016, x71977, x57785);
  nand n59017(x59017, x25749, x85987);
  nand n59018(x59018, x71982, x59003);
  nand n59019(x59019, x25749, x85988);
  nand n59020(x59020, x59019, x59018);
  nand n59021(x59021, x71982, x85989);
  nand n59022(x59022, x25749, x59008);
  nand n59023(x59023, x59022, x59021);
  nand n59024(x59024, x71982, x59011);
  nand n59025(x59025, x25749, x59013);
  nand n59026(x59026, x59025, x59024);
  nand n59027(x59027, x71982, x85988);
  nand n59028(x59028, x25749, x85989);
  nand n59029(x59029, x59028, x59027);
  nand n59030(x59030, x71982, x59008);
  nand n59031(x59031, x25749, x59011);
  nand n59032(x59032, x59031, x59030);
  nand n59033(x59033, x71982, x59015);
  nand n59034(x59034, x25749, x85990);
  nand n59035(x59035, x59034, x59033);
  nand n59036(x59036, x71987, x85991);
  nand n59037(x59037, x25772, x59020);
  nand n59038(x59038, x59037, x26027);
  nand n59039(x59039, x71987, x59023);
  nand n59040(x59040, x25772, x59026);
  nand n59041(x59041, x59040, x59039);
  nand n59042(x59042, x71987, x59029);
  nand n59043(x59043, x25772, x59032);
  nand n59044(x59044, x59043, x59042);
  nand n59045(x59045, x71987, x59035);
  nand n59046(x59046, x25782, x85992);
  nand n59047(x59047, x71992, x59038);
  nand n59048(x59048, x25782, x59041);
  nand n59049(x59049, x59048, x59047);
  nand n59050(x59050, x71992, x59044);
  nand n59051(x59051, x25782, x85993);
  nand n59052(x59052, x59051, x59050);
  nand n59053(x59053, x25790, x85994);
  nand n59054(x59054, x71997, x59049);
  nand n59055(x59055, x25790, x59052);
  nand n59056(x59056, x59055, x59054);
  nand n59057(x59057, x72002, x85995);
  nand n59058(x59058, x25796, x59056);
  nand n59059(x59059, x59058, x59057);
  nand n59060(x59060, x71977, x49825);
  nand n59061(x59061, x16876, x58718);
  nand n59062(x59062, x59061, x26053);
  nand n59063(x59063, x71977, x85909);
  nand n59064(x59064, x16876, x85861);
  nand n59065(x59065, x71977, x50807);
  nand n59066(x59066, x16876, x50807);
  nand n59067(x59067, x59066, x59065);
  nand n59068(x59068, x71977, x57970);
  nand n59069(x59069, x16876, x57932);
  nand n59070(x59070, x59069, x59068);
  nand n59071(x59071, x71977, x51055);
  nand n59072(x59072, x59061, x59071);
  nand n59073(x59073, x16876, x50038);
  nand n59074(x59074, x59073, x59071);
  nand n59075(x59075, x71977, x57789);
  nand n59076(x59076, x25749, x85996);
  nand n59077(x59077, x71982, x59062);
  nand n59078(x59078, x25749, x85997);
  nand n59079(x59079, x59078, x59077);
  nand n59080(x59080, x71982, x85998);
  nand n59081(x59081, x25749, x59067);
  nand n59082(x59082, x59081, x59080);
  nand n59083(x59083, x71982, x59070);
  nand n59084(x59084, x25749, x59072);
  nand n59085(x59085, x59084, x59083);
  nand n59086(x59086, x71982, x85997);
  nand n59087(x59087, x25749, x85998);
  nand n59088(x59088, x59087, x59086);
  nand n59089(x59089, x71982, x59067);
  nand n59090(x59090, x25749, x59070);
  nand n59091(x59091, x59090, x59089);
  nand n59092(x59092, x71982, x59074);
  nand n59093(x59093, x25749, x85999);
  nand n59094(x59094, x59093, x59092);
  nand n59095(x59095, x71987, x86000);
  nand n59096(x59096, x25772, x59079);
  nand n59097(x59097, x59096, x26090);
  nand n59098(x59098, x71987, x59082);
  nand n59099(x59099, x25772, x59085);
  nand n59100(x59100, x59099, x59098);
  nand n59101(x59101, x71987, x59088);
  nand n59102(x59102, x25772, x59091);
  nand n59103(x59103, x59102, x59101);
  nand n59104(x59104, x71987, x59094);
  nand n59105(x59105, x25782, x86001);
  nand n59106(x59106, x71992, x59097);
  nand n59107(x59107, x25782, x59100);
  nand n59108(x59108, x59107, x59106);
  nand n59109(x59109, x71992, x59103);
  nand n59110(x59110, x25782, x86002);
  nand n59111(x59111, x59110, x59109);
  nand n59112(x59112, x25790, x86003);
  nand n59113(x59113, x71997, x59108);
  nand n59114(x59114, x25790, x59111);
  nand n59115(x59115, x59114, x59113);
  nand n59116(x59116, x72002, x86004);
  nand n59117(x59117, x25796, x59115);
  nand n59118(x59118, x59117, x59116);
  nand n59119(x59119, x71977, x49827);
  nand n59120(x59120, x16876, x58721);
  nand n59121(x59121, x59120, x26116);
  nand n59122(x59122, x71977, x85910);
  nand n59123(x59123, x16876, x57437);
  nand n59124(x59124, x71977, x50812);
  nand n59125(x59125, x16876, x50812);
  nand n59126(x59126, x59125, x59124);
  nand n59127(x59127, x71977, x57972);
  nand n59128(x59128, x16876, x57933);
  nand n59129(x59129, x59128, x59127);
  nand n59130(x59130, x71977, x51103);
  nand n59131(x59131, x59120, x59130);
  nand n59132(x59132, x16876, x50044);
  nand n59133(x59133, x59132, x59130);
  nand n59134(x59134, x71977, x57793);
  nand n59135(x59135, x25749, x86005);
  nand n59136(x59136, x71982, x59121);
  nand n59137(x59137, x25749, x86006);
  nand n59138(x59138, x59137, x59136);
  nand n59139(x59139, x71982, x86007);
  nand n59140(x59140, x25749, x59126);
  nand n59141(x59141, x59140, x59139);
  nand n59142(x59142, x71982, x59129);
  nand n59143(x59143, x25749, x59131);
  nand n59144(x59144, x59143, x59142);
  nand n59145(x59145, x71982, x86006);
  nand n59146(x59146, x25749, x86007);
  nand n59147(x59147, x59146, x59145);
  nand n59148(x59148, x71982, x59126);
  nand n59149(x59149, x25749, x59129);
  nand n59150(x59150, x59149, x59148);
  nand n59151(x59151, x71982, x59133);
  nand n59152(x59152, x25749, x86008);
  nand n59153(x59153, x59152, x59151);
  nand n59154(x59154, x71987, x86009);
  nand n59155(x59155, x25772, x59138);
  nand n59156(x59156, x59155, x26153);
  nand n59157(x59157, x71987, x59141);
  nand n59158(x59158, x25772, x59144);
  nand n59159(x59159, x59158, x59157);
  nand n59160(x59160, x71987, x59147);
  nand n59161(x59161, x25772, x59150);
  nand n59162(x59162, x59161, x59160);
  nand n59163(x59163, x71987, x59153);
  nand n59164(x59164, x25782, x86010);
  nand n59165(x59165, x71992, x59156);
  nand n59166(x59166, x25782, x59159);
  nand n59167(x59167, x59166, x59165);
  nand n59168(x59168, x71992, x59162);
  nand n59169(x59169, x25782, x86011);
  nand n59170(x59170, x59169, x59168);
  nand n59171(x59171, x25790, x86012);
  nand n59172(x59172, x71997, x59167);
  nand n59173(x59173, x25790, x59170);
  nand n59174(x59174, x59173, x59172);
  nand n59175(x59175, x72002, x86013);
  nand n59176(x59176, x25796, x59174);
  nand n59177(x59177, x59176, x59175);
  nand n59178(x59178, x71977, x49829);
  nand n59179(x59179, x16876, x58724);
  nand n59180(x59180, x59179, x26179);
  nand n59181(x59181, x71977, x85911);
  nand n59182(x59182, x16876, x57441);
  nand n59183(x59183, x71977, x50817);
  nand n59184(x59184, x16876, x50817);
  nand n59185(x59185, x59184, x59183);
  nand n59186(x59186, x71977, x57974);
  nand n59187(x59187, x16876, x57934);
  nand n59188(x59188, x59187, x59186);
  nand n59189(x59189, x71977, x51158);
  nand n59190(x59190, x59179, x59189);
  nand n59191(x59191, x16876, x50050);
  nand n59192(x59192, x59191, x59189);
  nand n59193(x59193, x71977, x57797);
  nand n59194(x59194, x25749, x86014);
  nand n59195(x59195, x71982, x59180);
  nand n59196(x59196, x25749, x86015);
  nand n59197(x59197, x59196, x59195);
  nand n59198(x59198, x71982, x86016);
  nand n59199(x59199, x25749, x59185);
  nand n59200(x59200, x59199, x59198);
  nand n59201(x59201, x71982, x59188);
  nand n59202(x59202, x25749, x59190);
  nand n59203(x59203, x59202, x59201);
  nand n59204(x59204, x71982, x86015);
  nand n59205(x59205, x25749, x86016);
  nand n59206(x59206, x59205, x59204);
  nand n59207(x59207, x71982, x59185);
  nand n59208(x59208, x25749, x59188);
  nand n59209(x59209, x59208, x59207);
  nand n59210(x59210, x71982, x59192);
  nand n59211(x59211, x25749, x86017);
  nand n59212(x59212, x59211, x59210);
  nand n59213(x59213, x71987, x86018);
  nand n59214(x59214, x25772, x59197);
  nand n59215(x59215, x59214, x26216);
  nand n59216(x59216, x71987, x59200);
  nand n59217(x59217, x25772, x59203);
  nand n59218(x59218, x59217, x59216);
  nand n59219(x59219, x71987, x59206);
  nand n59220(x59220, x25772, x59209);
  nand n59221(x59221, x59220, x59219);
  nand n59222(x59222, x71987, x59212);
  nand n59223(x59223, x25782, x86019);
  nand n59224(x59224, x71992, x59215);
  nand n59225(x59225, x25782, x59218);
  nand n59226(x59226, x59225, x59224);
  nand n59227(x59227, x71992, x59221);
  nand n59228(x59228, x25782, x86020);
  nand n59229(x59229, x59228, x59227);
  nand n59230(x59230, x25790, x86021);
  nand n59231(x59231, x71997, x59226);
  nand n59232(x59232, x25790, x59229);
  nand n59233(x59233, x59232, x59231);
  nand n59234(x59234, x72002, x86022);
  nand n59235(x59235, x25796, x59233);
  nand n59236(x59236, x59235, x59234);
  nand n59237(x59237, x71977, x49831);
  nand n59238(x59238, x16876, x58727);
  nand n59239(x59239, x59238, x26242);
  nand n59240(x59240, x71977, x85912);
  nand n59241(x59241, x16876, x57445);
  nand n59242(x59242, x71977, x50822);
  nand n59243(x59243, x16876, x50822);
  nand n59244(x59244, x59243, x59242);
  nand n59245(x59245, x71977, x57976);
  nand n59246(x59246, x16876, x57935);
  nand n59247(x59247, x59246, x59245);
  nand n59248(x59248, x71977, x51221);
  nand n59249(x59249, x59238, x59248);
  nand n59250(x59250, x16876, x50056);
  nand n59251(x59251, x59250, x59248);
  nand n59252(x59252, x71977, x57801);
  nand n59253(x59253, x25749, x86023);
  nand n59254(x59254, x71982, x59239);
  nand n59255(x59255, x25749, x86024);
  nand n59256(x59256, x59255, x59254);
  nand n59257(x59257, x71982, x86025);
  nand n59258(x59258, x25749, x59244);
  nand n59259(x59259, x59258, x59257);
  nand n59260(x59260, x71982, x59247);
  nand n59261(x59261, x25749, x59249);
  nand n59262(x59262, x59261, x59260);
  nand n59263(x59263, x71982, x86024);
  nand n59264(x59264, x25749, x86025);
  nand n59265(x59265, x59264, x59263);
  nand n59266(x59266, x71982, x59244);
  nand n59267(x59267, x25749, x59247);
  nand n59268(x59268, x59267, x59266);
  nand n59269(x59269, x71982, x59251);
  nand n59270(x59270, x25749, x86026);
  nand n59271(x59271, x59270, x59269);
  nand n59272(x59272, x71987, x86027);
  nand n59273(x59273, x25772, x59256);
  nand n59274(x59274, x59273, x26279);
  nand n59275(x59275, x71987, x59259);
  nand n59276(x59276, x25772, x59262);
  nand n59277(x59277, x59276, x59275);
  nand n59278(x59278, x71987, x59265);
  nand n59279(x59279, x25772, x59268);
  nand n59280(x59280, x59279, x59278);
  nand n59281(x59281, x71987, x59271);
  nand n59282(x59282, x25782, x86028);
  nand n59283(x59283, x71992, x59274);
  nand n59284(x59284, x25782, x59277);
  nand n59285(x59285, x59284, x59283);
  nand n59286(x59286, x71992, x59280);
  nand n59287(x59287, x25782, x86029);
  nand n59288(x59288, x59287, x59286);
  nand n59289(x59289, x25790, x86030);
  nand n59290(x59290, x71997, x59285);
  nand n59291(x59291, x25790, x59288);
  nand n59292(x59292, x59291, x59290);
  nand n59293(x59293, x72002, x86031);
  nand n59294(x59294, x25796, x59292);
  nand n59295(x59295, x59294, x59293);
  nand n59296(x59296, x71977, x49833);
  nand n59297(x59297, x16876, x58730);
  nand n59298(x59298, x59297, x26305);
  nand n59299(x59299, x71977, x85913);
  nand n59300(x59300, x16876, x57449);
  nand n59301(x59301, x71977, x50827);
  nand n59302(x59302, x16876, x50827);
  nand n59303(x59303, x59302, x59301);
  nand n59304(x59304, x71977, x57978);
  nand n59305(x59305, x16876, x57936);
  nand n59306(x59306, x59305, x59304);
  nand n59307(x59307, x71977, x51293);
  nand n59308(x59308, x59297, x59307);
  nand n59309(x59309, x16876, x50062);
  nand n59310(x59310, x59309, x59307);
  nand n59311(x59311, x71977, x57805);
  nand n59312(x59312, x25749, x86032);
  nand n59313(x59313, x71982, x59298);
  nand n59314(x59314, x25749, x86033);
  nand n59315(x59315, x59314, x59313);
  nand n59316(x59316, x71982, x86034);
  nand n59317(x59317, x25749, x59303);
  nand n59318(x59318, x59317, x59316);
  nand n59319(x59319, x71982, x59306);
  nand n59320(x59320, x25749, x59308);
  nand n59321(x59321, x59320, x59319);
  nand n59322(x59322, x71982, x86033);
  nand n59323(x59323, x25749, x86034);
  nand n59324(x59324, x59323, x59322);
  nand n59325(x59325, x71982, x59303);
  nand n59326(x59326, x25749, x59306);
  nand n59327(x59327, x59326, x59325);
  nand n59328(x59328, x71982, x59310);
  nand n59329(x59329, x25749, x86035);
  nand n59330(x59330, x59329, x59328);
  nand n59331(x59331, x71987, x86036);
  nand n59332(x59332, x25772, x59315);
  nand n59333(x59333, x59332, x26342);
  nand n59334(x59334, x71987, x59318);
  nand n59335(x59335, x25772, x59321);
  nand n59336(x59336, x59335, x59334);
  nand n59337(x59337, x71987, x59324);
  nand n59338(x59338, x25772, x59327);
  nand n59339(x59339, x59338, x59337);
  nand n59340(x59340, x71987, x59330);
  nand n59341(x59341, x25782, x86037);
  nand n59342(x59342, x71992, x59333);
  nand n59343(x59343, x25782, x59336);
  nand n59344(x59344, x59343, x59342);
  nand n59345(x59345, x71992, x59339);
  nand n59346(x59346, x25782, x86038);
  nand n59347(x59347, x59346, x59345);
  nand n59348(x59348, x25790, x86039);
  nand n59349(x59349, x71997, x59344);
  nand n59350(x59350, x25790, x59347);
  nand n59351(x59351, x59350, x59349);
  nand n59352(x59352, x72002, x86040);
  nand n59353(x59353, x25796, x59351);
  nand n59354(x59354, x59353, x59352);
  nand n59355(x59355, x71977, x49835);
  nand n59356(x59356, x16876, x58733);
  nand n59357(x59357, x59356, x26368);
  nand n59358(x59358, x71977, x85914);
  nand n59359(x59359, x16876, x57453);
  nand n59360(x59360, x71977, x50832);
  nand n59361(x59361, x16876, x50832);
  nand n59362(x59362, x59361, x59360);
  nand n59363(x59363, x71977, x57980);
  nand n59364(x59364, x16876, x57937);
  nand n59365(x59365, x59364, x59363);
  nand n59366(x59366, x71977, x51372);
  nand n59367(x59367, x59356, x59366);
  nand n59368(x59368, x16876, x50068);
  nand n59369(x59369, x59368, x59366);
  nand n59370(x59370, x71977, x57809);
  nand n59371(x59371, x25749, x86041);
  nand n59372(x59372, x71982, x59357);
  nand n59373(x59373, x25749, x86042);
  nand n59374(x59374, x59373, x59372);
  nand n59375(x59375, x71982, x86043);
  nand n59376(x59376, x25749, x59362);
  nand n59377(x59377, x59376, x59375);
  nand n59378(x59378, x71982, x59365);
  nand n59379(x59379, x25749, x59367);
  nand n59380(x59380, x59379, x59378);
  nand n59381(x59381, x71982, x86042);
  nand n59382(x59382, x25749, x86043);
  nand n59383(x59383, x59382, x59381);
  nand n59384(x59384, x71982, x59362);
  nand n59385(x59385, x25749, x59365);
  nand n59386(x59386, x59385, x59384);
  nand n59387(x59387, x71982, x59369);
  nand n59388(x59388, x25749, x86044);
  nand n59389(x59389, x59388, x59387);
  nand n59390(x59390, x71987, x86045);
  nand n59391(x59391, x25772, x59374);
  nand n59392(x59392, x59391, x26405);
  nand n59393(x59393, x71987, x59377);
  nand n59394(x59394, x25772, x59380);
  nand n59395(x59395, x59394, x59393);
  nand n59396(x59396, x71987, x59383);
  nand n59397(x59397, x25772, x59386);
  nand n59398(x59398, x59397, x59396);
  nand n59399(x59399, x71987, x59389);
  nand n59400(x59400, x25782, x86046);
  nand n59401(x59401, x71992, x59392);
  nand n59402(x59402, x25782, x59395);
  nand n59403(x59403, x59402, x59401);
  nand n59404(x59404, x71992, x59398);
  nand n59405(x59405, x25782, x86047);
  nand n59406(x59406, x59405, x59404);
  nand n59407(x59407, x25790, x86048);
  nand n59408(x59408, x71997, x59403);
  nand n59409(x59409, x25790, x59406);
  nand n59410(x59410, x59409, x59408);
  nand n59411(x59411, x72002, x86049);
  nand n59412(x59412, x25796, x59410);
  nand n59413(x59413, x59412, x59411);
  nand n59414(x59414, x71977, x49837);
  nand n59415(x59415, x16876, x58736);
  nand n59416(x59416, x59415, x26431);
  nand n59417(x59417, x71977, x85915);
  nand n59418(x59418, x16876, x57457);
  nand n59419(x59419, x71977, x50837);
  nand n59420(x59420, x16876, x50837);
  nand n59421(x59421, x59420, x59419);
  nand n59422(x59422, x71977, x57982);
  nand n59423(x59423, x16876, x57938);
  nand n59424(x59424, x59423, x59422);
  nand n59425(x59425, x71977, x51459);
  nand n59426(x59426, x59415, x59425);
  nand n59427(x59427, x16876, x50074);
  nand n59428(x59428, x59427, x59425);
  nand n59429(x59429, x71977, x57813);
  nand n59430(x59430, x25749, x86050);
  nand n59431(x59431, x71982, x59416);
  nand n59432(x59432, x25749, x86051);
  nand n59433(x59433, x59432, x59431);
  nand n59434(x59434, x71982, x86052);
  nand n59435(x59435, x25749, x59421);
  nand n59436(x59436, x59435, x59434);
  nand n59437(x59437, x71982, x59424);
  nand n59438(x59438, x25749, x59426);
  nand n59439(x59439, x59438, x59437);
  nand n59440(x59440, x71982, x86051);
  nand n59441(x59441, x25749, x86052);
  nand n59442(x59442, x59441, x59440);
  nand n59443(x59443, x71982, x59421);
  nand n59444(x59444, x25749, x59424);
  nand n59445(x59445, x59444, x59443);
  nand n59446(x59446, x71982, x59428);
  nand n59447(x59447, x25749, x86053);
  nand n59448(x59448, x59447, x59446);
  nand n59449(x59449, x71987, x86054);
  nand n59450(x59450, x25772, x59433);
  nand n59451(x59451, x59450, x26468);
  nand n59452(x59452, x71987, x59436);
  nand n59453(x59453, x25772, x59439);
  nand n59454(x59454, x59453, x59452);
  nand n59455(x59455, x71987, x59442);
  nand n59456(x59456, x25772, x59445);
  nand n59457(x59457, x59456, x59455);
  nand n59458(x59458, x71987, x59448);
  nand n59459(x59459, x25782, x86055);
  nand n59460(x59460, x71992, x59451);
  nand n59461(x59461, x25782, x59454);
  nand n59462(x59462, x59461, x59460);
  nand n59463(x59463, x71992, x59457);
  nand n59464(x59464, x25782, x86056);
  nand n59465(x59465, x59464, x59463);
  nand n59466(x59466, x25790, x86057);
  nand n59467(x59467, x71997, x59462);
  nand n59468(x59468, x25790, x59465);
  nand n59469(x59469, x59468, x59467);
  nand n59470(x59470, x72002, x86058);
  nand n59471(x59471, x25796, x59469);
  nand n59472(x59472, x59471, x59470);
  nand n59473(x59473, x71977, x49839);
  nand n59474(x59474, x16876, x58739);
  nand n59475(x59475, x59474, x26494);
  nand n59476(x59476, x71977, x85916);
  nand n59477(x59477, x16876, x57461);
  nand n59478(x59478, x71977, x50842);
  nand n59479(x59479, x16876, x50842);
  nand n59480(x59480, x59479, x59478);
  nand n59481(x59481, x71977, x57984);
  nand n59482(x59482, x16876, x57939);
  nand n59483(x59483, x59482, x59481);
  nand n59484(x59484, x71977, x51555);
  nand n59485(x59485, x59474, x59484);
  nand n59486(x59486, x16876, x50080);
  nand n59487(x59487, x59486, x59484);
  nand n59488(x59488, x71977, x57817);
  nand n59489(x59489, x25749, x86059);
  nand n59490(x59490, x71982, x59475);
  nand n59491(x59491, x25749, x86060);
  nand n59492(x59492, x59491, x59490);
  nand n59493(x59493, x71982, x86061);
  nand n59494(x59494, x25749, x59480);
  nand n59495(x59495, x59494, x59493);
  nand n59496(x59496, x71982, x59483);
  nand n59497(x59497, x25749, x59485);
  nand n59498(x59498, x59497, x59496);
  nand n59499(x59499, x71982, x86060);
  nand n59500(x59500, x25749, x86061);
  nand n59501(x59501, x59500, x59499);
  nand n59502(x59502, x71982, x59480);
  nand n59503(x59503, x25749, x59483);
  nand n59504(x59504, x59503, x59502);
  nand n59505(x59505, x71982, x59487);
  nand n59506(x59506, x25749, x86062);
  nand n59507(x59507, x59506, x59505);
  nand n59508(x59508, x71987, x86063);
  nand n59509(x59509, x25772, x59492);
  nand n59510(x59510, x59509, x26531);
  nand n59511(x59511, x71987, x59495);
  nand n59512(x59512, x25772, x59498);
  nand n59513(x59513, x59512, x59511);
  nand n59514(x59514, x71987, x59501);
  nand n59515(x59515, x25772, x59504);
  nand n59516(x59516, x59515, x59514);
  nand n59517(x59517, x71987, x59507);
  nand n59518(x59518, x25782, x86064);
  nand n59519(x59519, x71992, x59510);
  nand n59520(x59520, x25782, x59513);
  nand n59521(x59521, x59520, x59519);
  nand n59522(x59522, x71992, x59516);
  nand n59523(x59523, x25782, x86065);
  nand n59524(x59524, x59523, x59522);
  nand n59525(x59525, x25790, x86066);
  nand n59526(x59526, x71997, x59521);
  nand n59527(x59527, x25790, x59524);
  nand n59528(x59528, x59527, x59526);
  nand n59529(x59529, x72002, x86067);
  nand n59530(x59530, x25796, x59528);
  nand n59531(x59531, x59530, x59529);
  nand n59532(x59532, x71977, x49841);
  nand n59533(x59533, x16876, x58742);
  nand n59534(x59534, x59533, x26557);
  nand n59535(x59535, x71977, x85917);
  nand n59536(x59536, x16876, x57465);
  nand n59537(x59537, x71977, x50847);
  nand n59538(x59538, x16876, x50847);
  nand n59539(x59539, x59538, x59537);
  nand n59540(x59540, x71977, x57986);
  nand n59541(x59541, x16876, x57940);
  nand n59542(x59542, x59541, x59540);
  nand n59543(x59543, x71977, x51658);
  nand n59544(x59544, x59533, x59543);
  nand n59545(x59545, x16876, x50086);
  nand n59546(x59546, x59545, x59543);
  nand n59547(x59547, x71977, x57821);
  nand n59548(x59548, x25749, x86068);
  nand n59549(x59549, x71982, x59534);
  nand n59550(x59550, x25749, x86069);
  nand n59551(x59551, x59550, x59549);
  nand n59552(x59552, x71982, x86070);
  nand n59553(x59553, x25749, x59539);
  nand n59554(x59554, x59553, x59552);
  nand n59555(x59555, x71982, x59542);
  nand n59556(x59556, x25749, x59544);
  nand n59557(x59557, x59556, x59555);
  nand n59558(x59558, x71982, x86069);
  nand n59559(x59559, x25749, x86070);
  nand n59560(x59560, x59559, x59558);
  nand n59561(x59561, x71982, x59539);
  nand n59562(x59562, x25749, x59542);
  nand n59563(x59563, x59562, x59561);
  nand n59564(x59564, x71982, x59546);
  nand n59565(x59565, x25749, x86071);
  nand n59566(x59566, x59565, x59564);
  nand n59567(x59567, x71987, x86072);
  nand n59568(x59568, x25772, x59551);
  nand n59569(x59569, x59568, x26594);
  nand n59570(x59570, x71987, x59554);
  nand n59571(x59571, x25772, x59557);
  nand n59572(x59572, x59571, x59570);
  nand n59573(x59573, x71987, x59560);
  nand n59574(x59574, x25772, x59563);
  nand n59575(x59575, x59574, x59573);
  nand n59576(x59576, x71987, x59566);
  nand n59577(x59577, x25782, x86073);
  nand n59578(x59578, x71992, x59569);
  nand n59579(x59579, x25782, x59572);
  nand n59580(x59580, x59579, x59578);
  nand n59581(x59581, x71992, x59575);
  nand n59582(x59582, x25782, x86074);
  nand n59583(x59583, x59582, x59581);
  nand n59584(x59584, x25790, x86075);
  nand n59585(x59585, x71997, x59580);
  nand n59586(x59586, x25790, x59583);
  nand n59587(x59587, x59586, x59585);
  nand n59588(x59588, x72002, x86076);
  nand n59589(x59589, x25796, x59587);
  nand n59590(x59590, x59589, x59588);
  nand n59591(x59591, x71977, x49843);
  nand n59592(x59592, x16876, x58745);
  nand n59593(x59593, x59592, x26620);
  nand n59594(x59594, x71977, x85918);
  nand n59595(x59595, x16876, x57470);
  nand n59596(x59596, x71977, x50852);
  nand n59597(x59597, x16876, x50852);
  nand n59598(x59598, x59597, x59596);
  nand n59599(x59599, x71977, x57988);
  nand n59600(x59600, x16876, x57941);
  nand n59601(x59601, x59600, x59599);
  nand n59602(x59602, x71977, x51769);
  nand n59603(x59603, x59592, x59602);
  nand n59604(x59604, x16876, x50092);
  nand n59605(x59605, x59604, x59602);
  nand n59606(x59606, x71977, x57825);
  nand n59607(x59607, x25749, x86077);
  nand n59608(x59608, x71982, x59593);
  nand n59609(x59609, x25749, x86078);
  nand n59610(x59610, x59609, x59608);
  nand n59611(x59611, x71982, x86079);
  nand n59612(x59612, x25749, x59598);
  nand n59613(x59613, x59612, x59611);
  nand n59614(x59614, x71982, x59601);
  nand n59615(x59615, x25749, x59603);
  nand n59616(x59616, x59615, x59614);
  nand n59617(x59617, x71982, x86078);
  nand n59618(x59618, x25749, x86079);
  nand n59619(x59619, x59618, x59617);
  nand n59620(x59620, x71982, x59598);
  nand n59621(x59621, x25749, x59601);
  nand n59622(x59622, x59621, x59620);
  nand n59623(x59623, x71982, x59605);
  nand n59624(x59624, x25749, x86080);
  nand n59625(x59625, x59624, x59623);
  nand n59626(x59626, x71987, x86081);
  nand n59627(x59627, x25772, x59610);
  nand n59628(x59628, x59627, x26657);
  nand n59629(x59629, x71987, x59613);
  nand n59630(x59630, x25772, x59616);
  nand n59631(x59631, x59630, x59629);
  nand n59632(x59632, x71987, x59619);
  nand n59633(x59633, x25772, x59622);
  nand n59634(x59634, x59633, x59632);
  nand n59635(x59635, x71987, x59625);
  nand n59636(x59636, x25782, x86082);
  nand n59637(x59637, x71992, x59628);
  nand n59638(x59638, x25782, x59631);
  nand n59639(x59639, x59638, x59637);
  nand n59640(x59640, x71992, x59634);
  nand n59641(x59641, x25782, x86083);
  nand n59642(x59642, x59641, x59640);
  nand n59643(x59643, x25790, x86084);
  nand n59644(x59644, x71997, x59639);
  nand n59645(x59645, x25790, x59642);
  nand n59646(x59646, x59645, x59644);
  nand n59647(x59647, x72002, x86085);
  nand n59648(x59648, x25796, x59646);
  nand n59649(x59649, x59648, x59647);
  nand n59650(x59650, x71977, x49845);
  nand n59651(x59651, x16876, x58748);
  nand n59652(x59652, x59651, x26683);
  nand n59653(x59653, x71977, x85919);
  nand n59654(x59654, x16876, x57475);
  nand n59655(x59655, x71977, x50857);
  nand n59656(x59656, x16876, x50857);
  nand n59657(x59657, x59656, x59655);
  nand n59658(x59658, x71977, x57990);
  nand n59659(x59659, x16876, x57942);
  nand n59660(x59660, x59659, x59658);
  nand n59661(x59661, x71977, x51889);
  nand n59662(x59662, x59651, x59661);
  nand n59663(x59663, x16876, x50098);
  nand n59664(x59664, x59663, x59661);
  nand n59665(x59665, x71977, x57829);
  nand n59666(x59666, x25749, x86086);
  nand n59667(x59667, x71982, x59652);
  nand n59668(x59668, x25749, x86087);
  nand n59669(x59669, x59668, x59667);
  nand n59670(x59670, x71982, x86088);
  nand n59671(x59671, x25749, x59657);
  nand n59672(x59672, x59671, x59670);
  nand n59673(x59673, x71982, x59660);
  nand n59674(x59674, x25749, x59662);
  nand n59675(x59675, x59674, x59673);
  nand n59676(x59676, x71982, x86087);
  nand n59677(x59677, x25749, x86088);
  nand n59678(x59678, x59677, x59676);
  nand n59679(x59679, x71982, x59657);
  nand n59680(x59680, x25749, x59660);
  nand n59681(x59681, x59680, x59679);
  nand n59682(x59682, x71982, x59664);
  nand n59683(x59683, x25749, x86089);
  nand n59684(x59684, x59683, x59682);
  nand n59685(x59685, x71987, x86090);
  nand n59686(x59686, x25772, x59669);
  nand n59687(x59687, x59686, x26720);
  nand n59688(x59688, x71987, x59672);
  nand n59689(x59689, x25772, x59675);
  nand n59690(x59690, x59689, x59688);
  nand n59691(x59691, x71987, x59678);
  nand n59692(x59692, x25772, x59681);
  nand n59693(x59693, x59692, x59691);
  nand n59694(x59694, x71987, x59684);
  nand n59695(x59695, x25782, x86091);
  nand n59696(x59696, x71992, x59687);
  nand n59697(x59697, x25782, x59690);
  nand n59698(x59698, x59697, x59696);
  nand n59699(x59699, x71992, x59693);
  nand n59700(x59700, x25782, x86092);
  nand n59701(x59701, x59700, x59699);
  nand n59702(x59702, x25790, x86093);
  nand n59703(x59703, x71997, x59698);
  nand n59704(x59704, x25790, x59701);
  nand n59705(x59705, x59704, x59703);
  nand n59706(x59706, x72002, x86094);
  nand n59707(x59707, x25796, x59705);
  nand n59708(x59708, x59707, x59706);
  nand n59709(x59709, x71977, x49847);
  nand n59710(x59710, x16876, x85935);
  nand n59711(x59711, x59710, x26746);
  nand n59712(x59712, x71977, x58364);
  nand n59713(x59713, x16876, x57479);
  nand n59714(x59714, x71977, x50862);
  nand n59715(x59715, x16876, x50862);
  nand n59716(x59716, x59715, x59714);
  nand n59717(x59717, x71977, x57992);
  nand n59718(x59718, x16876, x57943);
  nand n59719(x59719, x59718, x59717);
  nand n59720(x59720, x71977, x57896);
  nand n59721(x59721, x59710, x59720);
  nand n59722(x59722, x16876, x50104);
  nand n59723(x59723, x59722, x59720);
  nand n59724(x59724, x71977, x57833);
  nand n59725(x59725, x25749, x86095);
  nand n59726(x59726, x71982, x59711);
  nand n59727(x59727, x25749, x86096);
  nand n59728(x59728, x59727, x59726);
  nand n59729(x59729, x71982, x86097);
  nand n59730(x59730, x25749, x59716);
  nand n59731(x59731, x59730, x59729);
  nand n59732(x59732, x71982, x59719);
  nand n59733(x59733, x25749, x59721);
  nand n59734(x59734, x59733, x59732);
  nand n59735(x59735, x71982, x86096);
  nand n59736(x59736, x25749, x86097);
  nand n59737(x59737, x59736, x59735);
  nand n59738(x59738, x71982, x59716);
  nand n59739(x59739, x25749, x59719);
  nand n59740(x59740, x59739, x59738);
  nand n59741(x59741, x71982, x59723);
  nand n59742(x59742, x25749, x86098);
  nand n59743(x59743, x59742, x59741);
  nand n59744(x59744, x71987, x86099);
  nand n59745(x59745, x25772, x59728);
  nand n59746(x59746, x59745, x26783);
  nand n59747(x59747, x71987, x59731);
  nand n59748(x59748, x25772, x59734);
  nand n59749(x59749, x59748, x59747);
  nand n59750(x59750, x71987, x59737);
  nand n59751(x59751, x25772, x59740);
  nand n59752(x59752, x59751, x59750);
  nand n59753(x59753, x71987, x59743);
  nand n59754(x59754, x25782, x86100);
  nand n59755(x59755, x71992, x59746);
  nand n59756(x59756, x25782, x59749);
  nand n59757(x59757, x59756, x59755);
  nand n59758(x59758, x71992, x59752);
  nand n59759(x59759, x25782, x86101);
  nand n59760(x59760, x59759, x59758);
  nand n59761(x59761, x25790, x86102);
  nand n59762(x59762, x71997, x59757);
  nand n59763(x59763, x25790, x59760);
  nand n59764(x59764, x59763, x59762);
  nand n59765(x59765, x72002, x86103);
  nand n59766(x59766, x25796, x59764);
  nand n59767(x59767, x59766, x59765);
  nand n59768(x59768, x71977, x49849);
  nand n59769(x59769, x16876, x85936);
  nand n59770(x59770, x59769, x26809);
  nand n59771(x59771, x71977, x58367);
  nand n59772(x59772, x16876, x57483);
  nand n59773(x59773, x71977, x50867);
  nand n59774(x59774, x16876, x50867);
  nand n59775(x59775, x59774, x59773);
  nand n59776(x59776, x71977, x57994);
  nand n59777(x59777, x16876, x57944);
  nand n59778(x59778, x59777, x59776);
  nand n59779(x59779, x71977, x57898);
  nand n59780(x59780, x59769, x59779);
  nand n59781(x59781, x16876, x50110);
  nand n59782(x59782, x59781, x59779);
  nand n59783(x59783, x71977, x57837);
  nand n59784(x59784, x25749, x86104);
  nand n59785(x59785, x71982, x59770);
  nand n59786(x59786, x25749, x86105);
  nand n59787(x59787, x59786, x59785);
  nand n59788(x59788, x71982, x86106);
  nand n59789(x59789, x25749, x59775);
  nand n59790(x59790, x59789, x59788);
  nand n59791(x59791, x71982, x59778);
  nand n59792(x59792, x25749, x59780);
  nand n59793(x59793, x59792, x59791);
  nand n59794(x59794, x71982, x86105);
  nand n59795(x59795, x25749, x86106);
  nand n59796(x59796, x59795, x59794);
  nand n59797(x59797, x71982, x59775);
  nand n59798(x59798, x25749, x59778);
  nand n59799(x59799, x59798, x59797);
  nand n59800(x59800, x71982, x59782);
  nand n59801(x59801, x25749, x86107);
  nand n59802(x59802, x59801, x59800);
  nand n59803(x59803, x71987, x86108);
  nand n59804(x59804, x25772, x59787);
  nand n59805(x59805, x59804, x26846);
  nand n59806(x59806, x71987, x59790);
  nand n59807(x59807, x25772, x59793);
  nand n59808(x59808, x59807, x59806);
  nand n59809(x59809, x71987, x59796);
  nand n59810(x59810, x25772, x59799);
  nand n59811(x59811, x59810, x59809);
  nand n59812(x59812, x71987, x59802);
  nand n59813(x59813, x25782, x86109);
  nand n59814(x59814, x71992, x59805);
  nand n59815(x59815, x25782, x59808);
  nand n59816(x59816, x59815, x59814);
  nand n59817(x59817, x71992, x59811);
  nand n59818(x59818, x25782, x86110);
  nand n59819(x59819, x59818, x59817);
  nand n59820(x59820, x25790, x86111);
  nand n59821(x59821, x71997, x59816);
  nand n59822(x59822, x25790, x59819);
  nand n59823(x59823, x59822, x59821);
  nand n59824(x59824, x72002, x86112);
  nand n59825(x59825, x25796, x59823);
  nand n59826(x59826, x59825, x59824);
  nand n59827(x59827, x71977, x49851);
  nand n59828(x59828, x16876, x85937);
  nand n59829(x59829, x59828, x26872);
  nand n59830(x59830, x71977, x58370);
  nand n59831(x59831, x16876, x57487);
  nand n59832(x59832, x71977, x50872);
  nand n59833(x59833, x16876, x50872);
  nand n59834(x59834, x59833, x59832);
  nand n59835(x59835, x71977, x57996);
  nand n59836(x59836, x16876, x57945);
  nand n59837(x59837, x59836, x59835);
  nand n59838(x59838, x71977, x57900);
  nand n59839(x59839, x59828, x59838);
  nand n59840(x59840, x16876, x50116);
  nand n59841(x59841, x59840, x59838);
  nand n59842(x59842, x71977, x57841);
  nand n59843(x59843, x25749, x86113);
  nand n59844(x59844, x71982, x59829);
  nand n59845(x59845, x25749, x86114);
  nand n59846(x59846, x59845, x59844);
  nand n59847(x59847, x71982, x86115);
  nand n59848(x59848, x25749, x59834);
  nand n59849(x59849, x59848, x59847);
  nand n59850(x59850, x71982, x59837);
  nand n59851(x59851, x25749, x59839);
  nand n59852(x59852, x59851, x59850);
  nand n59853(x59853, x71982, x86114);
  nand n59854(x59854, x25749, x86115);
  nand n59855(x59855, x59854, x59853);
  nand n59856(x59856, x71982, x59834);
  nand n59857(x59857, x25749, x59837);
  nand n59858(x59858, x59857, x59856);
  nand n59859(x59859, x71982, x59841);
  nand n59860(x59860, x25749, x86116);
  nand n59861(x59861, x59860, x59859);
  nand n59862(x59862, x71987, x86117);
  nand n59863(x59863, x25772, x59846);
  nand n59864(x59864, x59863, x26909);
  nand n59865(x59865, x71987, x59849);
  nand n59866(x59866, x25772, x59852);
  nand n59867(x59867, x59866, x59865);
  nand n59868(x59868, x71987, x59855);
  nand n59869(x59869, x25772, x59858);
  nand n59870(x59870, x59869, x59868);
  nand n59871(x59871, x71987, x59861);
  nand n59872(x59872, x25782, x86118);
  nand n59873(x59873, x71992, x59864);
  nand n59874(x59874, x25782, x59867);
  nand n59875(x59875, x59874, x59873);
  nand n59876(x59876, x71992, x59870);
  nand n59877(x59877, x25782, x86119);
  nand n59878(x59878, x59877, x59876);
  nand n59879(x59879, x25790, x86120);
  nand n59880(x59880, x71997, x59875);
  nand n59881(x59881, x25790, x59878);
  nand n59882(x59882, x59881, x59880);
  nand n59883(x59883, x72002, x86121);
  nand n59884(x59884, x25796, x59882);
  nand n59885(x59885, x59884, x59883);
  nand n59886(x59886, x71977, x49853);
  nand n59887(x59887, x16876, x85938);
  nand n59888(x59888, x59887, x26935);
  nand n59889(x59889, x71977, x58373);
  nand n59890(x59890, x16876, x57491);
  nand n59891(x59891, x71977, x50877);
  nand n59892(x59892, x16876, x50877);
  nand n59893(x59893, x59892, x59891);
  nand n59894(x59894, x71977, x57998);
  nand n59895(x59895, x16876, x57946);
  nand n59896(x59896, x59895, x59894);
  nand n59897(x59897, x71977, x57902);
  nand n59898(x59898, x59887, x59897);
  nand n59899(x59899, x16876, x50122);
  nand n59900(x59900, x59899, x59897);
  nand n59901(x59901, x71977, x57845);
  nand n59902(x59902, x25749, x86122);
  nand n59903(x59903, x71982, x59888);
  nand n59904(x59904, x25749, x86123);
  nand n59905(x59905, x59904, x59903);
  nand n59906(x59906, x71982, x86124);
  nand n59907(x59907, x25749, x59893);
  nand n59908(x59908, x59907, x59906);
  nand n59909(x59909, x71982, x59896);
  nand n59910(x59910, x25749, x59898);
  nand n59911(x59911, x59910, x59909);
  nand n59912(x59912, x71982, x86123);
  nand n59913(x59913, x25749, x86124);
  nand n59914(x59914, x59913, x59912);
  nand n59915(x59915, x71982, x59893);
  nand n59916(x59916, x25749, x59896);
  nand n59917(x59917, x59916, x59915);
  nand n59918(x59918, x71982, x59900);
  nand n59919(x59919, x25749, x86125);
  nand n59920(x59920, x59919, x59918);
  nand n59921(x59921, x71987, x86126);
  nand n59922(x59922, x25772, x59905);
  nand n59923(x59923, x59922, x26972);
  nand n59924(x59924, x71987, x59908);
  nand n59925(x59925, x25772, x59911);
  nand n59926(x59926, x59925, x59924);
  nand n59927(x59927, x71987, x59914);
  nand n59928(x59928, x25772, x59917);
  nand n59929(x59929, x59928, x59927);
  nand n59930(x59930, x71987, x59920);
  nand n59931(x59931, x25782, x86127);
  nand n59932(x59932, x71992, x59923);
  nand n59933(x59933, x25782, x59926);
  nand n59934(x59934, x59933, x59932);
  nand n59935(x59935, x71992, x59929);
  nand n59936(x59936, x25782, x86128);
  nand n59937(x59937, x59936, x59935);
  nand n59938(x59938, x25790, x86129);
  nand n59939(x59939, x71997, x59934);
  nand n59940(x59940, x25790, x59937);
  nand n59941(x59941, x59940, x59939);
  nand n59942(x59942, x72002, x86130);
  nand n59943(x59943, x25796, x59941);
  nand n59944(x59944, x59943, x59942);
  nand n59945(x59945, x71977, x49855);
  nand n59946(x59946, x16876, x85939);
  nand n59947(x59947, x59946, x26998);
  nand n59948(x59948, x71977, x58376);
  nand n59949(x59949, x16876, x57495);
  nand n59950(x59950, x71977, x50882);
  nand n59951(x59951, x16876, x50882);
  nand n59952(x59952, x59951, x59950);
  nand n59953(x59953, x71977, x58000);
  nand n59954(x59954, x16876, x57947);
  nand n59955(x59955, x59954, x59953);
  nand n59956(x59956, x71977, x57904);
  nand n59957(x59957, x59946, x59956);
  nand n59958(x59958, x16876, x50128);
  nand n59959(x59959, x59958, x59956);
  nand n59960(x59960, x71977, x57849);
  nand n59961(x59961, x25749, x86131);
  nand n59962(x59962, x71982, x59947);
  nand n59963(x59963, x25749, x86132);
  nand n59964(x59964, x59963, x59962);
  nand n59965(x59965, x71982, x86133);
  nand n59966(x59966, x25749, x59952);
  nand n59967(x59967, x59966, x59965);
  nand n59968(x59968, x71982, x59955);
  nand n59969(x59969, x25749, x59957);
  nand n59970(x59970, x59969, x59968);
  nand n59971(x59971, x71982, x86132);
  nand n59972(x59972, x25749, x86133);
  nand n59973(x59973, x59972, x59971);
  nand n59974(x59974, x71982, x59952);
  nand n59975(x59975, x25749, x59955);
  nand n59976(x59976, x59975, x59974);
  nand n59977(x59977, x71982, x59959);
  nand n59978(x59978, x25749, x86134);
  nand n59979(x59979, x59978, x59977);
  nand n59980(x59980, x71987, x86135);
  nand n59981(x59981, x25772, x59964);
  nand n59982(x59982, x59981, x27035);
  nand n59983(x59983, x71987, x59967);
  nand n59984(x59984, x25772, x59970);
  nand n59985(x59985, x59984, x59983);
  nand n59986(x59986, x71987, x59973);
  nand n59987(x59987, x25772, x59976);
  nand n59988(x59988, x59987, x59986);
  nand n59989(x59989, x71987, x59979);
  nand n59990(x59990, x25782, x86136);
  nand n59991(x59991, x71992, x59982);
  nand n59992(x59992, x25782, x59985);
  nand n59993(x59993, x59992, x59991);
  nand n59994(x59994, x71992, x59988);
  nand n59995(x59995, x25782, x86137);
  nand n59996(x59996, x59995, x59994);
  nand n59997(x59997, x25790, x86138);
  nand n59998(x59998, x71997, x59993);
  nand n59999(x59999, x25790, x59996);
  nand n60000(x60000, x59999, x59998);
  nand n60001(x60001, x72002, x86139);
  nand n60002(x60002, x25796, x60000);
  nand n60003(x60003, x60002, x60001);
  nand n60004(x60004, x71977, x49857);
  nand n60005(x60005, x16876, x85940);
  nand n60006(x60006, x60005, x27061);
  nand n60007(x60007, x71977, x58379);
  nand n60008(x60008, x16876, x57499);
  nand n60009(x60009, x71977, x50887);
  nand n60010(x60010, x16876, x50887);
  nand n60011(x60011, x60010, x60009);
  nand n60012(x60012, x71977, x58002);
  nand n60013(x60013, x16876, x57948);
  nand n60014(x60014, x60013, x60012);
  nand n60015(x60015, x71977, x57906);
  nand n60016(x60016, x60005, x60015);
  nand n60017(x60017, x16876, x50134);
  nand n60018(x60018, x60017, x60015);
  nand n60019(x60019, x71977, x57853);
  nand n60020(x60020, x25749, x86140);
  nand n60021(x60021, x71982, x60006);
  nand n60022(x60022, x25749, x86141);
  nand n60023(x60023, x60022, x60021);
  nand n60024(x60024, x71982, x86142);
  nand n60025(x60025, x25749, x60011);
  nand n60026(x60026, x60025, x60024);
  nand n60027(x60027, x71982, x60014);
  nand n60028(x60028, x25749, x60016);
  nand n60029(x60029, x60028, x60027);
  nand n60030(x60030, x71982, x86141);
  nand n60031(x60031, x25749, x86142);
  nand n60032(x60032, x60031, x60030);
  nand n60033(x60033, x71982, x60011);
  nand n60034(x60034, x25749, x60014);
  nand n60035(x60035, x60034, x60033);
  nand n60036(x60036, x71982, x60018);
  nand n60037(x60037, x25749, x86143);
  nand n60038(x60038, x60037, x60036);
  nand n60039(x60039, x71987, x86144);
  nand n60040(x60040, x25772, x60023);
  nand n60041(x60041, x60040, x27098);
  nand n60042(x60042, x71987, x60026);
  nand n60043(x60043, x25772, x60029);
  nand n60044(x60044, x60043, x60042);
  nand n60045(x60045, x71987, x60032);
  nand n60046(x60046, x25772, x60035);
  nand n60047(x60047, x60046, x60045);
  nand n60048(x60048, x71987, x60038);
  nand n60049(x60049, x25782, x86145);
  nand n60050(x60050, x71992, x60041);
  nand n60051(x60051, x25782, x60044);
  nand n60052(x60052, x60051, x60050);
  nand n60053(x60053, x71992, x60047);
  nand n60054(x60054, x25782, x86146);
  nand n60055(x60055, x60054, x60053);
  nand n60056(x60056, x25790, x86147);
  nand n60057(x60057, x71997, x60052);
  nand n60058(x60058, x25790, x60055);
  nand n60059(x60059, x60058, x60057);
  nand n60060(x60060, x72002, x86148);
  nand n60061(x60061, x25796, x60059);
  nand n60062(x60062, x60061, x60060);
  nand n60063(x60063, x71977, x49859);
  nand n60064(x60064, x16876, x85941);
  nand n60065(x60065, x60064, x27124);
  nand n60066(x60066, x71977, x58382);
  nand n60067(x60067, x16876, x57504);
  nand n60068(x60068, x71977, x50892);
  nand n60069(x60069, x16876, x50892);
  nand n60070(x60070, x60069, x60068);
  nand n60071(x60071, x71977, x58004);
  nand n60072(x60072, x16876, x57949);
  nand n60073(x60073, x60072, x60071);
  nand n60074(x60074, x71977, x57908);
  nand n60075(x60075, x60064, x60074);
  nand n60076(x60076, x16876, x50140);
  nand n60077(x60077, x60076, x60074);
  nand n60078(x60078, x71977, x57857);
  nand n60079(x60079, x25749, x86149);
  nand n60080(x60080, x71982, x60065);
  nand n60081(x60081, x25749, x86150);
  nand n60082(x60082, x60081, x60080);
  nand n60083(x60083, x71982, x86151);
  nand n60084(x60084, x25749, x60070);
  nand n60085(x60085, x60084, x60083);
  nand n60086(x60086, x71982, x60073);
  nand n60087(x60087, x25749, x60075);
  nand n60088(x60088, x60087, x60086);
  nand n60089(x60089, x71982, x86150);
  nand n60090(x60090, x25749, x86151);
  nand n60091(x60091, x60090, x60089);
  nand n60092(x60092, x71982, x60070);
  nand n60093(x60093, x25749, x60073);
  nand n60094(x60094, x60093, x60092);
  nand n60095(x60095, x71982, x60077);
  nand n60096(x60096, x25749, x86152);
  nand n60097(x60097, x60096, x60095);
  nand n60098(x60098, x71987, x86153);
  nand n60099(x60099, x25772, x60082);
  nand n60100(x60100, x60099, x27161);
  nand n60101(x60101, x71987, x60085);
  nand n60102(x60102, x25772, x60088);
  nand n60103(x60103, x60102, x60101);
  nand n60104(x60104, x71987, x60091);
  nand n60105(x60105, x25772, x60094);
  nand n60106(x60106, x60105, x60104);
  nand n60107(x60107, x71987, x60097);
  nand n60108(x60108, x25782, x86154);
  nand n60109(x60109, x71992, x60100);
  nand n60110(x60110, x25782, x60103);
  nand n60111(x60111, x60110, x60109);
  nand n60112(x60112, x71992, x60106);
  nand n60113(x60113, x25782, x86155);
  nand n60114(x60114, x60113, x60112);
  nand n60115(x60115, x25790, x86156);
  nand n60116(x60116, x71997, x60111);
  nand n60117(x60117, x25790, x60114);
  nand n60118(x60118, x60117, x60116);
  nand n60119(x60119, x72002, x86157);
  nand n60120(x60120, x25796, x60118);
  nand n60121(x60121, x60120, x60119);
  nand n60122(x60122, x71977, x49861);
  nand n60123(x60123, x16876, x85942);
  nand n60124(x60124, x60123, x27187);
  nand n60125(x60125, x71977, x58385);
  nand n60126(x60126, x16876, x57509);
  nand n60127(x60127, x71977, x50897);
  nand n60128(x60128, x16876, x50897);
  nand n60129(x60129, x60128, x60127);
  nand n60130(x60130, x71977, x58006);
  nand n60131(x60131, x16876, x57950);
  nand n60132(x60132, x60131, x60130);
  nand n60133(x60133, x71977, x57910);
  nand n60134(x60134, x60123, x60133);
  nand n60135(x60135, x16876, x50146);
  nand n60136(x60136, x60135, x60133);
  nand n60137(x60137, x71977, x57861);
  nand n60138(x60138, x25749, x86158);
  nand n60139(x60139, x71982, x60124);
  nand n60140(x60140, x25749, x86159);
  nand n60141(x60141, x60140, x60139);
  nand n60142(x60142, x71982, x86160);
  nand n60143(x60143, x25749, x60129);
  nand n60144(x60144, x60143, x60142);
  nand n60145(x60145, x71982, x60132);
  nand n60146(x60146, x25749, x60134);
  nand n60147(x60147, x60146, x60145);
  nand n60148(x60148, x71982, x86159);
  nand n60149(x60149, x25749, x86160);
  nand n60150(x60150, x60149, x60148);
  nand n60151(x60151, x71982, x60129);
  nand n60152(x60152, x25749, x60132);
  nand n60153(x60153, x60152, x60151);
  nand n60154(x60154, x71982, x60136);
  nand n60155(x60155, x25749, x86161);
  nand n60156(x60156, x60155, x60154);
  nand n60157(x60157, x71987, x86162);
  nand n60158(x60158, x25772, x60141);
  nand n60159(x60159, x60158, x27224);
  nand n60160(x60160, x71987, x60144);
  nand n60161(x60161, x25772, x60147);
  nand n60162(x60162, x60161, x60160);
  nand n60163(x60163, x71987, x60150);
  nand n60164(x60164, x25772, x60153);
  nand n60165(x60165, x60164, x60163);
  nand n60166(x60166, x71987, x60156);
  nand n60167(x60167, x25782, x86163);
  nand n60168(x60168, x71992, x60159);
  nand n60169(x60169, x25782, x60162);
  nand n60170(x60170, x60169, x60168);
  nand n60171(x60171, x71992, x60165);
  nand n60172(x60172, x25782, x86164);
  nand n60173(x60173, x60172, x60171);
  nand n60174(x60174, x25790, x86165);
  nand n60175(x60175, x71997, x60170);
  nand n60176(x60176, x25790, x60173);
  nand n60177(x60177, x60176, x60175);
  nand n60178(x60178, x72002, x86166);
  nand n60179(x60179, x25796, x60177);
  nand n60180(x60180, x60179, x60178);
  nand n60181(x60181, x71977, x49863);
  nand n60182(x60182, x16876, x85943);
  nand n60183(x60183, x60182, x27250);
  nand n60184(x60184, x71977, x58388);
  nand n60185(x60185, x16876, x57514);
  nand n60186(x60186, x71977, x50902);
  nand n60187(x60187, x16876, x50902);
  nand n60188(x60188, x60187, x60186);
  nand n60189(x60189, x71977, x58008);
  nand n60190(x60190, x16876, x57951);
  nand n60191(x60191, x60190, x60189);
  nand n60192(x60192, x71977, x57912);
  nand n60193(x60193, x60182, x60192);
  nand n60194(x60194, x16876, x50152);
  nand n60195(x60195, x60194, x60192);
  nand n60196(x60196, x71977, x57865);
  nand n60197(x60197, x25749, x86167);
  nand n60198(x60198, x71982, x60183);
  nand n60199(x60199, x25749, x86168);
  nand n60200(x60200, x60199, x60198);
  nand n60201(x60201, x71982, x86169);
  nand n60202(x60202, x25749, x60188);
  nand n60203(x60203, x60202, x60201);
  nand n60204(x60204, x71982, x60191);
  nand n60205(x60205, x25749, x60193);
  nand n60206(x60206, x60205, x60204);
  nand n60207(x60207, x71982, x86168);
  nand n60208(x60208, x25749, x86169);
  nand n60209(x60209, x60208, x60207);
  nand n60210(x60210, x71982, x60188);
  nand n60211(x60211, x25749, x60191);
  nand n60212(x60212, x60211, x60210);
  nand n60213(x60213, x71982, x60195);
  nand n60214(x60214, x25749, x86170);
  nand n60215(x60215, x60214, x60213);
  nand n60216(x60216, x71987, x86171);
  nand n60217(x60217, x25772, x60200);
  nand n60218(x60218, x60217, x27287);
  nand n60219(x60219, x71987, x60203);
  nand n60220(x60220, x25772, x60206);
  nand n60221(x60221, x60220, x60219);
  nand n60222(x60222, x71987, x60209);
  nand n60223(x60223, x25772, x60212);
  nand n60224(x60224, x60223, x60222);
  nand n60225(x60225, x71987, x60215);
  nand n60226(x60226, x25782, x86172);
  nand n60227(x60227, x71992, x60218);
  nand n60228(x60228, x25782, x60221);
  nand n60229(x60229, x60228, x60227);
  nand n60230(x60230, x71992, x60224);
  nand n60231(x60231, x25782, x86173);
  nand n60232(x60232, x60231, x60230);
  nand n60233(x60233, x25790, x86174);
  nand n60234(x60234, x71997, x60229);
  nand n60235(x60235, x25790, x60232);
  nand n60236(x60236, x60235, x60234);
  nand n60237(x60237, x72002, x86175);
  nand n60238(x60238, x25796, x60236);
  nand n60239(x60239, x60238, x60237);
  nand n60240(x60240, x71977, x49865);
  nand n60241(x60241, x16876, x85944);
  nand n60242(x60242, x60241, x27313);
  nand n60243(x60243, x71977, x58391);
  nand n60244(x60244, x16876, x57519);
  nand n60245(x60245, x71977, x50907);
  nand n60246(x60246, x16876, x50907);
  nand n60247(x60247, x60246, x60245);
  nand n60248(x60248, x71977, x58010);
  nand n60249(x60249, x16876, x57952);
  nand n60250(x60250, x60249, x60248);
  nand n60251(x60251, x71977, x57914);
  nand n60252(x60252, x60241, x60251);
  nand n60253(x60253, x16876, x50158);
  nand n60254(x60254, x60253, x60251);
  nand n60255(x60255, x71977, x57869);
  nand n60256(x60256, x25749, x86176);
  nand n60257(x60257, x71982, x60242);
  nand n60258(x60258, x25749, x86177);
  nand n60259(x60259, x60258, x60257);
  nand n60260(x60260, x71982, x86178);
  nand n60261(x60261, x25749, x60247);
  nand n60262(x60262, x60261, x60260);
  nand n60263(x60263, x71982, x60250);
  nand n60264(x60264, x25749, x60252);
  nand n60265(x60265, x60264, x60263);
  nand n60266(x60266, x71982, x86177);
  nand n60267(x60267, x25749, x86178);
  nand n60268(x60268, x60267, x60266);
  nand n60269(x60269, x71982, x60247);
  nand n60270(x60270, x25749, x60250);
  nand n60271(x60271, x60270, x60269);
  nand n60272(x60272, x71982, x60254);
  nand n60273(x60273, x25749, x86179);
  nand n60274(x60274, x60273, x60272);
  nand n60275(x60275, x71987, x86180);
  nand n60276(x60276, x25772, x60259);
  nand n60277(x60277, x60276, x27350);
  nand n60278(x60278, x71987, x60262);
  nand n60279(x60279, x25772, x60265);
  nand n60280(x60280, x60279, x60278);
  nand n60281(x60281, x71987, x60268);
  nand n60282(x60282, x25772, x60271);
  nand n60283(x60283, x60282, x60281);
  nand n60284(x60284, x71987, x60274);
  nand n60285(x60285, x25782, x86181);
  nand n60286(x60286, x71992, x60277);
  nand n60287(x60287, x25782, x60280);
  nand n60288(x60288, x60287, x60286);
  nand n60289(x60289, x71992, x60283);
  nand n60290(x60290, x25782, x86182);
  nand n60291(x60291, x60290, x60289);
  nand n60292(x60292, x25790, x86183);
  nand n60293(x60293, x71997, x60288);
  nand n60294(x60294, x25790, x60291);
  nand n60295(x60295, x60294, x60293);
  nand n60296(x60296, x72002, x86184);
  nand n60297(x60297, x25796, x60295);
  nand n60298(x60298, x60297, x60296);
  nand n60299(x60299, x71977, x49867);
  nand n60300(x60300, x16876, x85945);
  nand n60301(x60301, x60300, x27376);
  nand n60302(x60302, x71977, x58394);
  nand n60303(x60303, x16876, x57524);
  nand n60304(x60304, x71977, x50912);
  nand n60305(x60305, x16876, x50912);
  nand n60306(x60306, x60305, x60304);
  nand n60307(x60307, x71977, x58012);
  nand n60308(x60308, x16876, x57953);
  nand n60309(x60309, x60308, x60307);
  nand n60310(x60310, x71977, x57916);
  nand n60311(x60311, x60300, x60310);
  nand n60312(x60312, x16876, x50164);
  nand n60313(x60313, x60312, x60310);
  nand n60314(x60314, x71977, x57873);
  nand n60315(x60315, x25749, x86185);
  nand n60316(x60316, x71982, x60301);
  nand n60317(x60317, x25749, x86186);
  nand n60318(x60318, x60317, x60316);
  nand n60319(x60319, x71982, x86187);
  nand n60320(x60320, x25749, x60306);
  nand n60321(x60321, x60320, x60319);
  nand n60322(x60322, x71982, x60309);
  nand n60323(x60323, x25749, x60311);
  nand n60324(x60324, x60323, x60322);
  nand n60325(x60325, x71982, x86186);
  nand n60326(x60326, x25749, x86187);
  nand n60327(x60327, x60326, x60325);
  nand n60328(x60328, x71982, x60306);
  nand n60329(x60329, x25749, x60309);
  nand n60330(x60330, x60329, x60328);
  nand n60331(x60331, x71982, x60313);
  nand n60332(x60332, x25749, x86188);
  nand n60333(x60333, x60332, x60331);
  nand n60334(x60334, x71987, x86189);
  nand n60335(x60335, x25772, x60318);
  nand n60336(x60336, x60335, x27413);
  nand n60337(x60337, x71987, x60321);
  nand n60338(x60338, x25772, x60324);
  nand n60339(x60339, x60338, x60337);
  nand n60340(x60340, x71987, x60327);
  nand n60341(x60341, x25772, x60330);
  nand n60342(x60342, x60341, x60340);
  nand n60343(x60343, x71987, x60333);
  nand n60344(x60344, x25782, x86190);
  nand n60345(x60345, x71992, x60336);
  nand n60346(x60346, x25782, x60339);
  nand n60347(x60347, x60346, x60345);
  nand n60348(x60348, x71992, x60342);
  nand n60349(x60349, x25782, x86191);
  nand n60350(x60350, x60349, x60348);
  nand n60351(x60351, x25790, x86192);
  nand n60352(x60352, x71997, x60347);
  nand n60353(x60353, x25790, x60350);
  nand n60354(x60354, x60353, x60352);
  nand n60355(x60355, x72002, x86193);
  nand n60356(x60356, x25796, x60354);
  nand n60357(x60357, x60356, x60355);
  nand n60358(x60358, x71977, x49869);
  nand n60359(x60359, x16876, x85946);
  nand n60360(x60360, x60359, x27439);
  nand n60361(x60361, x71977, x58397);
  nand n60362(x60362, x16876, x57529);
  nand n60363(x60363, x71977, x50917);
  nand n60364(x60364, x16876, x50917);
  nand n60365(x60365, x60364, x60363);
  nand n60366(x60366, x71977, x58014);
  nand n60367(x60367, x16876, x57954);
  nand n60368(x60368, x60367, x60366);
  nand n60369(x60369, x71977, x57918);
  nand n60370(x60370, x60359, x60369);
  nand n60371(x60371, x16876, x50170);
  nand n60372(x60372, x60371, x60369);
  nand n60373(x60373, x71977, x57877);
  nand n60374(x60374, x25749, x86194);
  nand n60375(x60375, x71982, x60360);
  nand n60376(x60376, x25749, x86195);
  nand n60377(x60377, x60376, x60375);
  nand n60378(x60378, x71982, x86196);
  nand n60379(x60379, x25749, x60365);
  nand n60380(x60380, x60379, x60378);
  nand n60381(x60381, x71982, x60368);
  nand n60382(x60382, x25749, x60370);
  nand n60383(x60383, x60382, x60381);
  nand n60384(x60384, x71982, x86195);
  nand n60385(x60385, x25749, x86196);
  nand n60386(x60386, x60385, x60384);
  nand n60387(x60387, x71982, x60365);
  nand n60388(x60388, x25749, x60368);
  nand n60389(x60389, x60388, x60387);
  nand n60390(x60390, x71982, x60372);
  nand n60391(x60391, x25749, x86197);
  nand n60392(x60392, x60391, x60390);
  nand n60393(x60393, x71987, x86198);
  nand n60394(x60394, x25772, x60377);
  nand n60395(x60395, x60394, x27476);
  nand n60396(x60396, x71987, x60380);
  nand n60397(x60397, x25772, x60383);
  nand n60398(x60398, x60397, x60396);
  nand n60399(x60399, x71987, x60386);
  nand n60400(x60400, x25772, x60389);
  nand n60401(x60401, x60400, x60399);
  nand n60402(x60402, x71987, x60392);
  nand n60403(x60403, x25782, x86199);
  nand n60404(x60404, x71992, x60395);
  nand n60405(x60405, x25782, x60398);
  nand n60406(x60406, x60405, x60404);
  nand n60407(x60407, x71992, x60401);
  nand n60408(x60408, x25782, x86200);
  nand n60409(x60409, x60408, x60407);
  nand n60410(x60410, x25790, x86201);
  nand n60411(x60411, x71997, x60406);
  nand n60412(x60412, x25790, x60409);
  nand n60413(x60413, x60412, x60411);
  nand n60414(x60414, x72002, x86202);
  nand n60415(x60415, x25796, x60413);
  nand n60416(x60416, x60415, x60414);
  nand n60417(x60417, x71977, x49871);
  nand n60418(x60418, x16876, x85947);
  nand n60419(x60419, x60418, x27502);
  nand n60420(x60420, x71977, x58400);
  nand n60421(x60421, x16876, x57534);
  nand n60422(x60422, x71977, x50922);
  nand n60423(x60423, x16876, x50922);
  nand n60424(x60424, x60423, x60422);
  nand n60425(x60425, x71977, x58016);
  nand n60426(x60426, x16876, x57955);
  nand n60427(x60427, x60426, x60425);
  nand n60428(x60428, x71977, x57920);
  nand n60429(x60429, x60418, x60428);
  nand n60430(x60430, x16876, x50176);
  nand n60431(x60431, x60430, x60428);
  nand n60432(x60432, x71977, x57881);
  nand n60433(x60433, x25749, x86203);
  nand n60434(x60434, x71982, x60419);
  nand n60435(x60435, x25749, x86204);
  nand n60436(x60436, x60435, x60434);
  nand n60437(x60437, x71982, x86205);
  nand n60438(x60438, x25749, x60424);
  nand n60439(x60439, x60438, x60437);
  nand n60440(x60440, x71982, x60427);
  nand n60441(x60441, x25749, x60429);
  nand n60442(x60442, x60441, x60440);
  nand n60443(x60443, x71982, x86204);
  nand n60444(x60444, x25749, x86205);
  nand n60445(x60445, x60444, x60443);
  nand n60446(x60446, x71982, x60424);
  nand n60447(x60447, x25749, x60427);
  nand n60448(x60448, x60447, x60446);
  nand n60449(x60449, x71982, x60431);
  nand n60450(x60450, x25749, x86206);
  nand n60451(x60451, x60450, x60449);
  nand n60452(x60452, x71987, x86207);
  nand n60453(x60453, x25772, x60436);
  nand n60454(x60454, x60453, x27539);
  nand n60455(x60455, x71987, x60439);
  nand n60456(x60456, x25772, x60442);
  nand n60457(x60457, x60456, x60455);
  nand n60458(x60458, x71987, x60445);
  nand n60459(x60459, x25772, x60448);
  nand n60460(x60460, x60459, x60458);
  nand n60461(x60461, x71987, x60451);
  nand n60462(x60462, x25782, x86208);
  nand n60463(x60463, x71992, x60454);
  nand n60464(x60464, x25782, x60457);
  nand n60465(x60465, x60464, x60463);
  nand n60466(x60466, x71992, x60460);
  nand n60467(x60467, x25782, x86209);
  nand n60468(x60468, x60467, x60466);
  nand n60469(x60469, x25790, x86210);
  nand n60470(x60470, x71997, x60465);
  nand n60471(x60471, x25790, x60468);
  nand n60472(x60472, x60471, x60470);
  nand n60473(x60473, x72002, x86211);
  nand n60474(x60474, x25796, x60472);
  nand n60475(x60475, x60474, x60473);
  nand n60476(x60476, x71977, x49873);
  nand n60477(x60477, x16876, x85948);
  nand n60478(x60478, x60477, x27565);
  nand n60479(x60479, x71977, x58403);
  nand n60480(x60480, x16876, x57539);
  nand n60481(x60481, x71977, x50927);
  nand n60482(x60482, x16876, x50927);
  nand n60483(x60483, x60482, x60481);
  nand n60484(x60484, x71977, x58018);
  nand n60485(x60485, x16876, x57956);
  nand n60486(x60486, x60485, x60484);
  nand n60487(x60487, x71977, x57922);
  nand n60488(x60488, x60477, x60487);
  nand n60489(x60489, x16876, x50182);
  nand n60490(x60490, x60489, x60487);
  nand n60491(x60491, x71977, x57885);
  nand n60492(x60492, x25749, x86212);
  nand n60493(x60493, x71982, x60478);
  nand n60494(x60494, x25749, x86213);
  nand n60495(x60495, x60494, x60493);
  nand n60496(x60496, x71982, x86214);
  nand n60497(x60497, x25749, x60483);
  nand n60498(x60498, x60497, x60496);
  nand n60499(x60499, x71982, x60486);
  nand n60500(x60500, x25749, x60488);
  nand n60501(x60501, x60500, x60499);
  nand n60502(x60502, x71982, x86213);
  nand n60503(x60503, x25749, x86214);
  nand n60504(x60504, x60503, x60502);
  nand n60505(x60505, x71982, x60483);
  nand n60506(x60506, x25749, x60486);
  nand n60507(x60507, x60506, x60505);
  nand n60508(x60508, x71982, x60490);
  nand n60509(x60509, x25749, x86215);
  nand n60510(x60510, x60509, x60508);
  nand n60511(x60511, x71987, x86216);
  nand n60512(x60512, x25772, x60495);
  nand n60513(x60513, x60512, x27602);
  nand n60514(x60514, x71987, x60498);
  nand n60515(x60515, x25772, x60501);
  nand n60516(x60516, x60515, x60514);
  nand n60517(x60517, x71987, x60504);
  nand n60518(x60518, x25772, x60507);
  nand n60519(x60519, x60518, x60517);
  nand n60520(x60520, x71987, x60510);
  nand n60521(x60521, x25782, x86217);
  nand n60522(x60522, x71992, x60513);
  nand n60523(x60523, x25782, x60516);
  nand n60524(x60524, x60523, x60522);
  nand n60525(x60525, x71992, x60519);
  nand n60526(x60526, x25782, x86218);
  nand n60527(x60527, x60526, x60525);
  nand n60528(x60528, x25790, x86219);
  nand n60529(x60529, x71997, x60524);
  nand n60530(x60530, x25790, x60527);
  nand n60531(x60531, x60530, x60529);
  nand n60532(x60532, x72002, x86220);
  nand n60533(x60533, x25796, x60531);
  nand n60534(x60534, x60533, x60532);
  nand n60535(x60535, x71977, x49875);
  nand n60536(x60536, x16876, x85949);
  nand n60537(x60537, x60536, x27628);
  nand n60538(x60538, x71977, x58406);
  nand n60539(x60539, x16876, x57544);
  nand n60540(x60540, x71977, x50932);
  nand n60541(x60541, x16876, x50932);
  nand n60542(x60542, x60541, x60540);
  nand n60543(x60543, x71977, x58020);
  nand n60544(x60544, x16876, x57957);
  nand n60545(x60545, x60544, x60543);
  nand n60546(x60546, x71977, x57924);
  nand n60547(x60547, x60536, x60546);
  nand n60548(x60548, x16876, x50188);
  nand n60549(x60549, x60548, x60546);
  nand n60550(x60550, x71977, x57889);
  nand n60551(x60551, x25749, x86221);
  nand n60552(x60552, x71982, x60537);
  nand n60553(x60553, x25749, x86222);
  nand n60554(x60554, x60553, x60552);
  nand n60555(x60555, x71982, x86223);
  nand n60556(x60556, x25749, x60542);
  nand n60557(x60557, x60556, x60555);
  nand n60558(x60558, x71982, x60545);
  nand n60559(x60559, x25749, x60547);
  nand n60560(x60560, x60559, x60558);
  nand n60561(x60561, x71982, x86222);
  nand n60562(x60562, x25749, x86223);
  nand n60563(x60563, x60562, x60561);
  nand n60564(x60564, x71982, x60542);
  nand n60565(x60565, x25749, x60545);
  nand n60566(x60566, x60565, x60564);
  nand n60567(x60567, x71982, x60549);
  nand n60568(x60568, x25749, x86224);
  nand n60569(x60569, x60568, x60567);
  nand n60570(x60570, x71987, x86225);
  nand n60571(x60571, x25772, x60554);
  nand n60572(x60572, x60571, x27665);
  nand n60573(x60573, x71987, x60557);
  nand n60574(x60574, x25772, x60560);
  nand n60575(x60575, x60574, x60573);
  nand n60576(x60576, x71987, x60563);
  nand n60577(x60577, x25772, x60566);
  nand n60578(x60578, x60577, x60576);
  nand n60579(x60579, x71987, x60569);
  nand n60580(x60580, x25782, x86226);
  nand n60581(x60581, x71992, x60572);
  nand n60582(x60582, x25782, x60575);
  nand n60583(x60583, x60582, x60581);
  nand n60584(x60584, x71992, x60578);
  nand n60585(x60585, x25782, x86227);
  nand n60586(x60586, x60585, x60584);
  nand n60587(x60587, x25790, x86228);
  nand n60588(x60588, x71997, x60583);
  nand n60589(x60589, x25790, x60586);
  nand n60590(x60590, x60589, x60588);
  nand n60591(x60591, x72002, x86229);
  nand n60592(x60592, x25796, x60590);
  nand n60593(x60593, x60592, x60591);
  nand n60594(x60594, x71977, x49877);
  nand n60595(x60595, x16876, x85950);
  nand n60596(x60596, x60595, x27691);
  nand n60597(x60597, x71977, x58409);
  nand n60598(x60598, x16876, x57549);
  nand n60599(x60599, x71977, x50937);
  nand n60600(x60600, x16876, x50937);
  nand n60601(x60601, x60600, x60599);
  nand n60602(x60602, x71977, x58022);
  nand n60603(x60603, x16876, x57958);
  nand n60604(x60604, x60603, x60602);
  nand n60605(x60605, x71977, x57926);
  nand n60606(x60606, x60595, x60605);
  nand n60607(x60607, x16876, x50194);
  nand n60608(x60608, x60607, x60605);
  nand n60609(x60609, x71977, x57893);
  nand n60610(x60610, x25749, x86230);
  nand n60611(x60611, x71982, x60596);
  nand n60612(x60612, x25749, x86231);
  nand n60613(x60613, x60612, x60611);
  nand n60614(x60614, x71982, x86232);
  nand n60615(x60615, x25749, x60601);
  nand n60616(x60616, x60615, x60614);
  nand n60617(x60617, x71982, x60604);
  nand n60618(x60618, x25749, x60606);
  nand n60619(x60619, x60618, x60617);
  nand n60620(x60620, x71982, x86231);
  nand n60621(x60621, x25749, x86232);
  nand n60622(x60622, x60621, x60620);
  nand n60623(x60623, x71982, x60601);
  nand n60624(x60624, x25749, x60604);
  nand n60625(x60625, x60624, x60623);
  nand n60626(x60626, x71982, x60608);
  nand n60627(x60627, x25749, x86233);
  nand n60628(x60628, x60627, x60626);
  nand n60629(x60629, x71987, x86234);
  nand n60630(x60630, x25772, x60613);
  nand n60631(x60631, x60630, x27728);
  nand n60632(x60632, x71987, x60616);
  nand n60633(x60633, x25772, x60619);
  nand n60634(x60634, x60633, x60632);
  nand n60635(x60635, x71987, x60622);
  nand n60636(x60636, x25772, x60625);
  nand n60637(x60637, x60636, x60635);
  nand n60638(x60638, x71987, x60628);
  nand n60639(x60639, x25782, x86235);
  nand n60640(x60640, x71992, x60631);
  nand n60641(x60641, x25782, x60634);
  nand n60642(x60642, x60641, x60640);
  nand n60643(x60643, x71992, x60637);
  nand n60644(x60644, x25782, x86236);
  nand n60645(x60645, x60644, x60643);
  nand n60646(x60646, x25790, x86237);
  nand n60647(x60647, x71997, x60642);
  nand n60648(x60648, x25790, x60645);
  nand n60649(x60649, x60648, x60647);
  nand n60650(x60650, x72002, x86238);
  nand n60651(x60651, x25796, x60649);
  nand n60652(x60652, x60651, x60650);
  nand n60653(x60653, x16745, x58823);
  nand n60654(x60654, x68738, x60656);
  nand n60655(x60655, x60654, x60653);
  nand n60657(x60657, x16745, x58882);
  nand n60658(x60658, x68738, x60660);
  nand n60659(x60659, x60658, x60657);
  nand n60661(x60661, x16745, x58941);
  nand n60662(x60662, x68738, x60664);
  nand n60663(x60663, x60662, x60661);
  nand n60665(x60665, x16745, x59000);
  nand n60666(x60666, x68738, x60668);
  nand n60667(x60667, x60666, x60665);
  nand n60669(x60669, x16745, x59059);
  nand n60670(x60670, x68738, x60672);
  nand n60671(x60671, x60670, x60669);
  nand n60673(x60673, x16745, x59118);
  nand n60674(x60674, x68738, x60676);
  nand n60675(x60675, x60674, x60673);
  nand n60677(x60677, x16745, x59177);
  nand n60678(x60678, x68738, x60680);
  nand n60679(x60679, x60678, x60677);
  nand n60681(x60681, x16745, x59236);
  nand n60682(x60682, x68738, x60684);
  nand n60683(x60683, x60682, x60681);
  nand n60685(x60685, x16745, x59295);
  nand n60686(x60686, x68738, x60688);
  nand n60687(x60687, x60686, x60685);
  nand n60689(x60689, x16745, x59354);
  nand n60690(x60690, x68738, x60692);
  nand n60691(x60691, x60690, x60689);
  nand n60693(x60693, x16745, x59413);
  nand n60694(x60694, x68738, x60696);
  nand n60695(x60695, x60694, x60693);
  nand n60697(x60697, x16745, x59472);
  nand n60698(x60698, x68738, x60700);
  nand n60699(x60699, x60698, x60697);
  nand n60701(x60701, x16745, x59531);
  nand n60702(x60702, x68738, x60704);
  nand n60703(x60703, x60702, x60701);
  nand n60705(x60705, x16745, x59590);
  nand n60706(x60706, x68738, x60708);
  nand n60707(x60707, x60706, x60705);
  nand n60709(x60709, x16745, x59649);
  nand n60710(x60710, x68738, x60712);
  nand n60711(x60711, x60710, x60709);
  nand n60713(x60713, x16745, x59708);
  nand n60714(x60714, x68738, x60716);
  nand n60715(x60715, x60714, x60713);
  nand n60717(x60717, x16745, x59767);
  nand n60718(x60718, x68738, x60720);
  nand n60719(x60719, x60718, x60717);
  nand n60721(x60721, x16745, x59826);
  nand n60722(x60722, x68738, x60724);
  nand n60723(x60723, x60722, x60721);
  nand n60725(x60725, x16745, x59885);
  nand n60726(x60726, x68738, x60728);
  nand n60727(x60727, x60726, x60725);
  nand n60729(x60729, x16745, x59944);
  nand n60730(x60730, x68738, x60732);
  nand n60731(x60731, x60730, x60729);
  nand n60733(x60733, x16745, x60003);
  nand n60734(x60734, x68738, x60736);
  nand n60735(x60735, x60734, x60733);
  nand n60737(x60737, x16745, x60062);
  nand n60738(x60738, x68738, x60740);
  nand n60739(x60739, x60738, x60737);
  nand n60741(x60741, x16745, x60121);
  nand n60742(x60742, x68738, x60744);
  nand n60743(x60743, x60742, x60741);
  nand n60745(x60745, x16745, x60180);
  nand n60746(x60746, x68738, x60748);
  nand n60747(x60747, x60746, x60745);
  nand n60749(x60749, x16745, x60239);
  nand n60750(x60750, x68738, x60752);
  nand n60751(x60751, x60750, x60749);
  nand n60753(x60753, x16745, x60298);
  nand n60754(x60754, x68738, x60756);
  nand n60755(x60755, x60754, x60753);
  nand n60757(x60757, x16745, x60357);
  nand n60758(x60758, x68738, x60760);
  nand n60759(x60759, x60758, x60757);
  nand n60761(x60761, x16745, x60416);
  nand n60762(x60762, x68738, x60764);
  nand n60763(x60763, x60762, x60761);
  nand n60765(x60765, x16745, x60475);
  nand n60766(x60766, x68738, x60768);
  nand n60767(x60767, x60766, x60765);
  nand n60769(x60769, x16745, x60534);
  nand n60770(x60770, x68738, x60772);
  nand n60771(x60771, x60770, x60769);
  nand n60773(x60773, x16745, x60593);
  nand n60774(x60774, x68738, x60776);
  nand n60775(x60775, x60774, x60773);
  nand n60777(x60777, x16745, x60652);
  nand n60778(x60778, x68738, x60780);
  nand n60779(x60779, x60778, x60777);
  nand n60781(x60781, x16745, x83352);
  nand n60782(x60782, x68738, x60784);
  nand n60783(x60783, x60782, x60781);
  nand n60785(x60785, x16745, x71947);
  nand n60786(x60786, x68738, x60788);
  nand n60787(x60787, x60786, x60785);
  nand n60789(x60789, x16745, x71952);
  nand n60790(x60790, x68738, x60792);
  nand n60791(x60791, x60790, x60789);
  nand n60793(x60793, x16745, x71957);
  nand n60794(x60794, x68738, x60796);
  nand n60795(x60795, x60794, x60793);
  nand n60797(x60797, x16745, x71962);
  nand n60798(x60798, x68738, x60800);
  nand n60799(x60799, x60798, x60797);
  nand n60801(x60801, x16745, x71967);
  nand n60802(x60802, x68738, x60804);
  nand n60803(x60803, x60802, x60801);
  nand n60805(x60805, x16745, x71972);
  nand n60806(x60806, x68738, x60808);
  nand n60807(x60807, x60806, x60805);
  nand n60809(x60809, x16745, x72007);
  nand n60810(x60810, x68738, x60812);
  nand n60811(x60811, x60810, x60809);
  nand n60813(x60813, x16745, x72012);
  nand n60814(x60814, x68738, x60816);
  nand n60815(x60815, x60814, x60813);
  nand n60817(x60817, x16745, x72017);
  nand n60818(x60818, x68738, x60820);
  nand n60819(x60819, x60818, x60817);
  nand n60821(x60821, x16745, x72022);
  nand n60822(x60822, x68738, x60824);
  nand n60823(x60823, x60822, x60821);
  nand n60825(x60825, x16745, x72027);
  nand n60826(x60826, x68738, x60828);
  nand n60827(x60827, x60826, x60825);
  nand n60829(x60829, x16745, x72032);
  nand n60830(x60830, x68738, x60832);
  nand n60831(x60831, x60830, x60829);
  nand n60833(x60833, x16745, x72037);
  nand n60834(x60834, x68738, x60836);
  nand n60835(x60835, x60834, x60833);
  nand n60837(x60837, x16745, x72042);
  nand n60838(x60838, x68738, x60840);
  nand n60839(x60839, x60838, x60837);
  nand n60841(x60841, x68738, x83352);
  nand n60845(x60845, x60844, x60843);
  nand n60848(x60848, x60847, x60846);
  nand n60851(x60851, x60850, x60849);
  nand n60854(x60854, x60853, x60852);
  nand n60857(x60857, x60856, x60855);
  nand n60860(x60860, x60859, x60858);
  nand n60863(x60863, x60862, x60861);
  nand n60866(x60866, x60865, x60864);
  nand n60869(x60869, x60868, x60867);
  nand n60872(x60872, x60871, x60870);
  nand n60875(x60875, x60874, x60873);
  nand n60878(x60878, x60877, x60876);
  nand n60881(x60881, x60880, x60879);
  nand n60884(x60884, x60883, x60882);
  nand n60887(x60887, x60886, x60885);
  nand n60890(x60890, x60889, x60888);
  nand n60893(x60893, x60892, x60891);
  nand n60896(x60896, x60895, x60894);
  nand n60899(x60899, x60898, x60897);
  nand n60902(x60902, x60901, x60900);
  nand n60905(x60905, x60904, x60903);
  nand n60908(x60908, x60907, x60906);
  nand n60911(x60911, x60910, x60909);
  nand n60914(x60914, x60913, x60912);
  nand n60917(x60917, x60916, x60915);
  nand n60920(x60920, x60919, x60918);
  nand n60923(x60923, x60922, x60921);
  nand n60926(x60926, x60925, x60924);
  nand n60929(x60929, x60928, x60927);
  nand n60932(x60932, x60931, x60930);
  nand n60935(x60935, x60934, x60933);
  nand n60936(x60936, x74452, x74455);
  nand n60940(x60940, x60939, x60938);
  nand n60941(x60941, x60940, x60936);
  nand n60945(x60945, x60944, x60943);
  nand n60946(x60946, x74122, x74257);
  nand n60947(x60947, x60944, x60939);
  nand n60948(x60948, x60947, x60946);
  nand n60949(x60949, x74122, x60942);
  nand n60950(x60950, x60944, x60940);
  nand n60951(x60951, x60950, x60949);
  nand n60952(x60952, x74122, x60937);
  nand n60953(x60953, x60944, x60935);
  nand n60954(x60954, x60953, x60952);
  nand n60956(x60956, x60955, x86239);
  nand n60957(x60957, x74125, x60948);
  nand n60958(x60958, x60955, x60951);
  nand n60959(x60959, x60958, x60957);
  nand n60960(x60960, x74125, x60954);
  nand n60961(x60961, x74128, x86240);
  nand n60963(x60963, x60962, x60959);
  nand n60964(x60964, x60963, x60961);
  nand n60965(x60965, x74128, x86241);
  nand n60966(x60966, x74131, x60964);
  nand n60968(x60968, x60967, x86242);
  nand n60969(x60969, x60968, x60966);
  nand n60971(x60971, x60970, x60969);
  nand n60972(x60972, x74137, x86243);
  nand n60973(x60973, x60842, x86244);
  nand n60974(x60974, x68739, x60976);
  nand n60975(x60975, x60974, x60973);
  nand n60979(x60979, x60978, x60977);
  nand n60982(x60982, x60981, x60980);
  nand n60985(x60985, x60984, x60983);
  nand n60988(x60988, x60987, x60986);
  nand n60991(x60991, x60990, x60989);
  nand n60994(x60994, x60993, x60992);
  nand n60997(x60997, x60996, x60995);
  nand n61000(x61000, x60999, x60998);
  nand n61003(x61003, x61002, x61001);
  nand n61006(x61006, x61005, x61004);
  nand n61009(x61009, x61008, x61007);
  nand n61012(x61012, x61011, x61010);
  nand n61015(x61015, x61014, x61013);
  nand n61018(x61018, x61017, x61016);
  nand n61021(x61021, x61020, x61019);
  nand n61024(x61024, x61023, x61022);
  nand n61027(x61027, x61026, x61025);
  nand n61030(x61030, x61029, x61028);
  nand n61033(x61033, x61032, x61031);
  nand n61036(x61036, x61035, x61034);
  nand n61039(x61039, x61038, x61037);
  nand n61042(x61042, x61041, x61040);
  nand n61045(x61045, x61044, x61043);
  nand n61048(x61048, x61047, x61046);
  nand n61051(x61051, x61050, x61049);
  nand n61054(x61054, x61053, x61052);
  nand n61057(x61057, x61056, x61055);
  nand n61060(x61060, x61059, x61058);
  nand n61063(x61063, x61062, x61061);
  nand n61066(x61066, x61065, x61064);
  nand n61069(x61069, x61068, x61067);
  nand n61070(x61070, x74746, x74749);
  nand n61074(x61074, x61073, x61072);
  nand n61075(x61075, x61074, x61070);
  nand n61078(x61078, x60944, x61077);
  nand n61079(x61079, x74122, x74551);
  nand n61080(x61080, x60944, x61073);
  nand n61081(x61081, x61080, x61079);
  nand n61082(x61082, x74122, x61076);
  nand n61083(x61083, x60944, x61074);
  nand n61084(x61084, x61083, x61082);
  nand n61085(x61085, x74122, x61071);
  nand n61086(x61086, x60944, x61069);
  nand n61087(x61087, x61086, x61085);
  nand n61088(x61088, x60955, x86245);
  nand n61089(x61089, x74125, x61081);
  nand n61090(x61090, x60955, x61084);
  nand n61091(x61091, x61090, x61089);
  nand n61092(x61092, x74125, x61087);
  nand n61093(x61093, x74128, x86246);
  nand n61094(x61094, x60962, x61091);
  nand n61095(x61095, x61094, x61093);
  nand n61096(x61096, x74128, x86247);
  nand n61097(x61097, x74131, x61095);
  nand n61098(x61098, x60967, x86248);
  nand n61099(x61099, x61098, x61097);
  nand n61100(x61100, x60970, x61099);
  nand n61101(x61101, x74137, x86249);
  nand n61102(x61102, x60842, x86250);
  nand n61103(x61103, x68739, x61105);
  nand n61104(x61104, x61103, x61102);
  nand n61108(x61108, x61107, x61106);
  nand n61111(x61111, x61110, x61109);
  nand n61114(x61114, x61113, x61112);
  nand n61117(x61117, x61116, x61115);
  nand n61120(x61120, x61119, x61118);
  nand n61123(x61123, x61122, x61121);
  nand n61126(x61126, x61125, x61124);
  nand n61129(x61129, x61128, x61127);
  nand n61132(x61132, x61131, x61130);
  nand n61135(x61135, x61134, x61133);
  nand n61138(x61138, x61137, x61136);
  nand n61141(x61141, x61140, x61139);
  nand n61144(x61144, x61143, x61142);
  nand n61147(x61147, x61146, x61145);
  nand n61150(x61150, x61149, x61148);
  nand n61153(x61153, x61152, x61151);
  nand n61156(x61156, x61155, x61154);
  nand n61159(x61159, x61158, x61157);
  nand n61162(x61162, x61161, x61160);
  nand n61165(x61165, x61164, x61163);
  nand n61168(x61168, x61167, x61166);
  nand n61171(x61171, x61170, x61169);
  nand n61174(x61174, x61173, x61172);
  nand n61177(x61177, x61176, x61175);
  nand n61180(x61180, x61179, x61178);
  nand n61183(x61183, x61182, x61181);
  nand n61186(x61186, x61185, x61184);
  nand n61189(x61189, x61188, x61187);
  nand n61192(x61192, x61191, x61190);
  nand n61195(x61195, x61194, x61193);
  nand n61198(x61198, x61197, x61196);
  nand n61199(x61199, x75040, x75043);
  nand n61203(x61203, x61202, x61201);
  nand n61204(x61204, x61203, x61199);
  nand n61207(x61207, x60944, x61206);
  nand n61208(x61208, x74122, x74845);
  nand n61209(x61209, x60944, x61202);
  nand n61210(x61210, x61209, x61208);
  nand n61211(x61211, x74122, x61205);
  nand n61212(x61212, x60944, x61203);
  nand n61213(x61213, x61212, x61211);
  nand n61214(x61214, x74122, x61200);
  nand n61215(x61215, x60944, x61198);
  nand n61216(x61216, x61215, x61214);
  nand n61217(x61217, x60955, x86251);
  nand n61218(x61218, x74125, x61210);
  nand n61219(x61219, x60955, x61213);
  nand n61220(x61220, x61219, x61218);
  nand n61221(x61221, x74125, x61216);
  nand n61222(x61222, x74128, x86252);
  nand n61223(x61223, x60962, x61220);
  nand n61224(x61224, x61223, x61222);
  nand n61225(x61225, x74128, x86253);
  nand n61226(x61226, x74131, x61224);
  nand n61227(x61227, x60967, x86254);
  nand n61228(x61228, x61227, x61226);
  nand n61229(x61229, x60970, x61228);
  nand n61230(x61230, x74137, x86255);
  nand n61231(x61231, x60842, x86256);
  nand n61232(x61232, x68739, x61234);
  nand n61233(x61233, x61232, x61231);
  nand n61237(x61237, x61236, x61235);
  nand n61240(x61240, x61239, x61238);
  nand n61243(x61243, x61242, x61241);
  nand n61246(x61246, x61245, x61244);
  nand n61249(x61249, x61248, x61247);
  nand n61252(x61252, x61251, x61250);
  nand n61255(x61255, x61254, x61253);
  nand n61258(x61258, x61257, x61256);
  nand n61261(x61261, x61260, x61259);
  nand n61264(x61264, x61263, x61262);
  nand n61267(x61267, x61266, x61265);
  nand n61270(x61270, x61269, x61268);
  nand n61273(x61273, x61272, x61271);
  nand n61276(x61276, x61275, x61274);
  nand n61279(x61279, x61278, x61277);
  nand n61282(x61282, x61281, x61280);
  nand n61285(x61285, x61284, x61283);
  nand n61288(x61288, x61287, x61286);
  nand n61291(x61291, x61290, x61289);
  nand n61294(x61294, x61293, x61292);
  nand n61297(x61297, x61296, x61295);
  nand n61300(x61300, x61299, x61298);
  nand n61303(x61303, x61302, x61301);
  nand n61306(x61306, x61305, x61304);
  nand n61309(x61309, x61308, x61307);
  nand n61312(x61312, x61311, x61310);
  nand n61315(x61315, x61314, x61313);
  nand n61318(x61318, x61317, x61316);
  nand n61321(x61321, x61320, x61319);
  nand n61324(x61324, x61323, x61322);
  nand n61327(x61327, x61326, x61325);
  nand n61328(x61328, x75334, x75337);
  nand n61332(x61332, x61331, x61330);
  nand n61333(x61333, x61332, x61328);
  nand n61336(x61336, x60944, x61335);
  nand n61337(x61337, x74122, x75139);
  nand n61338(x61338, x60944, x61331);
  nand n61339(x61339, x61338, x61337);
  nand n61340(x61340, x74122, x61334);
  nand n61341(x61341, x60944, x61332);
  nand n61342(x61342, x61341, x61340);
  nand n61343(x61343, x74122, x61329);
  nand n61344(x61344, x60944, x61327);
  nand n61345(x61345, x61344, x61343);
  nand n61346(x61346, x60955, x86257);
  nand n61347(x61347, x74125, x61339);
  nand n61348(x61348, x60955, x61342);
  nand n61349(x61349, x61348, x61347);
  nand n61350(x61350, x74125, x61345);
  nand n61351(x61351, x74128, x86258);
  nand n61352(x61352, x60962, x61349);
  nand n61353(x61353, x61352, x61351);
  nand n61354(x61354, x74128, x86259);
  nand n61355(x61355, x74131, x61353);
  nand n61356(x61356, x60967, x86260);
  nand n61357(x61357, x61356, x61355);
  nand n61358(x61358, x60970, x61357);
  nand n61359(x61359, x74137, x86261);
  nand n61360(x61360, x60842, x86262);
  nand n61361(x61361, x68739, x61363);
  nand n61362(x61362, x61361, x61360);
  nand n61364(x61364, x60842, x83357);
  nand n61365(x61365, x68739, x61367);
  nand n61366(x61366, x61365, x61364);
  nand n61368(x61368, x60842, x74104);
  nand n61369(x61369, x68739, x61371);
  nand n61370(x61370, x61369, x61368);
  nand n61372(x61372, x60842, x74107);
  nand n61373(x61373, x68739, x61375);
  nand n61374(x61374, x61373, x61372);
  nand n61376(x61376, x60842, x74110);
  nand n61377(x61377, x68739, x61379);
  nand n61378(x61378, x61377, x61376);
  nand n61380(x61380, x60842, x74113);
  nand n61381(x61381, x68739, x61383);
  nand n61382(x61382, x61381, x61380);
  nand n61384(x61384, x60842, x74116);
  nand n61385(x61385, x68739, x61387);
  nand n61386(x61386, x61385, x61384);
  nand n61388(x61388, x60842, x74119);
  nand n61389(x61389, x68739, x61391);
  nand n61390(x61390, x61389, x61388);
  nand n61392(x61392, x60842, x74140);
  nand n61393(x61393, x68739, x61395);
  nand n61394(x61394, x61393, x61392);
  nand n61396(x61396, x60842, x74143);
  nand n61397(x61397, x68739, x61399);
  nand n61398(x61398, x61397, x61396);
  nand n61400(x61400, x60842, x74146);
  nand n61401(x61401, x68739, x61403);
  nand n61402(x61402, x61401, x61400);
  nand n61404(x61404, x60842, x74149);
  nand n61405(x61405, x68739, x61407);
  nand n61406(x61406, x61405, x61404);
  nand n61408(x61408, x60842, x74152);
  nand n61409(x61409, x68739, x61411);
  nand n61410(x61410, x61409, x61408);
  nand n61412(x61412, x60842, x74155);
  nand n61413(x61413, x68739, x61415);
  nand n61414(x61414, x61413, x61412);
  nand n61416(x61416, x60842, x74158);
  nand n61417(x61417, x68739, x61419);
  nand n61418(x61418, x61417, x61416);
  nand n61420(x61420, x60842, x74161);
  nand n61421(x61421, x68739, x61423);
  nand n61422(x61422, x61421, x61420);
  nand n61424(x61424, x68739, x83357);
  nand n61426(x61426, x61684, x61425);
  nand n61685(x61685, x75436, x75340);
  nand n61687(x61687, x61686, x75595);
  nand n61688(x61688, x61687, x61685);
  nand n61689(x61689, x75436, x75343);
  nand n61690(x61690, x61686, x75598);
  nand n61691(x61691, x61690, x61689);
  nand n61692(x61692, x75436, x75346);
  nand n61693(x61693, x61686, x75601);
  nand n61694(x61694, x61693, x61692);
  nand n61695(x61695, x75436, x75349);
  nand n61696(x61696, x61686, x75604);
  nand n61697(x61697, x61696, x61695);
  nand n61698(x61698, x75436, x75352);
  nand n61699(x61699, x61686, x75607);
  nand n61700(x61700, x61699, x61698);
  nand n61701(x61701, x75436, x75355);
  nand n61702(x61702, x61686, x75610);
  nand n61703(x61703, x61702, x61701);
  nand n61704(x61704, x75436, x75358);
  nand n61705(x61705, x61686, x75613);
  nand n61706(x61706, x61705, x61704);
  nand n61707(x61707, x75436, x75361);
  nand n61708(x61708, x61686, x75616);
  nand n61709(x61709, x61708, x61707);
  nand n61710(x61710, x75436, x75364);
  nand n61711(x61711, x61686, x75619);
  nand n61712(x61712, x61711, x61710);
  nand n61713(x61713, x75436, x75367);
  nand n61714(x61714, x61686, x75622);
  nand n61715(x61715, x61714, x61713);
  nand n61716(x61716, x75436, x75370);
  nand n61717(x61717, x61686, x75625);
  nand n61718(x61718, x61717, x61716);
  nand n61719(x61719, x75436, x75373);
  nand n61720(x61720, x61686, x75628);
  nand n61721(x61721, x61720, x61719);
  nand n61722(x61722, x75436, x75376);
  nand n61723(x61723, x61686, x75631);
  nand n61724(x61724, x61723, x61722);
  nand n61725(x61725, x75436, x75379);
  nand n61726(x61726, x61686, x75634);
  nand n61727(x61727, x61726, x61725);
  nand n61728(x61728, x75436, x75382);
  nand n61729(x61729, x61686, x75637);
  nand n61730(x61730, x61729, x61728);
  nand n61731(x61731, x75436, x75385);
  nand n61732(x61732, x61686, x75640);
  nand n61733(x61733, x61732, x61731);
  nand n61734(x61734, x75436, x75388);
  nand n61735(x61735, x61686, x75643);
  nand n61736(x61736, x61735, x61734);
  nand n61737(x61737, x75436, x75391);
  nand n61738(x61738, x61686, x75646);
  nand n61739(x61739, x61738, x61737);
  nand n61740(x61740, x75436, x75394);
  nand n61741(x61741, x61686, x75649);
  nand n61742(x61742, x61741, x61740);
  nand n61743(x61743, x75436, x75397);
  nand n61744(x61744, x61686, x75652);
  nand n61745(x61745, x61744, x61743);
  nand n61746(x61746, x75436, x75400);
  nand n61747(x61747, x61686, x75655);
  nand n61748(x61748, x61747, x61746);
  nand n61749(x61749, x75436, x75403);
  nand n61750(x61750, x61686, x75658);
  nand n61751(x61751, x61750, x61749);
  nand n61752(x61752, x75436, x75406);
  nand n61753(x61753, x61686, x75661);
  nand n61754(x61754, x61753, x61752);
  nand n61755(x61755, x75436, x75409);
  nand n61756(x61756, x61686, x75664);
  nand n61757(x61757, x61756, x61755);
  nand n61758(x61758, x75436, x75412);
  nand n61759(x61759, x61686, x75667);
  nand n61760(x61760, x61759, x61758);
  nand n61761(x61761, x75436, x75415);
  nand n61762(x61762, x61686, x75670);
  nand n61763(x61763, x61762, x61761);
  nand n61764(x61764, x75436, x75418);
  nand n61765(x61765, x61686, x75673);
  nand n61766(x61766, x61765, x61764);
  nand n61767(x61767, x75436, x75421);
  nand n61768(x61768, x61686, x75676);
  nand n61769(x61769, x61768, x61767);
  nand n61770(x61770, x75436, x75424);
  nand n61771(x61771, x61686, x75679);
  nand n61772(x61772, x61771, x61770);
  nand n61773(x61773, x75436, x75427);
  nand n61774(x61774, x61686, x75682);
  nand n61775(x61775, x61774, x61773);
  nand n61776(x61776, x75436, x75430);
  nand n61777(x61777, x61686, x75685);
  nand n61778(x61778, x61777, x61776);
  nand n61779(x61779, x75436, x75433);
  nand n61780(x61780, x61686, x75688);
  nand n61781(x61781, x61780, x61779);
  nand n61782(x61782, x61686, x75889);
  nand n61783(x61783, x61782, x61685);
  nand n61784(x61784, x61686, x75892);
  nand n61785(x61785, x61784, x61689);
  nand n61786(x61786, x61686, x75895);
  nand n61787(x61787, x61786, x61692);
  nand n61788(x61788, x61686, x75898);
  nand n61789(x61789, x61788, x61695);
  nand n61790(x61790, x61686, x75901);
  nand n61791(x61791, x61790, x61698);
  nand n61792(x61792, x61686, x75904);
  nand n61793(x61793, x61792, x61701);
  nand n61794(x61794, x61686, x75907);
  nand n61795(x61795, x61794, x61704);
  nand n61796(x61796, x61686, x75910);
  nand n61797(x61797, x61796, x61707);
  nand n61798(x61798, x61686, x75913);
  nand n61799(x61799, x61798, x61710);
  nand n61800(x61800, x61686, x75916);
  nand n61801(x61801, x61800, x61713);
  nand n61802(x61802, x61686, x75919);
  nand n61803(x61803, x61802, x61716);
  nand n61804(x61804, x61686, x75922);
  nand n61805(x61805, x61804, x61719);
  nand n61806(x61806, x61686, x75925);
  nand n61807(x61807, x61806, x61722);
  nand n61808(x61808, x61686, x75928);
  nand n61809(x61809, x61808, x61725);
  nand n61810(x61810, x61686, x75931);
  nand n61811(x61811, x61810, x61728);
  nand n61812(x61812, x61686, x75934);
  nand n61813(x61813, x61812, x61731);
  nand n61814(x61814, x61686, x75937);
  nand n61815(x61815, x61814, x61734);
  nand n61816(x61816, x61686, x75940);
  nand n61817(x61817, x61816, x61737);
  nand n61818(x61818, x61686, x75943);
  nand n61819(x61819, x61818, x61740);
  nand n61820(x61820, x61686, x75946);
  nand n61821(x61821, x61820, x61743);
  nand n61822(x61822, x61686, x75949);
  nand n61823(x61823, x61822, x61746);
  nand n61824(x61824, x61686, x75952);
  nand n61825(x61825, x61824, x61749);
  nand n61826(x61826, x61686, x75955);
  nand n61827(x61827, x61826, x61752);
  nand n61828(x61828, x61686, x75958);
  nand n61829(x61829, x61828, x61755);
  nand n61830(x61830, x61686, x75961);
  nand n61831(x61831, x61830, x61758);
  nand n61832(x61832, x61686, x75964);
  nand n61833(x61833, x61832, x61761);
  nand n61834(x61834, x61686, x75967);
  nand n61835(x61835, x61834, x61764);
  nand n61836(x61836, x61686, x75970);
  nand n61837(x61837, x61836, x61767);
  nand n61838(x61838, x61686, x75973);
  nand n61839(x61839, x61838, x61770);
  nand n61840(x61840, x61686, x75976);
  nand n61841(x61841, x61840, x61773);
  nand n61842(x61842, x61686, x75979);
  nand n61843(x61843, x61842, x61776);
  nand n61844(x61844, x61686, x75982);
  nand n61845(x61845, x61844, x61779);
  nand n61846(x61846, x61686, x76183);
  nand n61847(x61847, x61846, x61685);
  nand n61848(x61848, x61686, x76186);
  nand n61849(x61849, x61848, x61689);
  nand n61850(x61850, x61686, x76189);
  nand n61851(x61851, x61850, x61692);
  nand n61852(x61852, x61686, x76192);
  nand n61853(x61853, x61852, x61695);
  nand n61854(x61854, x61686, x76195);
  nand n61855(x61855, x61854, x61698);
  nand n61856(x61856, x61686, x76198);
  nand n61857(x61857, x61856, x61701);
  nand n61858(x61858, x61686, x76201);
  nand n61859(x61859, x61858, x61704);
  nand n61860(x61860, x61686, x76204);
  nand n61861(x61861, x61860, x61707);
  nand n61862(x61862, x61686, x76207);
  nand n61863(x61863, x61862, x61710);
  nand n61864(x61864, x61686, x76210);
  nand n61865(x61865, x61864, x61713);
  nand n61866(x61866, x61686, x76213);
  nand n61867(x61867, x61866, x61716);
  nand n61868(x61868, x61686, x76216);
  nand n61869(x61869, x61868, x61719);
  nand n61870(x61870, x61686, x76219);
  nand n61871(x61871, x61870, x61722);
  nand n61872(x61872, x61686, x76222);
  nand n61873(x61873, x61872, x61725);
  nand n61874(x61874, x61686, x76225);
  nand n61875(x61875, x61874, x61728);
  nand n61876(x61876, x61686, x76228);
  nand n61877(x61877, x61876, x61731);
  nand n61878(x61878, x61686, x76231);
  nand n61879(x61879, x61878, x61734);
  nand n61880(x61880, x61686, x76234);
  nand n61881(x61881, x61880, x61737);
  nand n61882(x61882, x61686, x76237);
  nand n61883(x61883, x61882, x61740);
  nand n61884(x61884, x61686, x76240);
  nand n61885(x61885, x61884, x61743);
  nand n61886(x61886, x61686, x76243);
  nand n61887(x61887, x61886, x61746);
  nand n61888(x61888, x61686, x76246);
  nand n61889(x61889, x61888, x61749);
  nand n61890(x61890, x61686, x76249);
  nand n61891(x61891, x61890, x61752);
  nand n61892(x61892, x61686, x76252);
  nand n61893(x61893, x61892, x61755);
  nand n61894(x61894, x61686, x76255);
  nand n61895(x61895, x61894, x61758);
  nand n61896(x61896, x61686, x76258);
  nand n61897(x61897, x61896, x61761);
  nand n61898(x61898, x61686, x76261);
  nand n61899(x61899, x61898, x61764);
  nand n61900(x61900, x61686, x76264);
  nand n61901(x61901, x61900, x61767);
  nand n61902(x61902, x61686, x76267);
  nand n61903(x61903, x61902, x61770);
  nand n61904(x61904, x61686, x76270);
  nand n61905(x61905, x61904, x61773);
  nand n61906(x61906, x61686, x76273);
  nand n61907(x61907, x61906, x61776);
  nand n61908(x61908, x61686, x76276);
  nand n61909(x61909, x61908, x61779);
  nand n61910(x61910, x61686, x76477);
  nand n61911(x61911, x61910, x61685);
  nand n61912(x61912, x61686, x76480);
  nand n61913(x61913, x61912, x61689);
  nand n61914(x61914, x61686, x76483);
  nand n61915(x61915, x61914, x61692);
  nand n61916(x61916, x61686, x76486);
  nand n61917(x61917, x61916, x61695);
  nand n61918(x61918, x61686, x76489);
  nand n61919(x61919, x61918, x61698);
  nand n61920(x61920, x61686, x76492);
  nand n61921(x61921, x61920, x61701);
  nand n61922(x61922, x61686, x76495);
  nand n61923(x61923, x61922, x61704);
  nand n61924(x61924, x61686, x76498);
  nand n61925(x61925, x61924, x61707);
  nand n61926(x61926, x61686, x76501);
  nand n61927(x61927, x61926, x61710);
  nand n61928(x61928, x61686, x76504);
  nand n61929(x61929, x61928, x61713);
  nand n61930(x61930, x61686, x76507);
  nand n61931(x61931, x61930, x61716);
  nand n61932(x61932, x61686, x76510);
  nand n61933(x61933, x61932, x61719);
  nand n61934(x61934, x61686, x76513);
  nand n61935(x61935, x61934, x61722);
  nand n61936(x61936, x61686, x76516);
  nand n61937(x61937, x61936, x61725);
  nand n61938(x61938, x61686, x76519);
  nand n61939(x61939, x61938, x61728);
  nand n61940(x61940, x61686, x76522);
  nand n61941(x61941, x61940, x61731);
  nand n61942(x61942, x61686, x76525);
  nand n61943(x61943, x61942, x61734);
  nand n61944(x61944, x61686, x76528);
  nand n61945(x61945, x61944, x61737);
  nand n61946(x61946, x61686, x76531);
  nand n61947(x61947, x61946, x61740);
  nand n61948(x61948, x61686, x76534);
  nand n61949(x61949, x61948, x61743);
  nand n61950(x61950, x61686, x76537);
  nand n61951(x61951, x61950, x61746);
  nand n61952(x61952, x61686, x76540);
  nand n61953(x61953, x61952, x61749);
  nand n61954(x61954, x61686, x76543);
  nand n61955(x61955, x61954, x61752);
  nand n61956(x61956, x61686, x76546);
  nand n61957(x61957, x61956, x61755);
  nand n61958(x61958, x61686, x76549);
  nand n61959(x61959, x61958, x61758);
  nand n61960(x61960, x61686, x76552);
  nand n61961(x61961, x61960, x61761);
  nand n61962(x61962, x61686, x76555);
  nand n61963(x61963, x61962, x61764);
  nand n61964(x61964, x61686, x76558);
  nand n61965(x61965, x61964, x61767);
  nand n61966(x61966, x61686, x76561);
  nand n61967(x61967, x61966, x61770);
  nand n61968(x61968, x61686, x76564);
  nand n61969(x61969, x61968, x61773);
  nand n61970(x61970, x61686, x76567);
  nand n61971(x61971, x61970, x61776);
  nand n61972(x61972, x61686, x76570);
  nand n61973(x61973, x61972, x61779);
  nand n61974(x61974, x75457, x61428);
  nand n61976(x61976, x61975, x61556);
  nand n61977(x61977, x61976, x61974);
  nand n61978(x61978, x61427, x61977);
  nand n61979(x61979, x61426, x61981);
  nand n61980(x61980, x61979, x61978);
  nand n61982(x61982, x75457, x61429);
  nand n61983(x61983, x61975, x61557);
  nand n61984(x61984, x61983, x61982);
  nand n61985(x61985, x61427, x61984);
  nand n61986(x61986, x61426, x61988);
  nand n61987(x61987, x61986, x61985);
  nand n61989(x61989, x75457, x61430);
  nand n61990(x61990, x61975, x61558);
  nand n61991(x61991, x61990, x61989);
  nand n61992(x61992, x61427, x61991);
  nand n61993(x61993, x61426, x61995);
  nand n61994(x61994, x61993, x61992);
  nand n61996(x61996, x75457, x61431);
  nand n61997(x61997, x61975, x61559);
  nand n61998(x61998, x61997, x61996);
  nand n61999(x61999, x61427, x61998);
  nand n62000(x62000, x61426, x62002);
  nand n62001(x62001, x62000, x61999);
  nand n62003(x62003, x75457, x61432);
  nand n62004(x62004, x61975, x61560);
  nand n62005(x62005, x62004, x62003);
  nand n62006(x62006, x61427, x62005);
  nand n62007(x62007, x61426, x62009);
  nand n62008(x62008, x62007, x62006);
  nand n62010(x62010, x75457, x61433);
  nand n62011(x62011, x61975, x61561);
  nand n62012(x62012, x62011, x62010);
  nand n62013(x62013, x61427, x62012);
  nand n62014(x62014, x61426, x62016);
  nand n62015(x62015, x62014, x62013);
  nand n62017(x62017, x75457, x61434);
  nand n62018(x62018, x61975, x61562);
  nand n62019(x62019, x62018, x62017);
  nand n62020(x62020, x61427, x62019);
  nand n62021(x62021, x61426, x62023);
  nand n62022(x62022, x62021, x62020);
  nand n62024(x62024, x75457, x61435);
  nand n62025(x62025, x61975, x61563);
  nand n62026(x62026, x62025, x62024);
  nand n62027(x62027, x61427, x62026);
  nand n62028(x62028, x61426, x62030);
  nand n62029(x62029, x62028, x62027);
  nand n62031(x62031, x75457, x61436);
  nand n62032(x62032, x61975, x61564);
  nand n62033(x62033, x62032, x62031);
  nand n62034(x62034, x61427, x62033);
  nand n62035(x62035, x61426, x62037);
  nand n62036(x62036, x62035, x62034);
  nand n62038(x62038, x75457, x61437);
  nand n62039(x62039, x61975, x61565);
  nand n62040(x62040, x62039, x62038);
  nand n62041(x62041, x61427, x62040);
  nand n62042(x62042, x61426, x62044);
  nand n62043(x62043, x62042, x62041);
  nand n62045(x62045, x75457, x61438);
  nand n62046(x62046, x61975, x61566);
  nand n62047(x62047, x62046, x62045);
  nand n62048(x62048, x61427, x62047);
  nand n62049(x62049, x61426, x62051);
  nand n62050(x62050, x62049, x62048);
  nand n62052(x62052, x75457, x61439);
  nand n62053(x62053, x61975, x61567);
  nand n62054(x62054, x62053, x62052);
  nand n62055(x62055, x61427, x62054);
  nand n62056(x62056, x61426, x62058);
  nand n62057(x62057, x62056, x62055);
  nand n62059(x62059, x75457, x61440);
  nand n62060(x62060, x61975, x61568);
  nand n62061(x62061, x62060, x62059);
  nand n62062(x62062, x61427, x62061);
  nand n62063(x62063, x61426, x62065);
  nand n62064(x62064, x62063, x62062);
  nand n62066(x62066, x75457, x61441);
  nand n62067(x62067, x61975, x61569);
  nand n62068(x62068, x62067, x62066);
  nand n62069(x62069, x61427, x62068);
  nand n62070(x62070, x61426, x62072);
  nand n62071(x62071, x62070, x62069);
  nand n62073(x62073, x75457, x61442);
  nand n62074(x62074, x61975, x61570);
  nand n62075(x62075, x62074, x62073);
  nand n62076(x62076, x61427, x62075);
  nand n62077(x62077, x61426, x62079);
  nand n62078(x62078, x62077, x62076);
  nand n62080(x62080, x75457, x61443);
  nand n62081(x62081, x61975, x61571);
  nand n62082(x62082, x62081, x62080);
  nand n62083(x62083, x61427, x62082);
  nand n62084(x62084, x61426, x62086);
  nand n62085(x62085, x62084, x62083);
  nand n62087(x62087, x75457, x61444);
  nand n62088(x62088, x61975, x61572);
  nand n62089(x62089, x62088, x62087);
  nand n62090(x62090, x61427, x62089);
  nand n62091(x62091, x61426, x62093);
  nand n62092(x62092, x62091, x62090);
  nand n62094(x62094, x75457, x61445);
  nand n62095(x62095, x61975, x61573);
  nand n62096(x62096, x62095, x62094);
  nand n62097(x62097, x61427, x62096);
  nand n62098(x62098, x61426, x62100);
  nand n62099(x62099, x62098, x62097);
  nand n62101(x62101, x75457, x61446);
  nand n62102(x62102, x61975, x61574);
  nand n62103(x62103, x62102, x62101);
  nand n62104(x62104, x61427, x62103);
  nand n62105(x62105, x61426, x62107);
  nand n62106(x62106, x62105, x62104);
  nand n62108(x62108, x75457, x61447);
  nand n62109(x62109, x61975, x61575);
  nand n62110(x62110, x62109, x62108);
  nand n62111(x62111, x61427, x62110);
  nand n62112(x62112, x61426, x62114);
  nand n62113(x62113, x62112, x62111);
  nand n62115(x62115, x75457, x61448);
  nand n62116(x62116, x61975, x61576);
  nand n62117(x62117, x62116, x62115);
  nand n62118(x62118, x61427, x62117);
  nand n62119(x62119, x61426, x62121);
  nand n62120(x62120, x62119, x62118);
  nand n62122(x62122, x75457, x61449);
  nand n62123(x62123, x61975, x61577);
  nand n62124(x62124, x62123, x62122);
  nand n62125(x62125, x61427, x62124);
  nand n62126(x62126, x61426, x62128);
  nand n62127(x62127, x62126, x62125);
  nand n62129(x62129, x75457, x61450);
  nand n62130(x62130, x61975, x61578);
  nand n62131(x62131, x62130, x62129);
  nand n62132(x62132, x61427, x62131);
  nand n62133(x62133, x61426, x62135);
  nand n62134(x62134, x62133, x62132);
  nand n62136(x62136, x75457, x61451);
  nand n62137(x62137, x61975, x61579);
  nand n62138(x62138, x62137, x62136);
  nand n62139(x62139, x61427, x62138);
  nand n62140(x62140, x61426, x62142);
  nand n62141(x62141, x62140, x62139);
  nand n62143(x62143, x75457, x61452);
  nand n62144(x62144, x61975, x61580);
  nand n62145(x62145, x62144, x62143);
  nand n62146(x62146, x61427, x62145);
  nand n62147(x62147, x61426, x62149);
  nand n62148(x62148, x62147, x62146);
  nand n62150(x62150, x75457, x61453);
  nand n62151(x62151, x61975, x61581);
  nand n62152(x62152, x62151, x62150);
  nand n62153(x62153, x61427, x62152);
  nand n62154(x62154, x61426, x62156);
  nand n62155(x62155, x62154, x62153);
  nand n62157(x62157, x75457, x61454);
  nand n62158(x62158, x61975, x61582);
  nand n62159(x62159, x62158, x62157);
  nand n62160(x62160, x61427, x62159);
  nand n62161(x62161, x61426, x62163);
  nand n62162(x62162, x62161, x62160);
  nand n62164(x62164, x75457, x61455);
  nand n62165(x62165, x61975, x61583);
  nand n62166(x62166, x62165, x62164);
  nand n62167(x62167, x61427, x62166);
  nand n62168(x62168, x61426, x62170);
  nand n62169(x62169, x62168, x62167);
  nand n62171(x62171, x75457, x61456);
  nand n62172(x62172, x61975, x61584);
  nand n62173(x62173, x62172, x62171);
  nand n62174(x62174, x61427, x62173);
  nand n62175(x62175, x61426, x62177);
  nand n62176(x62176, x62175, x62174);
  nand n62178(x62178, x75457, x61457);
  nand n62179(x62179, x61975, x61585);
  nand n62180(x62180, x62179, x62178);
  nand n62181(x62181, x61427, x62180);
  nand n62182(x62182, x61426, x62184);
  nand n62183(x62183, x62182, x62181);
  nand n62185(x62185, x75457, x61458);
  nand n62186(x62186, x61975, x61586);
  nand n62187(x62187, x62186, x62185);
  nand n62188(x62188, x61427, x62187);
  nand n62189(x62189, x61426, x62191);
  nand n62190(x62190, x62189, x62188);
  nand n62192(x62192, x75457, x61459);
  nand n62193(x62193, x61975, x61587);
  nand n62194(x62194, x62193, x62192);
  nand n62195(x62195, x61427, x62194);
  nand n62196(x62196, x61426, x62198);
  nand n62197(x62197, x62196, x62195);
  nand n62199(x62199, x75457, x61460);
  nand n62200(x62200, x61975, x61588);
  nand n62201(x62201, x62200, x62199);
  nand n62202(x62202, x61427, x62201);
  nand n62203(x62203, x61426, x62205);
  nand n62204(x62204, x62203, x62202);
  nand n62206(x62206, x75457, x61461);
  nand n62207(x62207, x61975, x61589);
  nand n62208(x62208, x62207, x62206);
  nand n62209(x62209, x61427, x62208);
  nand n62210(x62210, x61426, x62212);
  nand n62211(x62211, x62210, x62209);
  nand n62213(x62213, x75457, x61462);
  nand n62214(x62214, x61975, x61590);
  nand n62215(x62215, x62214, x62213);
  nand n62216(x62216, x61427, x62215);
  nand n62217(x62217, x61426, x62219);
  nand n62218(x62218, x62217, x62216);
  nand n62220(x62220, x75457, x61463);
  nand n62221(x62221, x61975, x61591);
  nand n62222(x62222, x62221, x62220);
  nand n62223(x62223, x61427, x62222);
  nand n62224(x62224, x61426, x62226);
  nand n62225(x62225, x62224, x62223);
  nand n62227(x62227, x75457, x61464);
  nand n62228(x62228, x61975, x61592);
  nand n62229(x62229, x62228, x62227);
  nand n62230(x62230, x61427, x62229);
  nand n62231(x62231, x61426, x62233);
  nand n62232(x62232, x62231, x62230);
  nand n62234(x62234, x75457, x61465);
  nand n62235(x62235, x61975, x61593);
  nand n62236(x62236, x62235, x62234);
  nand n62237(x62237, x61427, x62236);
  nand n62238(x62238, x61426, x62240);
  nand n62239(x62239, x62238, x62237);
  nand n62241(x62241, x75457, x61466);
  nand n62242(x62242, x61975, x61594);
  nand n62243(x62243, x62242, x62241);
  nand n62244(x62244, x61427, x62243);
  nand n62245(x62245, x61426, x62247);
  nand n62246(x62246, x62245, x62244);
  nand n62248(x62248, x75457, x61467);
  nand n62249(x62249, x61975, x61595);
  nand n62250(x62250, x62249, x62248);
  nand n62251(x62251, x61427, x62250);
  nand n62252(x62252, x61426, x62254);
  nand n62253(x62253, x62252, x62251);
  nand n62255(x62255, x75457, x61468);
  nand n62256(x62256, x61975, x61596);
  nand n62257(x62257, x62256, x62255);
  nand n62258(x62258, x61427, x62257);
  nand n62259(x62259, x61426, x62261);
  nand n62260(x62260, x62259, x62258);
  nand n62262(x62262, x75457, x61469);
  nand n62263(x62263, x61975, x61597);
  nand n62264(x62264, x62263, x62262);
  nand n62265(x62265, x61427, x62264);
  nand n62266(x62266, x61426, x62268);
  nand n62267(x62267, x62266, x62265);
  nand n62269(x62269, x75457, x61470);
  nand n62270(x62270, x61975, x61598);
  nand n62271(x62271, x62270, x62269);
  nand n62272(x62272, x61427, x62271);
  nand n62273(x62273, x61426, x62275);
  nand n62274(x62274, x62273, x62272);
  nand n62276(x62276, x75457, x61471);
  nand n62277(x62277, x61975, x61599);
  nand n62278(x62278, x62277, x62276);
  nand n62279(x62279, x61427, x62278);
  nand n62280(x62280, x61426, x62282);
  nand n62281(x62281, x62280, x62279);
  nand n62283(x62283, x75457, x61472);
  nand n62284(x62284, x61975, x61600);
  nand n62285(x62285, x62284, x62283);
  nand n62286(x62286, x61427, x62285);
  nand n62287(x62287, x61426, x62289);
  nand n62288(x62288, x62287, x62286);
  nand n62290(x62290, x75457, x61473);
  nand n62291(x62291, x61975, x61601);
  nand n62292(x62292, x62291, x62290);
  nand n62293(x62293, x61427, x62292);
  nand n62294(x62294, x61426, x62296);
  nand n62295(x62295, x62294, x62293);
  nand n62297(x62297, x75457, x61474);
  nand n62298(x62298, x61975, x61602);
  nand n62299(x62299, x62298, x62297);
  nand n62300(x62300, x61427, x62299);
  nand n62301(x62301, x61426, x62303);
  nand n62302(x62302, x62301, x62300);
  nand n62304(x62304, x75457, x61475);
  nand n62305(x62305, x61975, x61603);
  nand n62306(x62306, x62305, x62304);
  nand n62307(x62307, x61427, x62306);
  nand n62308(x62308, x61426, x62310);
  nand n62309(x62309, x62308, x62307);
  nand n62311(x62311, x75457, x61476);
  nand n62312(x62312, x61975, x61604);
  nand n62313(x62313, x62312, x62311);
  nand n62314(x62314, x61427, x62313);
  nand n62315(x62315, x61426, x62317);
  nand n62316(x62316, x62315, x62314);
  nand n62318(x62318, x75457, x61477);
  nand n62319(x62319, x61975, x61605);
  nand n62320(x62320, x62319, x62318);
  nand n62321(x62321, x61427, x62320);
  nand n62322(x62322, x61426, x62324);
  nand n62323(x62323, x62322, x62321);
  nand n62325(x62325, x75457, x61478);
  nand n62326(x62326, x61975, x61606);
  nand n62327(x62327, x62326, x62325);
  nand n62328(x62328, x61427, x62327);
  nand n62329(x62329, x61426, x62331);
  nand n62330(x62330, x62329, x62328);
  nand n62332(x62332, x75457, x61479);
  nand n62333(x62333, x61975, x61607);
  nand n62334(x62334, x62333, x62332);
  nand n62335(x62335, x61427, x62334);
  nand n62336(x62336, x61426, x62338);
  nand n62337(x62337, x62336, x62335);
  nand n62339(x62339, x75457, x61480);
  nand n62340(x62340, x61975, x61608);
  nand n62341(x62341, x62340, x62339);
  nand n62342(x62342, x61427, x62341);
  nand n62343(x62343, x61426, x62345);
  nand n62344(x62344, x62343, x62342);
  nand n62346(x62346, x75457, x61481);
  nand n62347(x62347, x61975, x61609);
  nand n62348(x62348, x62347, x62346);
  nand n62349(x62349, x61427, x62348);
  nand n62350(x62350, x61426, x62352);
  nand n62351(x62351, x62350, x62349);
  nand n62353(x62353, x75457, x61482);
  nand n62354(x62354, x61975, x61610);
  nand n62355(x62355, x62354, x62353);
  nand n62356(x62356, x61427, x62355);
  nand n62357(x62357, x61426, x62359);
  nand n62358(x62358, x62357, x62356);
  nand n62360(x62360, x75457, x61483);
  nand n62361(x62361, x61975, x61611);
  nand n62362(x62362, x62361, x62360);
  nand n62363(x62363, x61427, x62362);
  nand n62364(x62364, x61426, x62366);
  nand n62365(x62365, x62364, x62363);
  nand n62367(x62367, x75457, x61484);
  nand n62368(x62368, x61975, x61612);
  nand n62369(x62369, x62368, x62367);
  nand n62370(x62370, x61427, x62369);
  nand n62371(x62371, x61426, x62373);
  nand n62372(x62372, x62371, x62370);
  nand n62374(x62374, x75457, x61485);
  nand n62375(x62375, x61975, x61613);
  nand n62376(x62376, x62375, x62374);
  nand n62377(x62377, x61427, x62376);
  nand n62378(x62378, x61426, x62380);
  nand n62379(x62379, x62378, x62377);
  nand n62381(x62381, x75457, x61486);
  nand n62382(x62382, x61975, x61614);
  nand n62383(x62383, x62382, x62381);
  nand n62384(x62384, x61427, x62383);
  nand n62385(x62385, x61426, x62387);
  nand n62386(x62386, x62385, x62384);
  nand n62388(x62388, x75457, x61487);
  nand n62389(x62389, x61975, x61615);
  nand n62390(x62390, x62389, x62388);
  nand n62391(x62391, x61427, x62390);
  nand n62392(x62392, x61426, x62394);
  nand n62393(x62393, x62392, x62391);
  nand n62395(x62395, x75457, x61488);
  nand n62396(x62396, x61975, x61616);
  nand n62397(x62397, x62396, x62395);
  nand n62398(x62398, x61427, x62397);
  nand n62399(x62399, x61426, x62401);
  nand n62400(x62400, x62399, x62398);
  nand n62402(x62402, x75457, x61489);
  nand n62403(x62403, x61975, x61617);
  nand n62404(x62404, x62403, x62402);
  nand n62405(x62405, x61427, x62404);
  nand n62406(x62406, x61426, x62408);
  nand n62407(x62407, x62406, x62405);
  nand n62409(x62409, x75457, x61490);
  nand n62410(x62410, x61975, x61618);
  nand n62411(x62411, x62410, x62409);
  nand n62412(x62412, x61427, x62411);
  nand n62413(x62413, x61426, x62415);
  nand n62414(x62414, x62413, x62412);
  nand n62416(x62416, x75457, x61491);
  nand n62417(x62417, x61975, x61619);
  nand n62418(x62418, x62417, x62416);
  nand n62419(x62419, x61427, x62418);
  nand n62420(x62420, x61426, x62422);
  nand n62421(x62421, x62420, x62419);
  nand n62423(x62423, x75457, x61492);
  nand n62424(x62424, x61975, x61620);
  nand n62425(x62425, x62424, x62423);
  nand n62426(x62426, x61427, x62425);
  nand n62427(x62427, x61426, x62429);
  nand n62428(x62428, x62427, x62426);
  nand n62430(x62430, x75457, x61493);
  nand n62431(x62431, x61975, x61621);
  nand n62432(x62432, x62431, x62430);
  nand n62433(x62433, x61427, x62432);
  nand n62434(x62434, x61426, x62436);
  nand n62435(x62435, x62434, x62433);
  nand n62437(x62437, x75457, x61494);
  nand n62438(x62438, x61975, x61622);
  nand n62439(x62439, x62438, x62437);
  nand n62440(x62440, x61427, x62439);
  nand n62441(x62441, x61426, x62443);
  nand n62442(x62442, x62441, x62440);
  nand n62444(x62444, x75457, x61495);
  nand n62445(x62445, x61975, x61623);
  nand n62446(x62446, x62445, x62444);
  nand n62447(x62447, x61427, x62446);
  nand n62448(x62448, x61426, x62450);
  nand n62449(x62449, x62448, x62447);
  nand n62451(x62451, x75457, x61496);
  nand n62452(x62452, x61975, x61624);
  nand n62453(x62453, x62452, x62451);
  nand n62454(x62454, x61427, x62453);
  nand n62455(x62455, x61426, x62457);
  nand n62456(x62456, x62455, x62454);
  nand n62458(x62458, x75457, x61497);
  nand n62459(x62459, x61975, x61625);
  nand n62460(x62460, x62459, x62458);
  nand n62461(x62461, x61427, x62460);
  nand n62462(x62462, x61426, x62464);
  nand n62463(x62463, x62462, x62461);
  nand n62465(x62465, x75457, x61498);
  nand n62466(x62466, x61975, x61626);
  nand n62467(x62467, x62466, x62465);
  nand n62468(x62468, x61427, x62467);
  nand n62469(x62469, x61426, x62471);
  nand n62470(x62470, x62469, x62468);
  nand n62472(x62472, x75457, x61499);
  nand n62473(x62473, x61975, x61627);
  nand n62474(x62474, x62473, x62472);
  nand n62475(x62475, x61427, x62474);
  nand n62476(x62476, x61426, x62478);
  nand n62477(x62477, x62476, x62475);
  nand n62479(x62479, x75457, x61500);
  nand n62480(x62480, x61975, x61628);
  nand n62481(x62481, x62480, x62479);
  nand n62482(x62482, x61427, x62481);
  nand n62483(x62483, x61426, x62485);
  nand n62484(x62484, x62483, x62482);
  nand n62486(x62486, x75457, x61501);
  nand n62487(x62487, x61975, x61629);
  nand n62488(x62488, x62487, x62486);
  nand n62489(x62489, x61427, x62488);
  nand n62490(x62490, x61426, x62492);
  nand n62491(x62491, x62490, x62489);
  nand n62493(x62493, x75457, x61502);
  nand n62494(x62494, x61975, x61630);
  nand n62495(x62495, x62494, x62493);
  nand n62496(x62496, x61427, x62495);
  nand n62497(x62497, x61426, x62499);
  nand n62498(x62498, x62497, x62496);
  nand n62500(x62500, x75457, x61503);
  nand n62501(x62501, x61975, x61631);
  nand n62502(x62502, x62501, x62500);
  nand n62503(x62503, x61427, x62502);
  nand n62504(x62504, x61426, x62506);
  nand n62505(x62505, x62504, x62503);
  nand n62507(x62507, x75457, x61504);
  nand n62508(x62508, x61975, x61632);
  nand n62509(x62509, x62508, x62507);
  nand n62510(x62510, x61427, x62509);
  nand n62511(x62511, x61426, x62513);
  nand n62512(x62512, x62511, x62510);
  nand n62514(x62514, x75457, x61505);
  nand n62515(x62515, x61975, x61633);
  nand n62516(x62516, x62515, x62514);
  nand n62517(x62517, x61427, x62516);
  nand n62518(x62518, x61426, x62520);
  nand n62519(x62519, x62518, x62517);
  nand n62521(x62521, x75457, x61506);
  nand n62522(x62522, x61975, x61634);
  nand n62523(x62523, x62522, x62521);
  nand n62524(x62524, x61427, x62523);
  nand n62525(x62525, x61426, x62527);
  nand n62526(x62526, x62525, x62524);
  nand n62528(x62528, x75457, x61507);
  nand n62529(x62529, x61975, x61635);
  nand n62530(x62530, x62529, x62528);
  nand n62531(x62531, x61427, x62530);
  nand n62532(x62532, x61426, x62534);
  nand n62533(x62533, x62532, x62531);
  nand n62535(x62535, x75457, x61508);
  nand n62536(x62536, x61975, x61636);
  nand n62537(x62537, x62536, x62535);
  nand n62538(x62538, x61427, x62537);
  nand n62539(x62539, x61426, x62541);
  nand n62540(x62540, x62539, x62538);
  nand n62542(x62542, x75457, x61509);
  nand n62543(x62543, x61975, x61637);
  nand n62544(x62544, x62543, x62542);
  nand n62545(x62545, x61427, x62544);
  nand n62546(x62546, x61426, x62548);
  nand n62547(x62547, x62546, x62545);
  nand n62549(x62549, x75457, x61510);
  nand n62550(x62550, x61975, x61638);
  nand n62551(x62551, x62550, x62549);
  nand n62552(x62552, x61427, x62551);
  nand n62553(x62553, x61426, x62555);
  nand n62554(x62554, x62553, x62552);
  nand n62556(x62556, x75457, x61511);
  nand n62557(x62557, x61975, x61639);
  nand n62558(x62558, x62557, x62556);
  nand n62559(x62559, x61427, x62558);
  nand n62560(x62560, x61426, x62562);
  nand n62561(x62561, x62560, x62559);
  nand n62563(x62563, x75457, x61512);
  nand n62564(x62564, x61975, x61640);
  nand n62565(x62565, x62564, x62563);
  nand n62566(x62566, x61427, x62565);
  nand n62567(x62567, x61426, x62569);
  nand n62568(x62568, x62567, x62566);
  nand n62570(x62570, x75457, x61513);
  nand n62571(x62571, x61975, x61641);
  nand n62572(x62572, x62571, x62570);
  nand n62573(x62573, x61427, x62572);
  nand n62574(x62574, x61426, x62576);
  nand n62575(x62575, x62574, x62573);
  nand n62577(x62577, x75457, x61514);
  nand n62578(x62578, x61975, x61642);
  nand n62579(x62579, x62578, x62577);
  nand n62580(x62580, x61427, x62579);
  nand n62581(x62581, x61426, x62583);
  nand n62582(x62582, x62581, x62580);
  nand n62584(x62584, x75457, x61515);
  nand n62585(x62585, x61975, x61643);
  nand n62586(x62586, x62585, x62584);
  nand n62587(x62587, x61427, x62586);
  nand n62588(x62588, x61426, x62590);
  nand n62589(x62589, x62588, x62587);
  nand n62591(x62591, x75457, x61516);
  nand n62592(x62592, x61975, x61644);
  nand n62593(x62593, x62592, x62591);
  nand n62594(x62594, x61427, x62593);
  nand n62595(x62595, x61426, x62597);
  nand n62596(x62596, x62595, x62594);
  nand n62598(x62598, x75457, x61517);
  nand n62599(x62599, x61975, x61645);
  nand n62600(x62600, x62599, x62598);
  nand n62601(x62601, x61427, x62600);
  nand n62602(x62602, x61426, x62604);
  nand n62603(x62603, x62602, x62601);
  nand n62605(x62605, x75457, x61518);
  nand n62606(x62606, x61975, x61646);
  nand n62607(x62607, x62606, x62605);
  nand n62608(x62608, x61427, x62607);
  nand n62609(x62609, x61426, x62611);
  nand n62610(x62610, x62609, x62608);
  nand n62612(x62612, x75457, x61519);
  nand n62613(x62613, x61975, x61647);
  nand n62614(x62614, x62613, x62612);
  nand n62615(x62615, x61427, x62614);
  nand n62616(x62616, x61426, x62618);
  nand n62617(x62617, x62616, x62615);
  nand n62619(x62619, x75457, x61520);
  nand n62620(x62620, x61975, x61648);
  nand n62621(x62621, x62620, x62619);
  nand n62622(x62622, x61427, x62621);
  nand n62623(x62623, x61426, x62625);
  nand n62624(x62624, x62623, x62622);
  nand n62626(x62626, x75457, x61521);
  nand n62627(x62627, x61975, x61649);
  nand n62628(x62628, x62627, x62626);
  nand n62629(x62629, x61427, x62628);
  nand n62630(x62630, x61426, x62632);
  nand n62631(x62631, x62630, x62629);
  nand n62633(x62633, x75457, x61522);
  nand n62634(x62634, x61975, x61650);
  nand n62635(x62635, x62634, x62633);
  nand n62636(x62636, x61427, x62635);
  nand n62637(x62637, x61426, x62639);
  nand n62638(x62638, x62637, x62636);
  nand n62640(x62640, x75457, x61523);
  nand n62641(x62641, x61975, x61651);
  nand n62642(x62642, x62641, x62640);
  nand n62643(x62643, x61427, x62642);
  nand n62644(x62644, x61426, x62646);
  nand n62645(x62645, x62644, x62643);
  nand n62647(x62647, x75457, x61524);
  nand n62648(x62648, x61975, x61652);
  nand n62649(x62649, x62648, x62647);
  nand n62650(x62650, x61427, x62649);
  nand n62651(x62651, x61426, x62653);
  nand n62652(x62652, x62651, x62650);
  nand n62654(x62654, x75457, x61525);
  nand n62655(x62655, x61975, x61653);
  nand n62656(x62656, x62655, x62654);
  nand n62657(x62657, x61427, x62656);
  nand n62658(x62658, x61426, x62660);
  nand n62659(x62659, x62658, x62657);
  nand n62661(x62661, x75457, x61526);
  nand n62662(x62662, x61975, x61654);
  nand n62663(x62663, x62662, x62661);
  nand n62664(x62664, x61427, x62663);
  nand n62665(x62665, x61426, x62667);
  nand n62666(x62666, x62665, x62664);
  nand n62668(x62668, x75457, x61527);
  nand n62669(x62669, x61975, x61655);
  nand n62670(x62670, x62669, x62668);
  nand n62671(x62671, x61427, x62670);
  nand n62672(x62672, x61426, x62674);
  nand n62673(x62673, x62672, x62671);
  nand n62675(x62675, x75457, x61528);
  nand n62676(x62676, x61975, x61656);
  nand n62677(x62677, x62676, x62675);
  nand n62678(x62678, x61427, x62677);
  nand n62679(x62679, x61426, x62681);
  nand n62680(x62680, x62679, x62678);
  nand n62682(x62682, x75457, x61529);
  nand n62683(x62683, x61975, x61657);
  nand n62684(x62684, x62683, x62682);
  nand n62685(x62685, x61427, x62684);
  nand n62686(x62686, x61426, x62688);
  nand n62687(x62687, x62686, x62685);
  nand n62689(x62689, x75457, x61530);
  nand n62690(x62690, x61975, x61658);
  nand n62691(x62691, x62690, x62689);
  nand n62692(x62692, x61427, x62691);
  nand n62693(x62693, x61426, x62695);
  nand n62694(x62694, x62693, x62692);
  nand n62696(x62696, x75457, x61531);
  nand n62697(x62697, x61975, x61659);
  nand n62698(x62698, x62697, x62696);
  nand n62699(x62699, x61427, x62698);
  nand n62700(x62700, x61426, x62702);
  nand n62701(x62701, x62700, x62699);
  nand n62703(x62703, x75457, x61532);
  nand n62704(x62704, x61975, x61660);
  nand n62705(x62705, x62704, x62703);
  nand n62706(x62706, x61427, x62705);
  nand n62707(x62707, x61426, x62709);
  nand n62708(x62708, x62707, x62706);
  nand n62710(x62710, x75457, x61533);
  nand n62711(x62711, x61975, x61661);
  nand n62712(x62712, x62711, x62710);
  nand n62713(x62713, x61427, x62712);
  nand n62714(x62714, x61426, x62716);
  nand n62715(x62715, x62714, x62713);
  nand n62717(x62717, x75457, x61534);
  nand n62718(x62718, x61975, x61662);
  nand n62719(x62719, x62718, x62717);
  nand n62720(x62720, x61427, x62719);
  nand n62721(x62721, x61426, x62723);
  nand n62722(x62722, x62721, x62720);
  nand n62724(x62724, x75457, x61535);
  nand n62725(x62725, x61975, x61663);
  nand n62726(x62726, x62725, x62724);
  nand n62727(x62727, x61427, x62726);
  nand n62728(x62728, x61426, x62730);
  nand n62729(x62729, x62728, x62727);
  nand n62731(x62731, x75457, x61536);
  nand n62732(x62732, x61975, x61664);
  nand n62733(x62733, x62732, x62731);
  nand n62734(x62734, x61427, x62733);
  nand n62735(x62735, x61426, x62737);
  nand n62736(x62736, x62735, x62734);
  nand n62738(x62738, x75457, x61537);
  nand n62739(x62739, x61975, x61665);
  nand n62740(x62740, x62739, x62738);
  nand n62741(x62741, x61427, x62740);
  nand n62742(x62742, x61426, x62744);
  nand n62743(x62743, x62742, x62741);
  nand n62745(x62745, x75457, x61538);
  nand n62746(x62746, x61975, x61666);
  nand n62747(x62747, x62746, x62745);
  nand n62748(x62748, x61427, x62747);
  nand n62749(x62749, x61426, x62751);
  nand n62750(x62750, x62749, x62748);
  nand n62752(x62752, x75457, x61539);
  nand n62753(x62753, x61975, x61667);
  nand n62754(x62754, x62753, x62752);
  nand n62755(x62755, x61427, x62754);
  nand n62756(x62756, x61426, x62758);
  nand n62757(x62757, x62756, x62755);
  nand n62759(x62759, x75457, x61540);
  nand n62760(x62760, x61975, x61668);
  nand n62761(x62761, x62760, x62759);
  nand n62762(x62762, x61427, x62761);
  nand n62763(x62763, x61426, x62765);
  nand n62764(x62764, x62763, x62762);
  nand n62766(x62766, x75457, x61541);
  nand n62767(x62767, x61975, x61669);
  nand n62768(x62768, x62767, x62766);
  nand n62769(x62769, x61427, x62768);
  nand n62770(x62770, x61426, x62772);
  nand n62771(x62771, x62770, x62769);
  nand n62773(x62773, x75457, x61542);
  nand n62774(x62774, x61975, x61670);
  nand n62775(x62775, x62774, x62773);
  nand n62776(x62776, x61427, x62775);
  nand n62777(x62777, x61426, x62779);
  nand n62778(x62778, x62777, x62776);
  nand n62780(x62780, x75457, x61543);
  nand n62781(x62781, x61975, x61671);
  nand n62782(x62782, x62781, x62780);
  nand n62783(x62783, x61427, x62782);
  nand n62784(x62784, x61426, x62786);
  nand n62785(x62785, x62784, x62783);
  nand n62787(x62787, x75457, x61544);
  nand n62788(x62788, x61975, x61672);
  nand n62789(x62789, x62788, x62787);
  nand n62790(x62790, x61427, x62789);
  nand n62791(x62791, x61426, x62793);
  nand n62792(x62792, x62791, x62790);
  nand n62794(x62794, x75457, x61545);
  nand n62795(x62795, x61975, x61673);
  nand n62796(x62796, x62795, x62794);
  nand n62797(x62797, x61427, x62796);
  nand n62798(x62798, x61426, x62800);
  nand n62799(x62799, x62798, x62797);
  nand n62801(x62801, x75457, x61546);
  nand n62802(x62802, x61975, x61674);
  nand n62803(x62803, x62802, x62801);
  nand n62804(x62804, x61427, x62803);
  nand n62805(x62805, x61426, x62807);
  nand n62806(x62806, x62805, x62804);
  nand n62808(x62808, x75457, x61547);
  nand n62809(x62809, x61975, x61675);
  nand n62810(x62810, x62809, x62808);
  nand n62811(x62811, x61427, x62810);
  nand n62812(x62812, x61426, x62814);
  nand n62813(x62813, x62812, x62811);
  nand n62815(x62815, x75457, x61548);
  nand n62816(x62816, x61975, x61676);
  nand n62817(x62817, x62816, x62815);
  nand n62818(x62818, x61427, x62817);
  nand n62819(x62819, x61426, x62821);
  nand n62820(x62820, x62819, x62818);
  nand n62822(x62822, x75457, x61549);
  nand n62823(x62823, x61975, x61677);
  nand n62824(x62824, x62823, x62822);
  nand n62825(x62825, x61427, x62824);
  nand n62826(x62826, x61426, x62828);
  nand n62827(x62827, x62826, x62825);
  nand n62829(x62829, x75457, x61550);
  nand n62830(x62830, x61975, x61678);
  nand n62831(x62831, x62830, x62829);
  nand n62832(x62832, x61427, x62831);
  nand n62833(x62833, x61426, x62835);
  nand n62834(x62834, x62833, x62832);
  nand n62836(x62836, x75457, x61551);
  nand n62837(x62837, x61975, x61679);
  nand n62838(x62838, x62837, x62836);
  nand n62839(x62839, x61427, x62838);
  nand n62840(x62840, x61426, x62842);
  nand n62841(x62841, x62840, x62839);
  nand n62843(x62843, x75457, x61552);
  nand n62844(x62844, x61975, x61680);
  nand n62845(x62845, x62844, x62843);
  nand n62846(x62846, x61427, x62845);
  nand n62847(x62847, x61426, x62849);
  nand n62848(x62848, x62847, x62846);
  nand n62850(x62850, x75457, x61553);
  nand n62851(x62851, x61975, x61681);
  nand n62852(x62852, x62851, x62850);
  nand n62853(x62853, x61427, x62852);
  nand n62854(x62854, x61426, x62856);
  nand n62855(x62855, x62854, x62853);
  nand n62857(x62857, x75457, x61554);
  nand n62858(x62858, x61975, x61682);
  nand n62859(x62859, x62858, x62857);
  nand n62860(x62860, x61427, x62859);
  nand n62861(x62861, x61426, x62863);
  nand n62862(x62862, x62861, x62860);
  nand n62864(x62864, x75457, x61555);
  nand n62865(x62865, x61975, x61683);
  nand n62866(x62866, x62865, x62864);
  nand n62867(x62867, x61427, x62866);
  nand n62868(x62868, x61426, x62870);
  nand n62869(x62869, x62868, x62867);
  nand n62871(x62871, x83362, x61684);
  nand n62872(x62872, x61427, x83362);
  nand n62874(x62874, x61427, x75439);
  nand n62875(x62875, x61426, x62877);
  nand n62876(x62876, x62875, x62874);
  nand n62878(x62878, x61427, x75442);
  nand n62879(x62879, x61426, x62881);
  nand n62880(x62880, x62879, x62878);
  nand n62882(x62882, x61427, x75445);
  nand n62883(x62883, x61426, x62885);
  nand n62884(x62884, x62883, x62882);
  nand n62886(x62886, x61427, x75448);
  nand n62887(x62887, x61426, x62889);
  nand n62888(x62888, x62887, x62886);
  nand n62890(x62890, x61427, x75451);
  nand n62891(x62891, x61426, x62893);
  nand n62892(x62892, x62891, x62890);
  nand n62894(x62894, x61427, x75454);
  nand n62895(x62895, x61426, x62897);
  nand n62896(x62896, x62895, x62894);
  nand n62898(x62898, x61427, x75475);
  nand n62899(x62899, x61426, x62901);
  nand n62900(x62900, x62899, x62898);
  nand n62902(x62902, x61427, x75478);
  nand n62903(x62903, x61426, x62905);
  nand n62904(x62904, x62903, x62902);
  nand n62906(x62906, x61427, x75481);
  nand n62907(x62907, x61426, x62909);
  nand n62908(x62908, x62907, x62906);
  nand n62910(x62910, x61427, x75484);
  nand n62911(x62911, x61426, x62913);
  nand n62912(x62912, x62911, x62910);
  nand n62914(x62914, x61427, x75487);
  nand n62915(x62915, x61426, x62917);
  nand n62916(x62916, x62915, x62914);
  nand n62918(x62918, x61427, x75490);
  nand n62919(x62919, x61426, x62921);
  nand n62920(x62920, x62919, x62918);
  nand n62922(x62922, x61427, x75493);
  nand n62923(x62923, x61426, x62925);
  nand n62924(x62924, x62923, x62922);
  nand n62926(x62926, x61427, x75496);
  nand n62927(x62927, x61426, x62929);
  nand n62928(x62928, x62927, x62926);
  nand n62930(x62930, x62871, x83362);
  nand n62932(x62932, x76792, x76834);
  nand n62934(x62934, x62933, x76930);
  nand n62935(x62935, x62934, x62932);
  nand n62936(x62936, x76792, x76837);
  nand n62937(x62937, x62933, x76933);
  nand n62938(x62938, x62937, x62936);
  nand n62939(x62939, x76792, x76840);
  nand n62940(x62940, x62933, x76936);
  nand n62941(x62941, x62940, x62939);
  nand n62942(x62942, x76792, x76843);
  nand n62943(x62943, x62933, x76939);
  nand n62944(x62944, x62943, x62942);
  nand n62945(x62945, x76792, x76846);
  nand n62946(x62946, x62933, x76942);
  nand n62947(x62947, x62946, x62945);
  nand n62948(x62948, x76792, x76849);
  nand n62949(x62949, x62933, x76945);
  nand n62950(x62950, x62949, x62948);
  nand n62951(x62951, x76792, x76852);
  nand n62952(x62952, x62933, x76948);
  nand n62953(x62953, x62952, x62951);
  nand n62954(x62954, x76792, x76855);
  nand n62955(x62955, x62933, x76951);
  nand n62956(x62956, x62955, x62954);
  nand n62957(x62957, x76792, x76858);
  nand n62958(x62958, x62933, x76954);
  nand n62959(x62959, x62958, x62957);
  nand n62960(x62960, x76792, x76861);
  nand n62961(x62961, x62933, x76957);
  nand n62962(x62962, x62961, x62960);
  nand n62963(x62963, x76792, x76864);
  nand n62964(x62964, x62933, x76960);
  nand n62965(x62965, x62964, x62963);
  nand n62966(x62966, x76792, x76867);
  nand n62967(x62967, x62933, x76963);
  nand n62968(x62968, x62967, x62966);
  nand n62969(x62969, x76792, x76870);
  nand n62970(x62970, x62933, x76966);
  nand n62971(x62971, x62970, x62969);
  nand n62972(x62972, x76792, x76873);
  nand n62973(x62973, x62933, x76969);
  nand n62974(x62974, x62973, x62972);
  nand n62975(x62975, x76792, x76876);
  nand n62976(x62976, x62933, x76972);
  nand n62977(x62977, x62976, x62975);
  nand n62978(x62978, x76792, x76879);
  nand n62979(x62979, x62933, x76975);
  nand n62980(x62980, x62979, x62978);
  nand n62981(x62981, x76792, x76882);
  nand n62982(x62982, x62933, x76978);
  nand n62983(x62983, x62982, x62981);
  nand n62984(x62984, x76792, x76885);
  nand n62985(x62985, x62933, x76981);
  nand n62986(x62986, x62985, x62984);
  nand n62987(x62987, x76792, x76888);
  nand n62988(x62988, x62933, x76984);
  nand n62989(x62989, x62988, x62987);
  nand n62990(x62990, x76792, x76891);
  nand n62991(x62991, x62933, x76987);
  nand n62992(x62992, x62991, x62990);
  nand n62993(x62993, x76792, x76894);
  nand n62994(x62994, x62933, x76990);
  nand n62995(x62995, x62994, x62993);
  nand n62996(x62996, x76792, x76897);
  nand n62997(x62997, x62933, x76993);
  nand n62998(x62998, x62997, x62996);
  nand n62999(x62999, x76792, x76900);
  nand n63000(x63000, x62933, x76996);
  nand n63001(x63001, x63000, x62999);
  nand n63002(x63002, x76792, x76903);
  nand n63003(x63003, x62933, x76999);
  nand n63004(x63004, x63003, x63002);
  nand n63005(x63005, x76792, x76906);
  nand n63006(x63006, x62933, x77002);
  nand n63007(x63007, x63006, x63005);
  nand n63008(x63008, x76792, x76909);
  nand n63009(x63009, x62933, x77005);
  nand n63010(x63010, x63009, x63008);
  nand n63011(x63011, x76792, x76912);
  nand n63012(x63012, x62933, x77008);
  nand n63013(x63013, x63012, x63011);
  nand n63014(x63014, x76792, x76915);
  nand n63015(x63015, x62933, x77011);
  nand n63016(x63016, x63015, x63014);
  nand n63017(x63017, x76792, x76918);
  nand n63018(x63018, x62933, x77014);
  nand n63019(x63019, x63018, x63017);
  nand n63020(x63020, x76792, x76921);
  nand n63021(x63021, x62933, x77017);
  nand n63022(x63022, x63021, x63020);
  nand n63023(x63023, x76792, x76924);
  nand n63024(x63024, x62933, x77020);
  nand n63025(x63025, x63024, x63023);
  nand n63026(x63026, x76675, x62935);
  nand n63029(x63029, x63028, x63027);
  nand n63030(x63030, x63029, x63026);
  nand n63031(x63031, x76678, x62938);
  nand n63034(x63034, x63033, x63032);
  nand n63035(x63035, x63034, x63031);
  nand n63037(x63037, x76681, x62941);
  nand n63040(x63040, x63039, x63038);
  nand n63041(x63041, x63040, x63037);
  nand n63043(x63043, x76684, x62944);
  nand n63046(x63046, x63045, x63044);
  nand n63047(x63047, x63046, x63043);
  nand n63049(x63049, x76687, x62947);
  nand n63052(x63052, x63051, x63050);
  nand n63053(x63053, x63052, x63049);
  nand n63055(x63055, x76690, x62950);
  nand n63058(x63058, x63057, x63056);
  nand n63059(x63059, x63058, x63055);
  nand n63061(x63061, x76693, x62953);
  nand n63064(x63064, x63063, x63062);
  nand n63065(x63065, x63064, x63061);
  nand n63067(x63067, x76696, x62956);
  nand n63070(x63070, x63069, x63068);
  nand n63071(x63071, x63070, x63067);
  nand n63073(x63073, x76699, x62959);
  nand n63076(x63076, x63075, x63074);
  nand n63077(x63077, x63076, x63073);
  nand n63079(x63079, x76702, x62962);
  nand n63082(x63082, x63081, x63080);
  nand n63083(x63083, x63082, x63079);
  nand n63085(x63085, x76705, x62965);
  nand n63088(x63088, x63087, x63086);
  nand n63089(x63089, x63088, x63085);
  nand n63091(x63091, x76708, x62968);
  nand n63094(x63094, x63093, x63092);
  nand n63095(x63095, x63094, x63091);
  nand n63097(x63097, x76711, x62971);
  nand n63100(x63100, x63099, x63098);
  nand n63101(x63101, x63100, x63097);
  nand n63103(x63103, x76714, x62974);
  nand n63106(x63106, x63105, x63104);
  nand n63107(x63107, x63106, x63103);
  nand n63109(x63109, x76717, x62977);
  nand n63112(x63112, x63111, x63110);
  nand n63113(x63113, x63112, x63109);
  nand n63115(x63115, x76720, x62980);
  nand n63118(x63118, x63117, x63116);
  nand n63119(x63119, x63118, x63115);
  nand n63121(x63121, x76723, x62983);
  nand n63124(x63124, x63123, x63122);
  nand n63125(x63125, x63124, x63121);
  nand n63127(x63127, x76726, x62986);
  nand n63130(x63130, x63129, x63128);
  nand n63131(x63131, x63130, x63127);
  nand n63133(x63133, x76729, x62989);
  nand n63136(x63136, x63135, x63134);
  nand n63137(x63137, x63136, x63133);
  nand n63139(x63139, x76732, x62992);
  nand n63142(x63142, x63141, x63140);
  nand n63143(x63143, x63142, x63139);
  nand n63145(x63145, x76735, x62995);
  nand n63148(x63148, x63147, x63146);
  nand n63149(x63149, x63148, x63145);
  nand n63151(x63151, x76738, x62998);
  nand n63154(x63154, x63153, x63152);
  nand n63155(x63155, x63154, x63151);
  nand n63157(x63157, x76741, x63001);
  nand n63160(x63160, x63159, x63158);
  nand n63161(x63161, x63160, x63157);
  nand n63163(x63163, x76744, x63004);
  nand n63166(x63166, x63165, x63164);
  nand n63167(x63167, x63166, x63163);
  nand n63169(x63169, x76747, x63007);
  nand n63172(x63172, x63171, x63170);
  nand n63173(x63173, x63172, x63169);
  nand n63175(x63175, x76750, x63010);
  nand n63178(x63178, x63177, x63176);
  nand n63179(x63179, x63178, x63175);
  nand n63181(x63181, x76753, x63013);
  nand n63184(x63184, x63183, x63182);
  nand n63185(x63185, x63184, x63181);
  nand n63187(x63187, x76756, x63016);
  nand n63190(x63190, x63189, x63188);
  nand n63191(x63191, x63190, x63187);
  nand n63193(x63193, x76759, x63019);
  nand n63196(x63196, x63195, x63194);
  nand n63197(x63197, x63196, x63193);
  nand n63199(x63199, x76762, x63022);
  nand n63202(x63202, x63201, x63200);
  nand n63203(x63203, x63202, x63199);
  nand n63205(x63205, x76765, x63025);
  nand n63208(x63208, x63207, x63206);
  nand n63209(x63209, x63208, x63205);
  nand n63240(x63240, x63036, x63211);
  nand n63241(x63241, x63240, x63031);
  nand n63242(x63242, x63042, x63212);
  nand n63243(x63243, x63242, x63037);
  nand n63244(x63244, x63042, x63036);
  nand n63246(x63246, x63048, x63213);
  nand n63247(x63247, x63246, x63043);
  nand n63248(x63248, x63048, x63042);
  nand n63250(x63250, x63054, x63214);
  nand n63251(x63251, x63250, x63049);
  nand n63252(x63252, x63054, x63048);
  nand n63254(x63254, x63060, x63215);
  nand n63255(x63255, x63254, x63055);
  nand n63256(x63256, x63060, x63054);
  nand n63258(x63258, x63066, x63216);
  nand n63259(x63259, x63258, x63061);
  nand n63260(x63260, x63066, x63060);
  nand n63262(x63262, x63072, x63217);
  nand n63263(x63263, x63262, x63067);
  nand n63264(x63264, x63072, x63066);
  nand n63266(x63266, x63078, x63218);
  nand n63267(x63267, x63266, x63073);
  nand n63268(x63268, x63078, x63072);
  nand n63270(x63270, x63084, x63219);
  nand n63271(x63271, x63270, x63079);
  nand n63272(x63272, x63084, x63078);
  nand n63274(x63274, x63090, x63220);
  nand n63275(x63275, x63274, x63085);
  nand n63276(x63276, x63090, x63084);
  nand n63278(x63278, x63096, x63221);
  nand n63279(x63279, x63278, x63091);
  nand n63280(x63280, x63096, x63090);
  nand n63282(x63282, x63102, x63222);
  nand n63283(x63283, x63282, x63097);
  nand n63284(x63284, x63102, x63096);
  nand n63286(x63286, x63108, x63223);
  nand n63287(x63287, x63286, x63103);
  nand n63288(x63288, x63108, x63102);
  nand n63290(x63290, x63114, x63224);
  nand n63291(x63291, x63290, x63109);
  nand n63292(x63292, x63114, x63108);
  nand n63294(x63294, x63120, x63225);
  nand n63295(x63295, x63294, x63115);
  nand n63296(x63296, x63120, x63114);
  nand n63298(x63298, x63126, x63226);
  nand n63299(x63299, x63298, x63121);
  nand n63300(x63300, x63126, x63120);
  nand n63302(x63302, x63132, x63227);
  nand n63303(x63303, x63302, x63127);
  nand n63304(x63304, x63132, x63126);
  nand n63306(x63306, x63138, x63228);
  nand n63307(x63307, x63306, x63133);
  nand n63308(x63308, x63138, x63132);
  nand n63310(x63310, x63144, x63229);
  nand n63311(x63311, x63310, x63139);
  nand n63312(x63312, x63144, x63138);
  nand n63314(x63314, x63150, x63230);
  nand n63315(x63315, x63314, x63145);
  nand n63316(x63316, x63150, x63144);
  nand n63318(x63318, x63156, x63231);
  nand n63319(x63319, x63318, x63151);
  nand n63320(x63320, x63156, x63150);
  nand n63322(x63322, x63162, x63232);
  nand n63323(x63323, x63322, x63157);
  nand n63324(x63324, x63162, x63156);
  nand n63326(x63326, x63168, x63233);
  nand n63327(x63327, x63326, x63163);
  nand n63328(x63328, x63168, x63162);
  nand n63330(x63330, x63174, x63234);
  nand n63331(x63331, x63330, x63169);
  nand n63332(x63332, x63174, x63168);
  nand n63334(x63334, x63180, x63235);
  nand n63335(x63335, x63334, x63175);
  nand n63336(x63336, x63180, x63174);
  nand n63338(x63338, x63186, x63236);
  nand n63339(x63339, x63338, x63181);
  nand n63340(x63340, x63186, x63180);
  nand n63342(x63342, x63192, x63237);
  nand n63343(x63343, x63342, x63187);
  nand n63344(x63344, x63192, x63186);
  nand n63346(x63346, x63198, x63238);
  nand n63347(x63347, x63346, x63193);
  nand n63348(x63348, x63198, x63192);
  nand n63350(x63350, x63204, x63239);
  nand n63351(x63351, x63350, x63199);
  nand n63352(x63352, x63204, x63198);
  nand n63355(x63355, x63245, x63211);
  nand n63357(x63357, x63355, x63356);
  nand n63358(x63358, x63249, x63241);
  nand n63360(x63360, x63358, x63359);
  nand n63361(x63361, x63253, x63243);
  nand n63363(x63363, x63361, x63362);
  nand n63364(x63364, x63253, x63245);
  nand n63366(x63366, x63257, x63247);
  nand n63368(x63368, x63366, x63367);
  nand n63369(x63369, x63257, x63249);
  nand n63371(x63371, x63261, x63251);
  nand n63373(x63373, x63371, x63372);
  nand n63374(x63374, x63261, x63253);
  nand n63376(x63376, x63265, x63255);
  nand n63378(x63378, x63376, x63377);
  nand n63379(x63379, x63265, x63257);
  nand n63381(x63381, x63269, x63259);
  nand n63383(x63383, x63381, x63382);
  nand n63384(x63384, x63269, x63261);
  nand n63386(x63386, x63273, x63263);
  nand n63388(x63388, x63386, x63387);
  nand n63389(x63389, x63273, x63265);
  nand n63391(x63391, x63277, x63267);
  nand n63393(x63393, x63391, x63392);
  nand n63394(x63394, x63277, x63269);
  nand n63396(x63396, x63281, x63271);
  nand n63398(x63398, x63396, x63397);
  nand n63399(x63399, x63281, x63273);
  nand n63401(x63401, x63285, x63275);
  nand n63403(x63403, x63401, x63402);
  nand n63404(x63404, x63285, x63277);
  nand n63406(x63406, x63289, x63279);
  nand n63408(x63408, x63406, x63407);
  nand n63409(x63409, x63289, x63281);
  nand n63411(x63411, x63293, x63283);
  nand n63413(x63413, x63411, x63412);
  nand n63414(x63414, x63293, x63285);
  nand n63416(x63416, x63297, x63287);
  nand n63418(x63418, x63416, x63417);
  nand n63419(x63419, x63297, x63289);
  nand n63421(x63421, x63301, x63291);
  nand n63423(x63423, x63421, x63422);
  nand n63424(x63424, x63301, x63293);
  nand n63426(x63426, x63305, x63295);
  nand n63428(x63428, x63426, x63427);
  nand n63429(x63429, x63305, x63297);
  nand n63431(x63431, x63309, x63299);
  nand n63433(x63433, x63431, x63432);
  nand n63434(x63434, x63309, x63301);
  nand n63436(x63436, x63313, x63303);
  nand n63438(x63438, x63436, x63437);
  nand n63439(x63439, x63313, x63305);
  nand n63441(x63441, x63317, x63307);
  nand n63443(x63443, x63441, x63442);
  nand n63444(x63444, x63317, x63309);
  nand n63446(x63446, x63321, x63311);
  nand n63448(x63448, x63446, x63447);
  nand n63449(x63449, x63321, x63313);
  nand n63451(x63451, x63325, x63315);
  nand n63453(x63453, x63451, x63452);
  nand n63454(x63454, x63325, x63317);
  nand n63456(x63456, x63329, x63319);
  nand n63458(x63458, x63456, x63457);
  nand n63459(x63459, x63329, x63321);
  nand n63461(x63461, x63333, x63323);
  nand n63463(x63463, x63461, x63462);
  nand n63464(x63464, x63333, x63325);
  nand n63466(x63466, x63337, x63327);
  nand n63468(x63468, x63466, x63467);
  nand n63469(x63469, x63337, x63329);
  nand n63471(x63471, x63341, x63331);
  nand n63473(x63473, x63471, x63472);
  nand n63474(x63474, x63341, x63333);
  nand n63476(x63476, x63345, x63335);
  nand n63478(x63478, x63476, x63477);
  nand n63479(x63479, x63345, x63337);
  nand n63481(x63481, x63349, x63339);
  nand n63483(x63483, x63481, x63482);
  nand n63484(x63484, x63349, x63341);
  nand n63486(x63486, x63353, x63343);
  nand n63488(x63488, x63486, x63487);
  nand n63489(x63489, x63353, x63345);
  nand n63492(x63492, x63365, x63211);
  nand n63494(x63494, x63492, x63493);
  nand n63495(x63495, x63370, x63241);
  nand n63497(x63497, x63495, x63496);
  nand n63498(x63498, x63375, x63357);
  nand n63500(x63500, x63498, x63499);
  nand n63501(x63501, x63380, x63360);
  nand n63503(x63503, x63501, x63502);
  nand n63504(x63504, x63385, x63363);
  nand n63506(x63506, x63504, x63505);
  nand n63507(x63507, x63385, x63365);
  nand n63509(x63509, x63390, x63368);
  nand n63511(x63511, x63509, x63510);
  nand n63512(x63512, x63390, x63370);
  nand n63514(x63514, x63395, x63373);
  nand n63516(x63516, x63514, x63515);
  nand n63517(x63517, x63395, x63375);
  nand n63519(x63519, x63400, x63378);
  nand n63521(x63521, x63519, x63520);
  nand n63522(x63522, x63400, x63380);
  nand n63524(x63524, x63405, x63383);
  nand n63526(x63526, x63524, x63525);
  nand n63527(x63527, x63405, x63385);
  nand n63529(x63529, x63410, x63388);
  nand n63531(x63531, x63529, x63530);
  nand n63532(x63532, x63410, x63390);
  nand n63534(x63534, x63415, x63393);
  nand n63536(x63536, x63534, x63535);
  nand n63537(x63537, x63415, x63395);
  nand n63539(x63539, x63420, x63398);
  nand n63541(x63541, x63539, x63540);
  nand n63542(x63542, x63420, x63400);
  nand n63544(x63544, x63425, x63403);
  nand n63546(x63546, x63544, x63545);
  nand n63547(x63547, x63425, x63405);
  nand n63549(x63549, x63430, x63408);
  nand n63551(x63551, x63549, x63550);
  nand n63552(x63552, x63430, x63410);
  nand n63554(x63554, x63435, x63413);
  nand n63556(x63556, x63554, x63555);
  nand n63557(x63557, x63435, x63415);
  nand n63559(x63559, x63440, x63418);
  nand n63561(x63561, x63559, x63560);
  nand n63562(x63562, x63440, x63420);
  nand n63564(x63564, x63445, x63423);
  nand n63566(x63566, x63564, x63565);
  nand n63567(x63567, x63445, x63425);
  nand n63569(x63569, x63450, x63428);
  nand n63571(x63571, x63569, x63570);
  nand n63572(x63572, x63450, x63430);
  nand n63574(x63574, x63455, x63433);
  nand n63576(x63576, x63574, x63575);
  nand n63577(x63577, x63455, x63435);
  nand n63579(x63579, x63460, x63438);
  nand n63581(x63581, x63579, x63580);
  nand n63582(x63582, x63460, x63440);
  nand n63584(x63584, x63465, x63443);
  nand n63586(x63586, x63584, x63585);
  nand n63587(x63587, x63465, x63445);
  nand n63589(x63589, x63470, x63448);
  nand n63591(x63591, x63589, x63590);
  nand n63592(x63592, x63470, x63450);
  nand n63594(x63594, x63475, x63453);
  nand n63596(x63596, x63594, x63595);
  nand n63597(x63597, x63475, x63455);
  nand n63599(x63599, x63480, x63458);
  nand n63601(x63601, x63599, x63600);
  nand n63602(x63602, x63480, x63460);
  nand n63604(x63604, x63485, x63463);
  nand n63606(x63606, x63604, x63605);
  nand n63607(x63607, x63485, x63465);
  nand n63609(x63609, x63490, x63468);
  nand n63611(x63611, x63609, x63610);
  nand n63612(x63612, x63490, x63470);
  nand n63615(x63615, x63508, x63211);
  nand n63617(x63617, x63615, x63616);
  nand n63618(x63618, x63513, x63241);
  nand n63620(x63620, x63618, x63619);
  nand n63621(x63621, x63518, x63357);
  nand n63623(x63623, x63621, x63622);
  nand n63624(x63624, x63523, x63360);
  nand n63626(x63626, x63624, x63625);
  nand n63627(x63627, x63528, x63494);
  nand n63629(x63629, x63627, x63628);
  nand n63630(x63630, x63533, x63497);
  nand n63632(x63632, x63630, x63631);
  nand n63633(x63633, x63538, x63500);
  nand n63635(x63635, x63633, x63634);
  nand n63636(x63636, x63543, x63503);
  nand n63638(x63638, x63636, x63637);
  nand n63639(x63639, x63548, x63506);
  nand n63641(x63641, x63639, x63640);
  nand n63642(x63642, x63548, x63508);
  nand n63644(x63644, x63553, x63511);
  nand n63646(x63646, x63644, x63645);
  nand n63647(x63647, x63553, x63513);
  nand n63649(x63649, x63558, x63516);
  nand n63651(x63651, x63649, x63650);
  nand n63652(x63652, x63558, x63518);
  nand n63654(x63654, x63563, x63521);
  nand n63656(x63656, x63654, x63655);
  nand n63657(x63657, x63563, x63523);
  nand n63659(x63659, x63568, x63526);
  nand n63661(x63661, x63659, x63660);
  nand n63662(x63662, x63568, x63528);
  nand n63664(x63664, x63573, x63531);
  nand n63666(x63666, x63664, x63665);
  nand n63667(x63667, x63573, x63533);
  nand n63669(x63669, x63578, x63536);
  nand n63671(x63671, x63669, x63670);
  nand n63672(x63672, x63578, x63538);
  nand n63674(x63674, x63583, x63541);
  nand n63676(x63676, x63674, x63675);
  nand n63677(x63677, x63583, x63543);
  nand n63679(x63679, x63588, x63546);
  nand n63681(x63681, x63679, x63680);
  nand n63682(x63682, x63588, x63548);
  nand n63684(x63684, x63593, x63551);
  nand n63686(x63686, x63684, x63685);
  nand n63687(x63687, x63593, x63553);
  nand n63689(x63689, x63598, x63556);
  nand n63691(x63691, x63689, x63690);
  nand n63692(x63692, x63598, x63558);
  nand n63694(x63694, x63603, x63561);
  nand n63696(x63696, x63694, x63695);
  nand n63697(x63697, x63603, x63563);
  nand n63699(x63699, x63608, x63566);
  nand n63701(x63701, x63699, x63700);
  nand n63702(x63702, x63608, x63568);
  nand n63704(x63704, x63613, x63571);
  nand n63706(x63706, x63704, x63705);
  nand n63707(x63707, x63613, x63573);
  nand n63710(x63710, x63643, x63211);
  nand n63712(x63712, x63710, x63711);
  nand n63713(x63713, x63648, x63241);
  nand n63715(x63715, x63713, x63714);
  nand n63716(x63716, x63653, x63357);
  nand n63718(x63718, x63716, x63717);
  nand n63719(x63719, x63658, x63360);
  nand n63721(x63721, x63719, x63720);
  nand n63722(x63722, x63663, x63494);
  nand n63724(x63724, x63722, x63723);
  nand n63725(x63725, x63668, x63497);
  nand n63727(x63727, x63725, x63726);
  nand n63728(x63728, x63673, x63500);
  nand n63730(x63730, x63728, x63729);
  nand n63731(x63731, x63678, x63503);
  nand n63733(x63733, x63731, x63732);
  nand n63734(x63734, x63683, x63617);
  nand n63736(x63736, x63734, x63735);
  nand n63737(x63737, x63688, x63620);
  nand n63739(x63739, x63737, x63738);
  nand n63740(x63740, x63693, x63623);
  nand n63742(x63742, x63740, x63741);
  nand n63743(x63743, x63698, x63626);
  nand n63745(x63745, x63743, x63744);
  nand n63746(x63746, x63703, x63629);
  nand n63748(x63748, x63746, x63747);
  nand n63749(x63749, x63708, x63632);
  nand n63751(x63751, x63749, x63750);
  nand n63752(x63752, x63035, x63026);
  nand n63753(x63753, x63752, x63240);
  nand n63754(x63754, x63042, x63241);
  nand n63755(x63755, x63041, x63354);
  nand n63756(x63756, x63755, x63754);
  nand n63758(x63758, x63048, x63357);
  nand n63760(x63760, x63047, x63759);
  nand n63761(x63761, x63760, x63758);
  nand n63763(x63763, x63054, x63360);
  nand n63764(x63764, x63053, x63491);
  nand n63765(x63765, x63764, x63763);
  nand n63767(x63767, x63060, x63494);
  nand n63769(x63769, x63059, x63768);
  nand n63770(x63770, x63769, x63767);
  nand n63772(x63772, x63066, x63497);
  nand n63774(x63774, x63065, x63773);
  nand n63775(x63775, x63774, x63772);
  nand n63777(x63777, x63072, x63500);
  nand n63779(x63779, x63071, x63778);
  nand n63780(x63780, x63779, x63777);
  nand n63782(x63782, x63078, x63503);
  nand n63783(x63783, x63077, x63614);
  nand n63784(x63784, x63783, x63782);
  nand n63786(x63786, x63084, x63617);
  nand n63788(x63788, x63083, x63787);
  nand n63789(x63789, x63788, x63786);
  nand n63791(x63791, x63090, x63620);
  nand n63793(x63793, x63089, x63792);
  nand n63794(x63794, x63793, x63791);
  nand n63795(x63795, x63096, x63623);
  nand n63797(x63797, x63095, x63796);
  nand n63798(x63798, x63797, x63795);
  nand n63799(x63799, x63102, x63626);
  nand n63801(x63801, x63101, x63800);
  nand n63802(x63802, x63801, x63799);
  nand n63803(x63803, x63108, x63629);
  nand n63805(x63805, x63107, x63804);
  nand n63806(x63806, x63805, x63803);
  nand n63807(x63807, x63114, x63632);
  nand n63809(x63809, x63113, x63808);
  nand n63810(x63810, x63809, x63807);
  nand n63811(x63811, x63120, x63635);
  nand n63813(x63813, x63119, x63812);
  nand n63814(x63814, x63813, x63811);
  nand n63815(x63815, x63126, x63638);
  nand n63816(x63816, x63125, x63709);
  nand n63817(x63817, x63816, x63815);
  nand n63818(x63818, x63132, x63712);
  nand n63820(x63820, x63131, x63819);
  nand n63821(x63821, x63820, x63818);
  nand n63822(x63822, x63138, x63715);
  nand n63824(x63824, x63137, x63823);
  nand n63825(x63825, x63824, x63822);
  nand n63826(x63826, x63144, x63718);
  nand n63828(x63828, x63143, x63827);
  nand n63829(x63829, x63828, x63826);
  nand n63830(x63830, x63150, x63721);
  nand n63832(x63832, x63149, x63831);
  nand n63833(x63833, x63832, x63830);
  nand n63834(x63834, x63156, x63724);
  nand n63836(x63836, x63155, x63835);
  nand n63837(x63837, x63836, x63834);
  nand n63838(x63838, x63162, x63727);
  nand n63840(x63840, x63161, x63839);
  nand n63841(x63841, x63840, x63838);
  nand n63842(x63842, x63168, x63730);
  nand n63844(x63844, x63167, x63843);
  nand n63845(x63845, x63844, x63842);
  nand n63846(x63846, x63174, x63733);
  nand n63848(x63848, x63173, x63847);
  nand n63849(x63849, x63848, x63846);
  nand n63850(x63850, x63180, x63736);
  nand n63852(x63852, x63179, x63851);
  nand n63853(x63853, x63852, x63850);
  nand n63854(x63854, x63186, x63739);
  nand n63856(x63856, x63185, x63855);
  nand n63857(x63857, x63856, x63854);
  nand n63858(x63858, x63192, x63742);
  nand n63860(x63860, x63191, x63859);
  nand n63861(x63861, x63860, x63858);
  nand n63862(x63862, x63198, x63745);
  nand n63864(x63864, x63197, x63863);
  nand n63865(x63865, x63864, x63862);
  nand n63866(x63866, x63204, x63748);
  nand n63868(x63868, x63203, x63867);
  nand n63869(x63869, x63868, x63866);
  nand n63870(x63870, x63210, x63751);
  nand n63872(x63872, x63209, x63871);
  nand n63873(x63873, x63872, x63870);
  nand n63874(x63874, x83367, x62933);
  nand n63913(x63913, x63908, x63877);
  nand n63915(x63915, x63914, x63876);
  nand n63916(x63916, x63915, x63913);
  nand n63917(x63917, x63908, x63878);
  nand n63918(x63918, x63914, x63877);
  nand n63919(x63919, x63918, x63917);
  nand n63920(x63920, x63908, x63879);
  nand n63921(x63921, x63914, x63878);
  nand n63922(x63922, x63921, x63920);
  nand n63923(x63923, x63908, x63880);
  nand n63924(x63924, x63914, x63879);
  nand n63925(x63925, x63924, x63923);
  nand n63926(x63926, x63908, x63881);
  nand n63927(x63927, x63914, x63880);
  nand n63928(x63928, x63927, x63926);
  nand n63929(x63929, x63908, x63882);
  nand n63930(x63930, x63914, x63881);
  nand n63931(x63931, x63930, x63929);
  nand n63932(x63932, x63908, x63883);
  nand n63933(x63933, x63914, x63882);
  nand n63934(x63934, x63933, x63932);
  nand n63935(x63935, x63908, x63884);
  nand n63936(x63936, x63914, x63883);
  nand n63937(x63937, x63936, x63935);
  nand n63938(x63938, x63908, x63885);
  nand n63939(x63939, x63914, x63884);
  nand n63940(x63940, x63939, x63938);
  nand n63941(x63941, x63908, x63886);
  nand n63942(x63942, x63914, x63885);
  nand n63943(x63943, x63942, x63941);
  nand n63944(x63944, x63908, x63887);
  nand n63945(x63945, x63914, x63886);
  nand n63946(x63946, x63945, x63944);
  nand n63947(x63947, x63908, x63888);
  nand n63948(x63948, x63914, x63887);
  nand n63949(x63949, x63948, x63947);
  nand n63950(x63950, x63908, x63889);
  nand n63951(x63951, x63914, x63888);
  nand n63952(x63952, x63951, x63950);
  nand n63953(x63953, x63908, x63890);
  nand n63954(x63954, x63914, x63889);
  nand n63955(x63955, x63954, x63953);
  nand n63956(x63956, x63908, x63891);
  nand n63957(x63957, x63914, x63890);
  nand n63958(x63958, x63957, x63956);
  nand n63959(x63959, x63908, x63892);
  nand n63960(x63960, x63914, x63891);
  nand n63961(x63961, x63960, x63959);
  nand n63962(x63962, x63908, x63893);
  nand n63963(x63963, x63914, x63892);
  nand n63964(x63964, x63963, x63962);
  nand n63965(x63965, x63908, x63894);
  nand n63966(x63966, x63914, x63893);
  nand n63967(x63967, x63966, x63965);
  nand n63968(x63968, x63908, x63895);
  nand n63969(x63969, x63914, x63894);
  nand n63970(x63970, x63969, x63968);
  nand n63971(x63971, x63908, x63896);
  nand n63972(x63972, x63914, x63895);
  nand n63973(x63973, x63972, x63971);
  nand n63974(x63974, x63908, x63897);
  nand n63975(x63975, x63914, x63896);
  nand n63976(x63976, x63975, x63974);
  nand n63977(x63977, x63908, x63898);
  nand n63978(x63978, x63914, x63897);
  nand n63979(x63979, x63978, x63977);
  nand n63980(x63980, x63908, x63899);
  nand n63981(x63981, x63914, x63898);
  nand n63982(x63982, x63981, x63980);
  nand n63983(x63983, x63908, x63900);
  nand n63984(x63984, x63914, x63899);
  nand n63985(x63985, x63984, x63983);
  nand n63986(x63986, x63908, x63901);
  nand n63987(x63987, x63914, x63900);
  nand n63988(x63988, x63987, x63986);
  nand n63989(x63989, x63908, x63902);
  nand n63990(x63990, x63914, x63901);
  nand n63991(x63991, x63990, x63989);
  nand n63992(x63992, x63908, x63903);
  nand n63993(x63993, x63914, x63902);
  nand n63994(x63994, x63993, x63992);
  nand n63995(x63995, x63908, x63904);
  nand n63996(x63996, x63914, x63903);
  nand n63997(x63997, x63996, x63995);
  nand n63998(x63998, x63908, x63905);
  nand n63999(x63999, x63914, x63904);
  nand n64000(x64000, x63999, x63998);
  nand n64001(x64001, x63908, x63906);
  nand n64002(x64002, x63914, x63905);
  nand n64003(x64003, x64002, x64001);
  nand n64004(x64004, x63908, x63907);
  nand n64005(x64005, x63914, x63906);
  nand n64006(x64006, x64005, x64004);
  nand n64007(x64007, x63914, x63907);
  nand n64008(x64008, x63909, x63922);
  nand n64010(x64010, x64009, x63916);
  nand n64011(x64011, x64010, x64008);
  nand n64012(x64012, x63909, x63925);
  nand n64013(x64013, x64009, x63919);
  nand n64014(x64014, x64013, x64012);
  nand n64015(x64015, x63909, x63928);
  nand n64016(x64016, x64009, x63922);
  nand n64017(x64017, x64016, x64015);
  nand n64018(x64018, x63909, x63931);
  nand n64019(x64019, x64009, x63925);
  nand n64020(x64020, x64019, x64018);
  nand n64021(x64021, x63909, x63934);
  nand n64022(x64022, x64009, x63928);
  nand n64023(x64023, x64022, x64021);
  nand n64024(x64024, x63909, x63937);
  nand n64025(x64025, x64009, x63931);
  nand n64026(x64026, x64025, x64024);
  nand n64027(x64027, x63909, x63940);
  nand n64028(x64028, x64009, x63934);
  nand n64029(x64029, x64028, x64027);
  nand n64030(x64030, x63909, x63943);
  nand n64031(x64031, x64009, x63937);
  nand n64032(x64032, x64031, x64030);
  nand n64033(x64033, x63909, x63946);
  nand n64034(x64034, x64009, x63940);
  nand n64035(x64035, x64034, x64033);
  nand n64036(x64036, x63909, x63949);
  nand n64037(x64037, x64009, x63943);
  nand n64038(x64038, x64037, x64036);
  nand n64039(x64039, x63909, x63952);
  nand n64040(x64040, x64009, x63946);
  nand n64041(x64041, x64040, x64039);
  nand n64042(x64042, x63909, x63955);
  nand n64043(x64043, x64009, x63949);
  nand n64044(x64044, x64043, x64042);
  nand n64045(x64045, x63909, x63958);
  nand n64046(x64046, x64009, x63952);
  nand n64047(x64047, x64046, x64045);
  nand n64048(x64048, x63909, x63961);
  nand n64049(x64049, x64009, x63955);
  nand n64050(x64050, x64049, x64048);
  nand n64051(x64051, x63909, x63964);
  nand n64052(x64052, x64009, x63958);
  nand n64053(x64053, x64052, x64051);
  nand n64054(x64054, x63909, x63967);
  nand n64055(x64055, x64009, x63961);
  nand n64056(x64056, x64055, x64054);
  nand n64057(x64057, x63909, x63970);
  nand n64058(x64058, x64009, x63964);
  nand n64059(x64059, x64058, x64057);
  nand n64060(x64060, x63909, x63973);
  nand n64061(x64061, x64009, x63967);
  nand n64062(x64062, x64061, x64060);
  nand n64063(x64063, x63909, x63976);
  nand n64064(x64064, x64009, x63970);
  nand n64065(x64065, x64064, x64063);
  nand n64066(x64066, x63909, x63979);
  nand n64067(x64067, x64009, x63973);
  nand n64068(x64068, x64067, x64066);
  nand n64069(x64069, x63909, x63982);
  nand n64070(x64070, x64009, x63976);
  nand n64071(x64071, x64070, x64069);
  nand n64072(x64072, x63909, x63985);
  nand n64073(x64073, x64009, x63979);
  nand n64074(x64074, x64073, x64072);
  nand n64075(x64075, x63909, x63988);
  nand n64076(x64076, x64009, x63982);
  nand n64077(x64077, x64076, x64075);
  nand n64078(x64078, x63909, x63991);
  nand n64079(x64079, x64009, x63985);
  nand n64080(x64080, x64079, x64078);
  nand n64081(x64081, x63909, x63994);
  nand n64082(x64082, x64009, x63988);
  nand n64083(x64083, x64082, x64081);
  nand n64084(x64084, x63909, x63997);
  nand n64085(x64085, x64009, x63991);
  nand n64086(x64086, x64085, x64084);
  nand n64087(x64087, x63909, x64000);
  nand n64088(x64088, x64009, x63994);
  nand n64089(x64089, x64088, x64087);
  nand n64090(x64090, x63909, x64003);
  nand n64091(x64091, x64009, x63997);
  nand n64092(x64092, x64091, x64090);
  nand n64093(x64093, x63909, x64006);
  nand n64094(x64094, x64009, x64000);
  nand n64095(x64095, x64094, x64093);
  nand n64096(x64096, x63909, x86266);
  nand n64097(x64097, x64009, x64003);
  nand n64098(x64098, x64097, x64096);
  nand n64099(x64099, x64009, x64006);
  nand n64100(x64100, x64009, x86266);
  nand n64101(x64101, x63910, x64023);
  nand n64103(x64103, x64102, x64011);
  nand n64104(x64104, x64103, x64101);
  nand n64105(x64105, x63910, x64026);
  nand n64106(x64106, x64102, x64014);
  nand n64107(x64107, x64106, x64105);
  nand n64108(x64108, x63910, x64029);
  nand n64109(x64109, x64102, x64017);
  nand n64110(x64110, x64109, x64108);
  nand n64111(x64111, x63910, x64032);
  nand n64112(x64112, x64102, x64020);
  nand n64113(x64113, x64112, x64111);
  nand n64114(x64114, x63910, x64035);
  nand n64115(x64115, x64102, x64023);
  nand n64116(x64116, x64115, x64114);
  nand n64117(x64117, x63910, x64038);
  nand n64118(x64118, x64102, x64026);
  nand n64119(x64119, x64118, x64117);
  nand n64120(x64120, x63910, x64041);
  nand n64121(x64121, x64102, x64029);
  nand n64122(x64122, x64121, x64120);
  nand n64123(x64123, x63910, x64044);
  nand n64124(x64124, x64102, x64032);
  nand n64125(x64125, x64124, x64123);
  nand n64126(x64126, x63910, x64047);
  nand n64127(x64127, x64102, x64035);
  nand n64128(x64128, x64127, x64126);
  nand n64129(x64129, x63910, x64050);
  nand n64130(x64130, x64102, x64038);
  nand n64131(x64131, x64130, x64129);
  nand n64132(x64132, x63910, x64053);
  nand n64133(x64133, x64102, x64041);
  nand n64134(x64134, x64133, x64132);
  nand n64135(x64135, x63910, x64056);
  nand n64136(x64136, x64102, x64044);
  nand n64137(x64137, x64136, x64135);
  nand n64138(x64138, x63910, x64059);
  nand n64139(x64139, x64102, x64047);
  nand n64140(x64140, x64139, x64138);
  nand n64141(x64141, x63910, x64062);
  nand n64142(x64142, x64102, x64050);
  nand n64143(x64143, x64142, x64141);
  nand n64144(x64144, x63910, x64065);
  nand n64145(x64145, x64102, x64053);
  nand n64146(x64146, x64145, x64144);
  nand n64147(x64147, x63910, x64068);
  nand n64148(x64148, x64102, x64056);
  nand n64149(x64149, x64148, x64147);
  nand n64150(x64150, x63910, x64071);
  nand n64151(x64151, x64102, x64059);
  nand n64152(x64152, x64151, x64150);
  nand n64153(x64153, x63910, x64074);
  nand n64154(x64154, x64102, x64062);
  nand n64155(x64155, x64154, x64153);
  nand n64156(x64156, x63910, x64077);
  nand n64157(x64157, x64102, x64065);
  nand n64158(x64158, x64157, x64156);
  nand n64159(x64159, x63910, x64080);
  nand n64160(x64160, x64102, x64068);
  nand n64161(x64161, x64160, x64159);
  nand n64162(x64162, x63910, x64083);
  nand n64163(x64163, x64102, x64071);
  nand n64164(x64164, x64163, x64162);
  nand n64165(x64165, x63910, x64086);
  nand n64166(x64166, x64102, x64074);
  nand n64167(x64167, x64166, x64165);
  nand n64168(x64168, x63910, x64089);
  nand n64169(x64169, x64102, x64077);
  nand n64170(x64170, x64169, x64168);
  nand n64171(x64171, x63910, x64092);
  nand n64172(x64172, x64102, x64080);
  nand n64173(x64173, x64172, x64171);
  nand n64174(x64174, x63910, x64095);
  nand n64175(x64175, x64102, x64083);
  nand n64176(x64176, x64175, x64174);
  nand n64177(x64177, x63910, x64098);
  nand n64178(x64178, x64102, x64086);
  nand n64179(x64179, x64178, x64177);
  nand n64180(x64180, x63910, x86267);
  nand n64181(x64181, x64102, x64089);
  nand n64182(x64182, x64181, x64180);
  nand n64183(x64183, x63910, x86268);
  nand n64184(x64184, x64102, x64092);
  nand n64185(x64185, x64184, x64183);
  nand n64186(x64186, x64102, x64095);
  nand n64187(x64187, x64102, x64098);
  nand n64188(x64188, x64102, x86267);
  nand n64189(x64189, x64102, x86268);
  nand n64190(x64190, x63911, x64128);
  nand n64192(x64192, x64191, x64104);
  nand n64193(x64193, x64192, x64190);
  nand n64194(x64194, x63911, x64131);
  nand n64195(x64195, x64191, x64107);
  nand n64196(x64196, x64195, x64194);
  nand n64197(x64197, x63911, x64134);
  nand n64198(x64198, x64191, x64110);
  nand n64199(x64199, x64198, x64197);
  nand n64200(x64200, x63911, x64137);
  nand n64201(x64201, x64191, x64113);
  nand n64202(x64202, x64201, x64200);
  nand n64203(x64203, x63911, x64140);
  nand n64204(x64204, x64191, x64116);
  nand n64205(x64205, x64204, x64203);
  nand n64206(x64206, x63911, x64143);
  nand n64207(x64207, x64191, x64119);
  nand n64208(x64208, x64207, x64206);
  nand n64209(x64209, x63911, x64146);
  nand n64210(x64210, x64191, x64122);
  nand n64211(x64211, x64210, x64209);
  nand n64212(x64212, x63911, x64149);
  nand n64213(x64213, x64191, x64125);
  nand n64214(x64214, x64213, x64212);
  nand n64215(x64215, x63911, x64152);
  nand n64216(x64216, x64191, x64128);
  nand n64217(x64217, x64216, x64215);
  nand n64218(x64218, x63911, x64155);
  nand n64219(x64219, x64191, x64131);
  nand n64220(x64220, x64219, x64218);
  nand n64221(x64221, x63911, x64158);
  nand n64222(x64222, x64191, x64134);
  nand n64223(x64223, x64222, x64221);
  nand n64224(x64224, x63911, x64161);
  nand n64225(x64225, x64191, x64137);
  nand n64226(x64226, x64225, x64224);
  nand n64227(x64227, x63911, x64164);
  nand n64228(x64228, x64191, x64140);
  nand n64229(x64229, x64228, x64227);
  nand n64230(x64230, x63911, x64167);
  nand n64231(x64231, x64191, x64143);
  nand n64232(x64232, x64231, x64230);
  nand n64233(x64233, x63911, x64170);
  nand n64234(x64234, x64191, x64146);
  nand n64235(x64235, x64234, x64233);
  nand n64236(x64236, x63911, x64173);
  nand n64237(x64237, x64191, x64149);
  nand n64238(x64238, x64237, x64236);
  nand n64239(x64239, x63911, x64176);
  nand n64240(x64240, x64191, x64152);
  nand n64241(x64241, x64240, x64239);
  nand n64242(x64242, x63911, x64179);
  nand n64243(x64243, x64191, x64155);
  nand n64244(x64244, x64243, x64242);
  nand n64245(x64245, x63911, x64182);
  nand n64246(x64246, x64191, x64158);
  nand n64247(x64247, x64246, x64245);
  nand n64248(x64248, x63911, x64185);
  nand n64249(x64249, x64191, x64161);
  nand n64250(x64250, x64249, x64248);
  nand n64251(x64251, x63911, x86269);
  nand n64252(x64252, x64191, x64164);
  nand n64253(x64253, x64252, x64251);
  nand n64254(x64254, x63911, x86270);
  nand n64255(x64255, x64191, x64167);
  nand n64256(x64256, x64255, x64254);
  nand n64257(x64257, x63911, x86271);
  nand n64258(x64258, x64191, x64170);
  nand n64259(x64259, x64258, x64257);
  nand n64260(x64260, x63911, x86272);
  nand n64261(x64261, x64191, x64173);
  nand n64262(x64262, x64261, x64260);
  nand n64263(x64263, x64191, x64176);
  nand n64264(x64264, x64191, x64179);
  nand n64265(x64265, x64191, x64182);
  nand n64266(x64266, x64191, x64185);
  nand n64267(x64267, x64191, x86269);
  nand n64268(x64268, x64191, x86270);
  nand n64269(x64269, x64191, x86271);
  nand n64270(x64270, x64191, x86272);
  nand n64271(x64271, x63912, x64241);
  nand n64273(x64273, x64272, x64193);
  nand n64274(x64274, x64273, x64271);
  nand n64275(x64275, x63912, x64244);
  nand n64276(x64276, x64272, x64196);
  nand n64277(x64277, x64276, x64275);
  nand n64278(x64278, x63912, x64247);
  nand n64279(x64279, x64272, x64199);
  nand n64280(x64280, x64279, x64278);
  nand n64281(x64281, x63912, x64250);
  nand n64282(x64282, x64272, x64202);
  nand n64283(x64283, x64282, x64281);
  nand n64284(x64284, x63912, x64253);
  nand n64285(x64285, x64272, x64205);
  nand n64286(x64286, x64285, x64284);
  nand n64287(x64287, x63912, x64256);
  nand n64288(x64288, x64272, x64208);
  nand n64289(x64289, x64288, x64287);
  nand n64290(x64290, x63912, x64259);
  nand n64291(x64291, x64272, x64211);
  nand n64292(x64292, x64291, x64290);
  nand n64293(x64293, x63912, x64262);
  nand n64294(x64294, x64272, x64214);
  nand n64295(x64295, x64294, x64293);
  nand n64296(x64296, x63912, x86273);
  nand n64297(x64297, x64272, x64217);
  nand n64298(x64298, x64297, x64296);
  nand n64299(x64299, x63912, x86274);
  nand n64300(x64300, x64272, x64220);
  nand n64301(x64301, x64300, x64299);
  nand n64302(x64302, x63912, x86275);
  nand n64303(x64303, x64272, x64223);
  nand n64304(x64304, x64303, x64302);
  nand n64305(x64305, x63912, x86276);
  nand n64306(x64306, x64272, x64226);
  nand n64307(x64307, x64306, x64305);
  nand n64308(x64308, x63912, x86277);
  nand n64309(x64309, x64272, x64229);
  nand n64310(x64310, x64309, x64308);
  nand n64311(x64311, x63912, x86278);
  nand n64312(x64312, x64272, x64232);
  nand n64313(x64313, x64312, x64311);
  nand n64314(x64314, x63912, x86279);
  nand n64315(x64315, x64272, x64235);
  nand n64316(x64316, x64315, x64314);
  nand n64317(x64317, x63912, x86280);
  nand n64318(x64318, x64272, x64238);
  nand n64319(x64319, x64318, x64317);
  nand n64320(x64320, x64272, x64241);
  nand n64321(x64321, x64272, x64244);
  nand n64322(x64322, x64272, x64247);
  nand n64323(x64323, x64272, x64250);
  nand n64324(x64324, x64272, x64253);
  nand n64325(x64325, x64272, x64256);
  nand n64326(x64326, x64272, x64259);
  nand n64327(x64327, x64272, x64262);
  nand n64328(x64328, x64272, x86273);
  nand n64329(x64329, x64272, x86274);
  nand n64330(x64330, x64272, x86275);
  nand n64331(x64331, x64272, x86276);
  nand n64332(x64332, x64272, x86277);
  nand n64333(x64333, x64272, x86278);
  nand n64334(x64334, x64272, x86279);
  nand n64335(x64335, x64272, x86280);
  nand n64336(x64336, x63869, x63873);
  nand n64338(x64338, x63861, x63865);
  nand n64340(x64340, x63853, x63857);
  nand n64342(x64342, x63845, x63849);
  nand n64344(x64344, x63837, x63841);
  nand n64346(x64346, x63829, x63833);
  nand n64348(x64348, x63821, x63825);
  nand n64350(x64350, x63814, x63817);
  nand n64352(x64352, x63806, x63810);
  nand n64354(x64354, x63798, x63802);
  nand n64356(x64356, x63789, x63794);
  nand n64358(x64358, x63780, x63784);
  nand n64360(x64360, x63770, x63775);
  nand n64362(x64362, x63761, x63765);
  nand n64364(x64364, x63753, x63756);
  nand n64366(x64366, x64337, x63030);
  nand n64368(x64368, x64341, x64339);
  nand n64370(x64370, x64345, x64343);
  nand n64372(x64372, x64349, x64347);
  nand n64374(x64374, x64353, x64351);
  nand n64376(x64376, x64357, x64355);
  nand n64378(x64378, x64361, x64359);
  nand n64380(x64380, x64365, x64363);
  nand n64382(x64382, x64369, x64367);
  nand n64384(x64384, x64373, x64371);
  nand n64386(x64386, x64377, x64375);
  nand n64388(x64388, x64381, x64379);
  nand n64390(x64390, x64385, x64383);
  nand n64392(x64392, x64389, x64387);
  nand n64394(x64394, x64393, x64391);
  nand n64396(x64396, x63875, x64395);
  nand n64398(x64398, x76792, x77128);
  nand n64399(x64399, x62933, x77224);
  nand n64400(x64400, x64399, x64398);
  nand n64401(x64401, x76792, x77131);
  nand n64402(x64402, x62933, x77227);
  nand n64403(x64403, x64402, x64401);
  nand n64404(x64404, x76792, x77134);
  nand n64405(x64405, x62933, x77230);
  nand n64406(x64406, x64405, x64404);
  nand n64407(x64407, x76792, x77137);
  nand n64408(x64408, x62933, x77233);
  nand n64409(x64409, x64408, x64407);
  nand n64410(x64410, x76792, x77140);
  nand n64411(x64411, x62933, x77236);
  nand n64412(x64412, x64411, x64410);
  nand n64413(x64413, x76792, x77143);
  nand n64414(x64414, x62933, x77239);
  nand n64415(x64415, x64414, x64413);
  nand n64416(x64416, x76792, x77146);
  nand n64417(x64417, x62933, x77242);
  nand n64418(x64418, x64417, x64416);
  nand n64419(x64419, x76792, x77149);
  nand n64420(x64420, x62933, x77245);
  nand n64421(x64421, x64420, x64419);
  nand n64422(x64422, x76792, x77152);
  nand n64423(x64423, x62933, x77248);
  nand n64424(x64424, x64423, x64422);
  nand n64425(x64425, x76792, x77155);
  nand n64426(x64426, x62933, x77251);
  nand n64427(x64427, x64426, x64425);
  nand n64428(x64428, x76675, x64400);
  nand n64430(x64430, x63028, x64429);
  nand n64431(x64431, x64430, x64428);
  nand n64432(x64432, x76678, x64403);
  nand n64434(x64434, x63033, x64433);
  nand n64435(x64435, x64434, x64432);
  nand n64437(x64437, x76681, x64406);
  nand n64439(x64439, x63039, x64438);
  nand n64440(x64440, x64439, x64437);
  nand n64442(x64442, x76684, x64409);
  nand n64444(x64444, x63045, x64443);
  nand n64445(x64445, x64444, x64442);
  nand n64447(x64447, x76687, x64412);
  nand n64449(x64449, x63051, x64448);
  nand n64450(x64450, x64449, x64447);
  nand n64452(x64452, x76690, x64415);
  nand n64454(x64454, x63057, x64453);
  nand n64455(x64455, x64454, x64452);
  nand n64457(x64457, x76693, x64418);
  nand n64459(x64459, x63063, x64458);
  nand n64460(x64460, x64459, x64457);
  nand n64462(x64462, x76696, x64421);
  nand n64464(x64464, x63069, x64463);
  nand n64465(x64465, x64464, x64462);
  nand n64467(x64467, x76699, x64424);
  nand n64469(x64469, x63075, x64468);
  nand n64470(x64470, x64469, x64467);
  nand n64472(x64472, x76702, x64427);
  nand n64474(x64474, x63081, x64473);
  nand n64475(x64475, x64474, x64472);
  nand n64485(x64485, x64436, x64477);
  nand n64486(x64486, x64485, x64432);
  nand n64487(x64487, x64441, x64478);
  nand n64488(x64488, x64487, x64437);
  nand n64489(x64489, x64441, x64436);
  nand n64491(x64491, x64446, x64479);
  nand n64492(x64492, x64491, x64442);
  nand n64493(x64493, x64446, x64441);
  nand n64495(x64495, x64451, x64480);
  nand n64496(x64496, x64495, x64447);
  nand n64497(x64497, x64451, x64446);
  nand n64499(x64499, x64456, x64481);
  nand n64500(x64500, x64499, x64452);
  nand n64501(x64501, x64456, x64451);
  nand n64503(x64503, x64461, x64482);
  nand n64504(x64504, x64503, x64457);
  nand n64505(x64505, x64461, x64456);
  nand n64507(x64507, x64466, x64483);
  nand n64508(x64508, x64507, x64462);
  nand n64509(x64509, x64466, x64461);
  nand n64511(x64511, x64471, x64484);
  nand n64512(x64512, x64511, x64467);
  nand n64513(x64513, x64471, x64466);
  nand n64516(x64516, x64490, x64477);
  nand n64518(x64518, x64516, x64517);
  nand n64519(x64519, x64494, x64486);
  nand n64521(x64521, x64519, x64520);
  nand n64522(x64522, x64498, x64488);
  nand n64524(x64524, x64522, x64523);
  nand n64525(x64525, x64498, x64490);
  nand n64527(x64527, x64502, x64492);
  nand n64529(x64529, x64527, x64528);
  nand n64530(x64530, x64502, x64494);
  nand n64532(x64532, x64506, x64496);
  nand n64534(x64534, x64532, x64533);
  nand n64535(x64535, x64506, x64498);
  nand n64537(x64537, x64510, x64500);
  nand n64539(x64539, x64537, x64538);
  nand n64540(x64540, x64510, x64502);
  nand n64542(x64542, x64514, x64504);
  nand n64544(x64544, x64542, x64543);
  nand n64545(x64545, x64514, x64506);
  nand n64548(x64548, x64526, x64477);
  nand n64550(x64550, x64548, x64549);
  nand n64551(x64551, x64531, x64486);
  nand n64553(x64553, x64551, x64552);
  nand n64554(x64554, x64536, x64518);
  nand n64556(x64556, x64554, x64555);
  nand n64557(x64557, x64541, x64521);
  nand n64559(x64559, x64557, x64558);
  nand n64560(x64560, x64546, x64524);
  nand n64562(x64562, x64560, x64561);
  nand n64563(x64563, x64546, x64526);
  nand n64566(x64566, x64564, x64477);
  nand n64568(x64568, x64566, x64567);
  nand n64569(x64569, x64435, x64428);
  nand n64570(x64570, x64569, x64485);
  nand n64571(x64571, x64441, x64486);
  nand n64572(x64572, x64440, x64515);
  nand n64573(x64573, x64572, x64571);
  nand n64575(x64575, x64446, x64518);
  nand n64577(x64577, x64445, x64576);
  nand n64578(x64578, x64577, x64575);
  nand n64580(x64580, x64451, x64521);
  nand n64581(x64581, x64450, x64547);
  nand n64582(x64582, x64581, x64580);
  nand n64584(x64584, x64456, x64550);
  nand n64586(x64586, x64455, x64585);
  nand n64587(x64587, x64586, x64584);
  nand n64589(x64589, x64461, x64553);
  nand n64591(x64591, x64460, x64590);
  nand n64592(x64592, x64591, x64589);
  nand n64594(x64594, x64466, x64556);
  nand n64596(x64596, x64465, x64595);
  nand n64597(x64597, x64596, x64594);
  nand n64599(x64599, x64471, x64559);
  nand n64600(x64600, x64470, x64565);
  nand n64601(x64601, x64600, x64599);
  nand n64603(x64603, x64476, x64568);
  nand n64605(x64605, x64475, x64604);
  nand n64606(x64606, x64605, x64603);
  nand n64645(x64645, x64640, x64609);
  nand n64647(x64647, x64646, x64608);
  nand n64648(x64648, x64647, x64645);
  nand n64649(x64649, x64640, x64610);
  nand n64650(x64650, x64646, x64609);
  nand n64651(x64651, x64650, x64649);
  nand n64652(x64652, x64640, x64611);
  nand n64653(x64653, x64646, x64610);
  nand n64654(x64654, x64653, x64652);
  nand n64655(x64655, x64640, x64612);
  nand n64656(x64656, x64646, x64611);
  nand n64657(x64657, x64656, x64655);
  nand n64658(x64658, x64640, x64613);
  nand n64659(x64659, x64646, x64612);
  nand n64660(x64660, x64659, x64658);
  nand n64661(x64661, x64640, x64614);
  nand n64662(x64662, x64646, x64613);
  nand n64663(x64663, x64662, x64661);
  nand n64664(x64664, x64640, x64615);
  nand n64665(x64665, x64646, x64614);
  nand n64666(x64666, x64665, x64664);
  nand n64667(x64667, x64640, x64616);
  nand n64668(x64668, x64646, x64615);
  nand n64669(x64669, x64668, x64667);
  nand n64670(x64670, x64640, x64617);
  nand n64671(x64671, x64646, x64616);
  nand n64672(x64672, x64671, x64670);
  nand n64673(x64673, x64640, x64618);
  nand n64674(x64674, x64646, x64617);
  nand n64675(x64675, x64674, x64673);
  nand n64676(x64676, x64640, x64619);
  nand n64677(x64677, x64646, x64618);
  nand n64678(x64678, x64677, x64676);
  nand n64679(x64679, x64640, x64620);
  nand n64680(x64680, x64646, x64619);
  nand n64681(x64681, x64680, x64679);
  nand n64682(x64682, x64640, x64621);
  nand n64683(x64683, x64646, x64620);
  nand n64684(x64684, x64683, x64682);
  nand n64685(x64685, x64640, x64622);
  nand n64686(x64686, x64646, x64621);
  nand n64687(x64687, x64686, x64685);
  nand n64688(x64688, x64640, x64623);
  nand n64689(x64689, x64646, x64622);
  nand n64690(x64690, x64689, x64688);
  nand n64691(x64691, x64640, x64624);
  nand n64692(x64692, x64646, x64623);
  nand n64693(x64693, x64692, x64691);
  nand n64694(x64694, x64640, x64625);
  nand n64695(x64695, x64646, x64624);
  nand n64696(x64696, x64695, x64694);
  nand n64697(x64697, x64640, x64626);
  nand n64698(x64698, x64646, x64625);
  nand n64699(x64699, x64698, x64697);
  nand n64700(x64700, x64640, x64627);
  nand n64701(x64701, x64646, x64626);
  nand n64702(x64702, x64701, x64700);
  nand n64703(x64703, x64640, x64628);
  nand n64704(x64704, x64646, x64627);
  nand n64705(x64705, x64704, x64703);
  nand n64706(x64706, x64640, x64629);
  nand n64707(x64707, x64646, x64628);
  nand n64708(x64708, x64707, x64706);
  nand n64709(x64709, x64640, x64630);
  nand n64710(x64710, x64646, x64629);
  nand n64711(x64711, x64710, x64709);
  nand n64712(x64712, x64640, x64631);
  nand n64713(x64713, x64646, x64630);
  nand n64714(x64714, x64713, x64712);
  nand n64715(x64715, x64640, x64632);
  nand n64716(x64716, x64646, x64631);
  nand n64717(x64717, x64716, x64715);
  nand n64718(x64718, x64640, x64633);
  nand n64719(x64719, x64646, x64632);
  nand n64720(x64720, x64719, x64718);
  nand n64721(x64721, x64640, x64634);
  nand n64722(x64722, x64646, x64633);
  nand n64723(x64723, x64722, x64721);
  nand n64724(x64724, x64640, x64635);
  nand n64725(x64725, x64646, x64634);
  nand n64726(x64726, x64725, x64724);
  nand n64727(x64727, x64640, x64636);
  nand n64728(x64728, x64646, x64635);
  nand n64729(x64729, x64728, x64727);
  nand n64730(x64730, x64640, x64637);
  nand n64731(x64731, x64646, x64636);
  nand n64732(x64732, x64731, x64730);
  nand n64733(x64733, x64640, x64638);
  nand n64734(x64734, x64646, x64637);
  nand n64735(x64735, x64734, x64733);
  nand n64736(x64736, x64640, x64639);
  nand n64737(x64737, x64646, x64638);
  nand n64738(x64738, x64737, x64736);
  nand n64739(x64739, x64646, x64639);
  nand n64740(x64740, x64641, x64654);
  nand n64742(x64742, x64741, x64648);
  nand n64743(x64743, x64742, x64740);
  nand n64744(x64744, x64641, x64657);
  nand n64745(x64745, x64741, x64651);
  nand n64746(x64746, x64745, x64744);
  nand n64747(x64747, x64641, x64660);
  nand n64748(x64748, x64741, x64654);
  nand n64749(x64749, x64748, x64747);
  nand n64750(x64750, x64641, x64663);
  nand n64751(x64751, x64741, x64657);
  nand n64752(x64752, x64751, x64750);
  nand n64753(x64753, x64641, x64666);
  nand n64754(x64754, x64741, x64660);
  nand n64755(x64755, x64754, x64753);
  nand n64756(x64756, x64641, x64669);
  nand n64757(x64757, x64741, x64663);
  nand n64758(x64758, x64757, x64756);
  nand n64759(x64759, x64641, x64672);
  nand n64760(x64760, x64741, x64666);
  nand n64761(x64761, x64760, x64759);
  nand n64762(x64762, x64641, x64675);
  nand n64763(x64763, x64741, x64669);
  nand n64764(x64764, x64763, x64762);
  nand n64765(x64765, x64641, x64678);
  nand n64766(x64766, x64741, x64672);
  nand n64767(x64767, x64766, x64765);
  nand n64768(x64768, x64641, x64681);
  nand n64769(x64769, x64741, x64675);
  nand n64770(x64770, x64769, x64768);
  nand n64771(x64771, x64641, x64684);
  nand n64772(x64772, x64741, x64678);
  nand n64773(x64773, x64772, x64771);
  nand n64774(x64774, x64641, x64687);
  nand n64775(x64775, x64741, x64681);
  nand n64776(x64776, x64775, x64774);
  nand n64777(x64777, x64641, x64690);
  nand n64778(x64778, x64741, x64684);
  nand n64779(x64779, x64778, x64777);
  nand n64780(x64780, x64641, x64693);
  nand n64781(x64781, x64741, x64687);
  nand n64782(x64782, x64781, x64780);
  nand n64783(x64783, x64641, x64696);
  nand n64784(x64784, x64741, x64690);
  nand n64785(x64785, x64784, x64783);
  nand n64786(x64786, x64641, x64699);
  nand n64787(x64787, x64741, x64693);
  nand n64788(x64788, x64787, x64786);
  nand n64789(x64789, x64641, x64702);
  nand n64790(x64790, x64741, x64696);
  nand n64791(x64791, x64790, x64789);
  nand n64792(x64792, x64641, x64705);
  nand n64793(x64793, x64741, x64699);
  nand n64794(x64794, x64793, x64792);
  nand n64795(x64795, x64641, x64708);
  nand n64796(x64796, x64741, x64702);
  nand n64797(x64797, x64796, x64795);
  nand n64798(x64798, x64641, x64711);
  nand n64799(x64799, x64741, x64705);
  nand n64800(x64800, x64799, x64798);
  nand n64801(x64801, x64641, x64714);
  nand n64802(x64802, x64741, x64708);
  nand n64803(x64803, x64802, x64801);
  nand n64804(x64804, x64641, x64717);
  nand n64805(x64805, x64741, x64711);
  nand n64806(x64806, x64805, x64804);
  nand n64807(x64807, x64641, x64720);
  nand n64808(x64808, x64741, x64714);
  nand n64809(x64809, x64808, x64807);
  nand n64810(x64810, x64641, x64723);
  nand n64811(x64811, x64741, x64717);
  nand n64812(x64812, x64811, x64810);
  nand n64813(x64813, x64641, x64726);
  nand n64814(x64814, x64741, x64720);
  nand n64815(x64815, x64814, x64813);
  nand n64816(x64816, x64641, x64729);
  nand n64817(x64817, x64741, x64723);
  nand n64818(x64818, x64817, x64816);
  nand n64819(x64819, x64641, x64732);
  nand n64820(x64820, x64741, x64726);
  nand n64821(x64821, x64820, x64819);
  nand n64822(x64822, x64641, x64735);
  nand n64823(x64823, x64741, x64729);
  nand n64824(x64824, x64823, x64822);
  nand n64825(x64825, x64641, x64738);
  nand n64826(x64826, x64741, x64732);
  nand n64827(x64827, x64826, x64825);
  nand n64828(x64828, x64641, x86299);
  nand n64829(x64829, x64741, x64735);
  nand n64830(x64830, x64829, x64828);
  nand n64831(x64831, x64741, x64738);
  nand n64832(x64832, x64741, x86299);
  nand n64833(x64833, x64642, x64755);
  nand n64835(x64835, x64834, x64743);
  nand n64836(x64836, x64835, x64833);
  nand n64837(x64837, x64642, x64758);
  nand n64838(x64838, x64834, x64746);
  nand n64839(x64839, x64838, x64837);
  nand n64840(x64840, x64642, x64761);
  nand n64841(x64841, x64834, x64749);
  nand n64842(x64842, x64841, x64840);
  nand n64843(x64843, x64642, x64764);
  nand n64844(x64844, x64834, x64752);
  nand n64845(x64845, x64844, x64843);
  nand n64846(x64846, x64642, x64767);
  nand n64847(x64847, x64834, x64755);
  nand n64848(x64848, x64847, x64846);
  nand n64849(x64849, x64642, x64770);
  nand n64850(x64850, x64834, x64758);
  nand n64851(x64851, x64850, x64849);
  nand n64852(x64852, x64642, x64773);
  nand n64853(x64853, x64834, x64761);
  nand n64854(x64854, x64853, x64852);
  nand n64855(x64855, x64642, x64776);
  nand n64856(x64856, x64834, x64764);
  nand n64857(x64857, x64856, x64855);
  nand n64858(x64858, x64642, x64779);
  nand n64859(x64859, x64834, x64767);
  nand n64860(x64860, x64859, x64858);
  nand n64861(x64861, x64642, x64782);
  nand n64862(x64862, x64834, x64770);
  nand n64863(x64863, x64862, x64861);
  nand n64864(x64864, x64642, x64785);
  nand n64865(x64865, x64834, x64773);
  nand n64866(x64866, x64865, x64864);
  nand n64867(x64867, x64642, x64788);
  nand n64868(x64868, x64834, x64776);
  nand n64869(x64869, x64868, x64867);
  nand n64870(x64870, x64642, x64791);
  nand n64871(x64871, x64834, x64779);
  nand n64872(x64872, x64871, x64870);
  nand n64873(x64873, x64642, x64794);
  nand n64874(x64874, x64834, x64782);
  nand n64875(x64875, x64874, x64873);
  nand n64876(x64876, x64642, x64797);
  nand n64877(x64877, x64834, x64785);
  nand n64878(x64878, x64877, x64876);
  nand n64879(x64879, x64642, x64800);
  nand n64880(x64880, x64834, x64788);
  nand n64881(x64881, x64880, x64879);
  nand n64882(x64882, x64642, x64803);
  nand n64883(x64883, x64834, x64791);
  nand n64884(x64884, x64883, x64882);
  nand n64885(x64885, x64642, x64806);
  nand n64886(x64886, x64834, x64794);
  nand n64887(x64887, x64886, x64885);
  nand n64888(x64888, x64642, x64809);
  nand n64889(x64889, x64834, x64797);
  nand n64890(x64890, x64889, x64888);
  nand n64891(x64891, x64642, x64812);
  nand n64892(x64892, x64834, x64800);
  nand n64893(x64893, x64892, x64891);
  nand n64894(x64894, x64642, x64815);
  nand n64895(x64895, x64834, x64803);
  nand n64896(x64896, x64895, x64894);
  nand n64897(x64897, x64642, x64818);
  nand n64898(x64898, x64834, x64806);
  nand n64899(x64899, x64898, x64897);
  nand n64900(x64900, x64642, x64821);
  nand n64901(x64901, x64834, x64809);
  nand n64902(x64902, x64901, x64900);
  nand n64903(x64903, x64642, x64824);
  nand n64904(x64904, x64834, x64812);
  nand n64905(x64905, x64904, x64903);
  nand n64906(x64906, x64642, x64827);
  nand n64907(x64907, x64834, x64815);
  nand n64908(x64908, x64907, x64906);
  nand n64909(x64909, x64642, x64830);
  nand n64910(x64910, x64834, x64818);
  nand n64911(x64911, x64910, x64909);
  nand n64912(x64912, x64642, x86300);
  nand n64913(x64913, x64834, x64821);
  nand n64914(x64914, x64913, x64912);
  nand n64915(x64915, x64642, x86301);
  nand n64916(x64916, x64834, x64824);
  nand n64917(x64917, x64916, x64915);
  nand n64918(x64918, x64834, x64827);
  nand n64919(x64919, x64834, x64830);
  nand n64920(x64920, x64834, x86300);
  nand n64921(x64921, x64834, x86301);
  nand n64922(x64922, x64643, x64860);
  nand n64924(x64924, x64923, x64836);
  nand n64925(x64925, x64924, x64922);
  nand n64926(x64926, x64643, x64863);
  nand n64927(x64927, x64923, x64839);
  nand n64928(x64928, x64927, x64926);
  nand n64929(x64929, x64643, x64866);
  nand n64930(x64930, x64923, x64842);
  nand n64931(x64931, x64930, x64929);
  nand n64932(x64932, x64643, x64869);
  nand n64933(x64933, x64923, x64845);
  nand n64934(x64934, x64933, x64932);
  nand n64935(x64935, x64643, x64872);
  nand n64936(x64936, x64923, x64848);
  nand n64937(x64937, x64936, x64935);
  nand n64938(x64938, x64643, x64875);
  nand n64939(x64939, x64923, x64851);
  nand n64940(x64940, x64939, x64938);
  nand n64941(x64941, x64643, x64878);
  nand n64942(x64942, x64923, x64854);
  nand n64943(x64943, x64942, x64941);
  nand n64944(x64944, x64643, x64881);
  nand n64945(x64945, x64923, x64857);
  nand n64946(x64946, x64945, x64944);
  nand n64947(x64947, x64643, x64884);
  nand n64948(x64948, x64923, x64860);
  nand n64949(x64949, x64948, x64947);
  nand n64950(x64950, x64643, x64887);
  nand n64951(x64951, x64923, x64863);
  nand n64952(x64952, x64951, x64950);
  nand n64953(x64953, x64643, x64890);
  nand n64954(x64954, x64923, x64866);
  nand n64955(x64955, x64954, x64953);
  nand n64956(x64956, x64643, x64893);
  nand n64957(x64957, x64923, x64869);
  nand n64958(x64958, x64957, x64956);
  nand n64959(x64959, x64643, x64896);
  nand n64960(x64960, x64923, x64872);
  nand n64961(x64961, x64960, x64959);
  nand n64962(x64962, x64643, x64899);
  nand n64963(x64963, x64923, x64875);
  nand n64964(x64964, x64963, x64962);
  nand n64965(x64965, x64643, x64902);
  nand n64966(x64966, x64923, x64878);
  nand n64967(x64967, x64966, x64965);
  nand n64968(x64968, x64643, x64905);
  nand n64969(x64969, x64923, x64881);
  nand n64970(x64970, x64969, x64968);
  nand n64971(x64971, x64643, x64908);
  nand n64972(x64972, x64923, x64884);
  nand n64973(x64973, x64972, x64971);
  nand n64974(x64974, x64643, x64911);
  nand n64975(x64975, x64923, x64887);
  nand n64976(x64976, x64975, x64974);
  nand n64977(x64977, x64643, x64914);
  nand n64978(x64978, x64923, x64890);
  nand n64979(x64979, x64978, x64977);
  nand n64980(x64980, x64643, x64917);
  nand n64981(x64981, x64923, x64893);
  nand n64982(x64982, x64981, x64980);
  nand n64983(x64983, x64643, x86302);
  nand n64984(x64984, x64923, x64896);
  nand n64985(x64985, x64984, x64983);
  nand n64986(x64986, x64643, x86303);
  nand n64987(x64987, x64923, x64899);
  nand n64988(x64988, x64987, x64986);
  nand n64989(x64989, x64643, x86304);
  nand n64990(x64990, x64923, x64902);
  nand n64991(x64991, x64990, x64989);
  nand n64992(x64992, x64643, x86305);
  nand n64993(x64993, x64923, x64905);
  nand n64994(x64994, x64993, x64992);
  nand n64995(x64995, x64923, x64908);
  nand n64996(x64996, x64923, x64911);
  nand n64997(x64997, x64923, x64914);
  nand n64998(x64998, x64923, x64917);
  nand n64999(x64999, x64923, x86302);
  nand n65000(x65000, x64923, x86303);
  nand n65001(x65001, x64923, x86304);
  nand n65002(x65002, x64923, x86305);
  nand n65003(x65003, x64644, x64973);
  nand n65005(x65005, x65004, x64925);
  nand n65006(x65006, x65005, x65003);
  nand n65007(x65007, x64644, x64976);
  nand n65008(x65008, x65004, x64928);
  nand n65009(x65009, x65008, x65007);
  nand n65010(x65010, x64644, x64979);
  nand n65011(x65011, x65004, x64931);
  nand n65012(x65012, x65011, x65010);
  nand n65013(x65013, x64644, x64982);
  nand n65014(x65014, x65004, x64934);
  nand n65015(x65015, x65014, x65013);
  nand n65016(x65016, x64644, x64985);
  nand n65017(x65017, x65004, x64937);
  nand n65018(x65018, x65017, x65016);
  nand n65019(x65019, x64644, x64988);
  nand n65020(x65020, x65004, x64940);
  nand n65021(x65021, x65020, x65019);
  nand n65022(x65022, x64644, x64991);
  nand n65023(x65023, x65004, x64943);
  nand n65024(x65024, x65023, x65022);
  nand n65025(x65025, x64644, x64994);
  nand n65026(x65026, x65004, x64946);
  nand n65027(x65027, x65026, x65025);
  nand n65028(x65028, x64644, x86306);
  nand n65029(x65029, x65004, x64949);
  nand n65030(x65030, x65029, x65028);
  nand n65031(x65031, x64644, x86307);
  nand n65032(x65032, x65004, x64952);
  nand n65033(x65033, x65032, x65031);
  nand n65034(x65034, x64644, x86308);
  nand n65035(x65035, x65004, x64955);
  nand n65036(x65036, x65035, x65034);
  nand n65037(x65037, x64644, x86309);
  nand n65038(x65038, x65004, x64958);
  nand n65039(x65039, x65038, x65037);
  nand n65040(x65040, x64644, x86310);
  nand n65041(x65041, x65004, x64961);
  nand n65042(x65042, x65041, x65040);
  nand n65043(x65043, x64644, x86311);
  nand n65044(x65044, x65004, x64964);
  nand n65045(x65045, x65044, x65043);
  nand n65046(x65046, x64644, x86312);
  nand n65047(x65047, x65004, x64967);
  nand n65048(x65048, x65047, x65046);
  nand n65049(x65049, x64644, x86313);
  nand n65050(x65050, x65004, x64970);
  nand n65051(x65051, x65050, x65049);
  nand n65052(x65052, x65004, x64973);
  nand n65053(x65053, x65004, x64976);
  nand n65054(x65054, x65004, x64979);
  nand n65055(x65055, x65004, x64982);
  nand n65056(x65056, x65004, x64985);
  nand n65057(x65057, x65004, x64988);
  nand n65058(x65058, x65004, x64991);
  nand n65059(x65059, x65004, x64994);
  nand n65060(x65060, x65004, x86306);
  nand n65061(x65061, x65004, x86307);
  nand n65062(x65062, x65004, x86308);
  nand n65063(x65063, x65004, x86309);
  nand n65064(x65064, x65004, x86310);
  nand n65065(x65065, x65004, x86311);
  nand n65066(x65066, x65004, x86312);
  nand n65067(x65067, x65004, x86313);
  nand n65068(x65068, x76792, x77422);
  nand n65069(x65069, x62933, x77518);
  nand n65070(x65070, x65069, x65068);
  nand n65071(x65071, x76792, x77425);
  nand n65072(x65072, x62933, x77521);
  nand n65073(x65073, x65072, x65071);
  nand n65074(x65074, x76792, x77428);
  nand n65075(x65075, x62933, x77524);
  nand n65076(x65076, x65075, x65074);
  nand n65077(x65077, x76792, x77431);
  nand n65078(x65078, x62933, x77527);
  nand n65079(x65079, x65078, x65077);
  nand n65080(x65080, x76792, x77434);
  nand n65081(x65081, x62933, x77530);
  nand n65082(x65082, x65081, x65080);
  nand n65083(x65083, x76792, x77437);
  nand n65084(x65084, x62933, x77533);
  nand n65085(x65085, x65084, x65083);
  nand n65086(x65086, x76792, x77440);
  nand n65087(x65087, x62933, x77536);
  nand n65088(x65088, x65087, x65086);
  nand n65089(x65089, x76792, x77443);
  nand n65090(x65090, x62933, x77539);
  nand n65091(x65091, x65090, x65089);
  nand n65092(x65092, x76792, x77446);
  nand n65093(x65093, x62933, x77542);
  nand n65094(x65094, x65093, x65092);
  nand n65095(x65095, x76792, x77449);
  nand n65096(x65096, x62933, x77545);
  nand n65097(x65097, x65096, x65095);
  nand n65098(x65098, x76675, x65070);
  nand n65100(x65100, x63028, x65099);
  nand n65101(x65101, x65100, x65098);
  nand n65102(x65102, x76678, x65073);
  nand n65104(x65104, x63033, x65103);
  nand n65105(x65105, x65104, x65102);
  nand n65107(x65107, x76681, x65076);
  nand n65109(x65109, x63039, x65108);
  nand n65110(x65110, x65109, x65107);
  nand n65112(x65112, x76684, x65079);
  nand n65114(x65114, x63045, x65113);
  nand n65115(x65115, x65114, x65112);
  nand n65117(x65117, x76687, x65082);
  nand n65119(x65119, x63051, x65118);
  nand n65120(x65120, x65119, x65117);
  nand n65122(x65122, x76690, x65085);
  nand n65124(x65124, x63057, x65123);
  nand n65125(x65125, x65124, x65122);
  nand n65127(x65127, x76693, x65088);
  nand n65129(x65129, x63063, x65128);
  nand n65130(x65130, x65129, x65127);
  nand n65132(x65132, x76696, x65091);
  nand n65134(x65134, x63069, x65133);
  nand n65135(x65135, x65134, x65132);
  nand n65137(x65137, x76699, x65094);
  nand n65139(x65139, x63075, x65138);
  nand n65140(x65140, x65139, x65137);
  nand n65142(x65142, x76702, x65097);
  nand n65144(x65144, x63081, x65143);
  nand n65145(x65145, x65144, x65142);
  nand n65155(x65155, x65106, x65147);
  nand n65156(x65156, x65155, x65102);
  nand n65157(x65157, x65111, x65148);
  nand n65158(x65158, x65157, x65107);
  nand n65159(x65159, x65111, x65106);
  nand n65161(x65161, x65116, x65149);
  nand n65162(x65162, x65161, x65112);
  nand n65163(x65163, x65116, x65111);
  nand n65165(x65165, x65121, x65150);
  nand n65166(x65166, x65165, x65117);
  nand n65167(x65167, x65121, x65116);
  nand n65169(x65169, x65126, x65151);
  nand n65170(x65170, x65169, x65122);
  nand n65171(x65171, x65126, x65121);
  nand n65173(x65173, x65131, x65152);
  nand n65174(x65174, x65173, x65127);
  nand n65175(x65175, x65131, x65126);
  nand n65177(x65177, x65136, x65153);
  nand n65178(x65178, x65177, x65132);
  nand n65179(x65179, x65136, x65131);
  nand n65181(x65181, x65141, x65154);
  nand n65182(x65182, x65181, x65137);
  nand n65183(x65183, x65141, x65136);
  nand n65186(x65186, x65160, x65147);
  nand n65188(x65188, x65186, x65187);
  nand n65189(x65189, x65164, x65156);
  nand n65191(x65191, x65189, x65190);
  nand n65192(x65192, x65168, x65158);
  nand n65194(x65194, x65192, x65193);
  nand n65195(x65195, x65168, x65160);
  nand n65197(x65197, x65172, x65162);
  nand n65199(x65199, x65197, x65198);
  nand n65200(x65200, x65172, x65164);
  nand n65202(x65202, x65176, x65166);
  nand n65204(x65204, x65202, x65203);
  nand n65205(x65205, x65176, x65168);
  nand n65207(x65207, x65180, x65170);
  nand n65209(x65209, x65207, x65208);
  nand n65210(x65210, x65180, x65172);
  nand n65212(x65212, x65184, x65174);
  nand n65214(x65214, x65212, x65213);
  nand n65215(x65215, x65184, x65176);
  nand n65218(x65218, x65196, x65147);
  nand n65220(x65220, x65218, x65219);
  nand n65221(x65221, x65201, x65156);
  nand n65223(x65223, x65221, x65222);
  nand n65224(x65224, x65206, x65188);
  nand n65226(x65226, x65224, x65225);
  nand n65227(x65227, x65211, x65191);
  nand n65229(x65229, x65227, x65228);
  nand n65230(x65230, x65216, x65194);
  nand n65232(x65232, x65230, x65231);
  nand n65233(x65233, x65216, x65196);
  nand n65236(x65236, x65234, x65147);
  nand n65238(x65238, x65236, x65237);
  nand n65239(x65239, x65105, x65098);
  nand n65240(x65240, x65239, x65155);
  nand n65241(x65241, x65111, x65156);
  nand n65242(x65242, x65110, x65185);
  nand n65243(x65243, x65242, x65241);
  nand n65245(x65245, x65116, x65188);
  nand n65247(x65247, x65115, x65246);
  nand n65248(x65248, x65247, x65245);
  nand n65250(x65250, x65121, x65191);
  nand n65251(x65251, x65120, x65217);
  nand n65252(x65252, x65251, x65250);
  nand n65254(x65254, x65126, x65220);
  nand n65256(x65256, x65125, x65255);
  nand n65257(x65257, x65256, x65254);
  nand n65259(x65259, x65131, x65223);
  nand n65261(x65261, x65130, x65260);
  nand n65262(x65262, x65261, x65259);
  nand n65264(x65264, x65136, x65226);
  nand n65266(x65266, x65135, x65265);
  nand n65267(x65267, x65266, x65264);
  nand n65269(x65269, x65141, x65229);
  nand n65270(x65270, x65140, x65235);
  nand n65271(x65271, x65270, x65269);
  nand n65273(x65273, x65146, x65238);
  nand n65275(x65275, x65145, x65274);
  nand n65276(x65276, x65275, x65273);
  nand n65315(x65315, x65310, x65279);
  nand n65317(x65317, x65316, x65278);
  nand n65318(x65318, x65317, x65315);
  nand n65319(x65319, x65310, x65280);
  nand n65320(x65320, x65316, x65279);
  nand n65321(x65321, x65320, x65319);
  nand n65322(x65322, x65310, x65281);
  nand n65323(x65323, x65316, x65280);
  nand n65324(x65324, x65323, x65322);
  nand n65325(x65325, x65310, x65282);
  nand n65326(x65326, x65316, x65281);
  nand n65327(x65327, x65326, x65325);
  nand n65328(x65328, x65310, x65283);
  nand n65329(x65329, x65316, x65282);
  nand n65330(x65330, x65329, x65328);
  nand n65331(x65331, x65310, x65284);
  nand n65332(x65332, x65316, x65283);
  nand n65333(x65333, x65332, x65331);
  nand n65334(x65334, x65310, x65285);
  nand n65335(x65335, x65316, x65284);
  nand n65336(x65336, x65335, x65334);
  nand n65337(x65337, x65310, x65286);
  nand n65338(x65338, x65316, x65285);
  nand n65339(x65339, x65338, x65337);
  nand n65340(x65340, x65310, x65287);
  nand n65341(x65341, x65316, x65286);
  nand n65342(x65342, x65341, x65340);
  nand n65343(x65343, x65310, x65288);
  nand n65344(x65344, x65316, x65287);
  nand n65345(x65345, x65344, x65343);
  nand n65346(x65346, x65310, x65289);
  nand n65347(x65347, x65316, x65288);
  nand n65348(x65348, x65347, x65346);
  nand n65349(x65349, x65310, x65290);
  nand n65350(x65350, x65316, x65289);
  nand n65351(x65351, x65350, x65349);
  nand n65352(x65352, x65310, x65291);
  nand n65353(x65353, x65316, x65290);
  nand n65354(x65354, x65353, x65352);
  nand n65355(x65355, x65310, x65292);
  nand n65356(x65356, x65316, x65291);
  nand n65357(x65357, x65356, x65355);
  nand n65358(x65358, x65310, x65293);
  nand n65359(x65359, x65316, x65292);
  nand n65360(x65360, x65359, x65358);
  nand n65361(x65361, x65310, x65294);
  nand n65362(x65362, x65316, x65293);
  nand n65363(x65363, x65362, x65361);
  nand n65364(x65364, x65310, x65295);
  nand n65365(x65365, x65316, x65294);
  nand n65366(x65366, x65365, x65364);
  nand n65367(x65367, x65310, x65296);
  nand n65368(x65368, x65316, x65295);
  nand n65369(x65369, x65368, x65367);
  nand n65370(x65370, x65310, x65297);
  nand n65371(x65371, x65316, x65296);
  nand n65372(x65372, x65371, x65370);
  nand n65373(x65373, x65310, x65298);
  nand n65374(x65374, x65316, x65297);
  nand n65375(x65375, x65374, x65373);
  nand n65376(x65376, x65310, x65299);
  nand n65377(x65377, x65316, x65298);
  nand n65378(x65378, x65377, x65376);
  nand n65379(x65379, x65310, x65300);
  nand n65380(x65380, x65316, x65299);
  nand n65381(x65381, x65380, x65379);
  nand n65382(x65382, x65310, x65301);
  nand n65383(x65383, x65316, x65300);
  nand n65384(x65384, x65383, x65382);
  nand n65385(x65385, x65310, x65302);
  nand n65386(x65386, x65316, x65301);
  nand n65387(x65387, x65386, x65385);
  nand n65388(x65388, x65310, x65303);
  nand n65389(x65389, x65316, x65302);
  nand n65390(x65390, x65389, x65388);
  nand n65391(x65391, x65310, x65304);
  nand n65392(x65392, x65316, x65303);
  nand n65393(x65393, x65392, x65391);
  nand n65394(x65394, x65310, x65305);
  nand n65395(x65395, x65316, x65304);
  nand n65396(x65396, x65395, x65394);
  nand n65397(x65397, x65310, x65306);
  nand n65398(x65398, x65316, x65305);
  nand n65399(x65399, x65398, x65397);
  nand n65400(x65400, x65310, x65307);
  nand n65401(x65401, x65316, x65306);
  nand n65402(x65402, x65401, x65400);
  nand n65403(x65403, x65310, x65308);
  nand n65404(x65404, x65316, x65307);
  nand n65405(x65405, x65404, x65403);
  nand n65406(x65406, x65310, x65309);
  nand n65407(x65407, x65316, x65308);
  nand n65408(x65408, x65407, x65406);
  nand n65409(x65409, x65316, x65309);
  nand n65410(x65410, x65311, x65324);
  nand n65412(x65412, x65411, x65318);
  nand n65413(x65413, x65412, x65410);
  nand n65414(x65414, x65311, x65327);
  nand n65415(x65415, x65411, x65321);
  nand n65416(x65416, x65415, x65414);
  nand n65417(x65417, x65311, x65330);
  nand n65418(x65418, x65411, x65324);
  nand n65419(x65419, x65418, x65417);
  nand n65420(x65420, x65311, x65333);
  nand n65421(x65421, x65411, x65327);
  nand n65422(x65422, x65421, x65420);
  nand n65423(x65423, x65311, x65336);
  nand n65424(x65424, x65411, x65330);
  nand n65425(x65425, x65424, x65423);
  nand n65426(x65426, x65311, x65339);
  nand n65427(x65427, x65411, x65333);
  nand n65428(x65428, x65427, x65426);
  nand n65429(x65429, x65311, x65342);
  nand n65430(x65430, x65411, x65336);
  nand n65431(x65431, x65430, x65429);
  nand n65432(x65432, x65311, x65345);
  nand n65433(x65433, x65411, x65339);
  nand n65434(x65434, x65433, x65432);
  nand n65435(x65435, x65311, x65348);
  nand n65436(x65436, x65411, x65342);
  nand n65437(x65437, x65436, x65435);
  nand n65438(x65438, x65311, x65351);
  nand n65439(x65439, x65411, x65345);
  nand n65440(x65440, x65439, x65438);
  nand n65441(x65441, x65311, x65354);
  nand n65442(x65442, x65411, x65348);
  nand n65443(x65443, x65442, x65441);
  nand n65444(x65444, x65311, x65357);
  nand n65445(x65445, x65411, x65351);
  nand n65446(x65446, x65445, x65444);
  nand n65447(x65447, x65311, x65360);
  nand n65448(x65448, x65411, x65354);
  nand n65449(x65449, x65448, x65447);
  nand n65450(x65450, x65311, x65363);
  nand n65451(x65451, x65411, x65357);
  nand n65452(x65452, x65451, x65450);
  nand n65453(x65453, x65311, x65366);
  nand n65454(x65454, x65411, x65360);
  nand n65455(x65455, x65454, x65453);
  nand n65456(x65456, x65311, x65369);
  nand n65457(x65457, x65411, x65363);
  nand n65458(x65458, x65457, x65456);
  nand n65459(x65459, x65311, x65372);
  nand n65460(x65460, x65411, x65366);
  nand n65461(x65461, x65460, x65459);
  nand n65462(x65462, x65311, x65375);
  nand n65463(x65463, x65411, x65369);
  nand n65464(x65464, x65463, x65462);
  nand n65465(x65465, x65311, x65378);
  nand n65466(x65466, x65411, x65372);
  nand n65467(x65467, x65466, x65465);
  nand n65468(x65468, x65311, x65381);
  nand n65469(x65469, x65411, x65375);
  nand n65470(x65470, x65469, x65468);
  nand n65471(x65471, x65311, x65384);
  nand n65472(x65472, x65411, x65378);
  nand n65473(x65473, x65472, x65471);
  nand n65474(x65474, x65311, x65387);
  nand n65475(x65475, x65411, x65381);
  nand n65476(x65476, x65475, x65474);
  nand n65477(x65477, x65311, x65390);
  nand n65478(x65478, x65411, x65384);
  nand n65479(x65479, x65478, x65477);
  nand n65480(x65480, x65311, x65393);
  nand n65481(x65481, x65411, x65387);
  nand n65482(x65482, x65481, x65480);
  nand n65483(x65483, x65311, x65396);
  nand n65484(x65484, x65411, x65390);
  nand n65485(x65485, x65484, x65483);
  nand n65486(x65486, x65311, x65399);
  nand n65487(x65487, x65411, x65393);
  nand n65488(x65488, x65487, x65486);
  nand n65489(x65489, x65311, x65402);
  nand n65490(x65490, x65411, x65396);
  nand n65491(x65491, x65490, x65489);
  nand n65492(x65492, x65311, x65405);
  nand n65493(x65493, x65411, x65399);
  nand n65494(x65494, x65493, x65492);
  nand n65495(x65495, x65311, x65408);
  nand n65496(x65496, x65411, x65402);
  nand n65497(x65497, x65496, x65495);
  nand n65498(x65498, x65311, x86332);
  nand n65499(x65499, x65411, x65405);
  nand n65500(x65500, x65499, x65498);
  nand n65501(x65501, x65411, x65408);
  nand n65502(x65502, x65411, x86332);
  nand n65503(x65503, x65312, x65425);
  nand n65505(x65505, x65504, x65413);
  nand n65506(x65506, x65505, x65503);
  nand n65507(x65507, x65312, x65428);
  nand n65508(x65508, x65504, x65416);
  nand n65509(x65509, x65508, x65507);
  nand n65510(x65510, x65312, x65431);
  nand n65511(x65511, x65504, x65419);
  nand n65512(x65512, x65511, x65510);
  nand n65513(x65513, x65312, x65434);
  nand n65514(x65514, x65504, x65422);
  nand n65515(x65515, x65514, x65513);
  nand n65516(x65516, x65312, x65437);
  nand n65517(x65517, x65504, x65425);
  nand n65518(x65518, x65517, x65516);
  nand n65519(x65519, x65312, x65440);
  nand n65520(x65520, x65504, x65428);
  nand n65521(x65521, x65520, x65519);
  nand n65522(x65522, x65312, x65443);
  nand n65523(x65523, x65504, x65431);
  nand n65524(x65524, x65523, x65522);
  nand n65525(x65525, x65312, x65446);
  nand n65526(x65526, x65504, x65434);
  nand n65527(x65527, x65526, x65525);
  nand n65528(x65528, x65312, x65449);
  nand n65529(x65529, x65504, x65437);
  nand n65530(x65530, x65529, x65528);
  nand n65531(x65531, x65312, x65452);
  nand n65532(x65532, x65504, x65440);
  nand n65533(x65533, x65532, x65531);
  nand n65534(x65534, x65312, x65455);
  nand n65535(x65535, x65504, x65443);
  nand n65536(x65536, x65535, x65534);
  nand n65537(x65537, x65312, x65458);
  nand n65538(x65538, x65504, x65446);
  nand n65539(x65539, x65538, x65537);
  nand n65540(x65540, x65312, x65461);
  nand n65541(x65541, x65504, x65449);
  nand n65542(x65542, x65541, x65540);
  nand n65543(x65543, x65312, x65464);
  nand n65544(x65544, x65504, x65452);
  nand n65545(x65545, x65544, x65543);
  nand n65546(x65546, x65312, x65467);
  nand n65547(x65547, x65504, x65455);
  nand n65548(x65548, x65547, x65546);
  nand n65549(x65549, x65312, x65470);
  nand n65550(x65550, x65504, x65458);
  nand n65551(x65551, x65550, x65549);
  nand n65552(x65552, x65312, x65473);
  nand n65553(x65553, x65504, x65461);
  nand n65554(x65554, x65553, x65552);
  nand n65555(x65555, x65312, x65476);
  nand n65556(x65556, x65504, x65464);
  nand n65557(x65557, x65556, x65555);
  nand n65558(x65558, x65312, x65479);
  nand n65559(x65559, x65504, x65467);
  nand n65560(x65560, x65559, x65558);
  nand n65561(x65561, x65312, x65482);
  nand n65562(x65562, x65504, x65470);
  nand n65563(x65563, x65562, x65561);
  nand n65564(x65564, x65312, x65485);
  nand n65565(x65565, x65504, x65473);
  nand n65566(x65566, x65565, x65564);
  nand n65567(x65567, x65312, x65488);
  nand n65568(x65568, x65504, x65476);
  nand n65569(x65569, x65568, x65567);
  nand n65570(x65570, x65312, x65491);
  nand n65571(x65571, x65504, x65479);
  nand n65572(x65572, x65571, x65570);
  nand n65573(x65573, x65312, x65494);
  nand n65574(x65574, x65504, x65482);
  nand n65575(x65575, x65574, x65573);
  nand n65576(x65576, x65312, x65497);
  nand n65577(x65577, x65504, x65485);
  nand n65578(x65578, x65577, x65576);
  nand n65579(x65579, x65312, x65500);
  nand n65580(x65580, x65504, x65488);
  nand n65581(x65581, x65580, x65579);
  nand n65582(x65582, x65312, x86333);
  nand n65583(x65583, x65504, x65491);
  nand n65584(x65584, x65583, x65582);
  nand n65585(x65585, x65312, x86334);
  nand n65586(x65586, x65504, x65494);
  nand n65587(x65587, x65586, x65585);
  nand n65588(x65588, x65504, x65497);
  nand n65589(x65589, x65504, x65500);
  nand n65590(x65590, x65504, x86333);
  nand n65591(x65591, x65504, x86334);
  nand n65592(x65592, x65313, x65530);
  nand n65594(x65594, x65593, x65506);
  nand n65595(x65595, x65594, x65592);
  nand n65596(x65596, x65313, x65533);
  nand n65597(x65597, x65593, x65509);
  nand n65598(x65598, x65597, x65596);
  nand n65599(x65599, x65313, x65536);
  nand n65600(x65600, x65593, x65512);
  nand n65601(x65601, x65600, x65599);
  nand n65602(x65602, x65313, x65539);
  nand n65603(x65603, x65593, x65515);
  nand n65604(x65604, x65603, x65602);
  nand n65605(x65605, x65313, x65542);
  nand n65606(x65606, x65593, x65518);
  nand n65607(x65607, x65606, x65605);
  nand n65608(x65608, x65313, x65545);
  nand n65609(x65609, x65593, x65521);
  nand n65610(x65610, x65609, x65608);
  nand n65611(x65611, x65313, x65548);
  nand n65612(x65612, x65593, x65524);
  nand n65613(x65613, x65612, x65611);
  nand n65614(x65614, x65313, x65551);
  nand n65615(x65615, x65593, x65527);
  nand n65616(x65616, x65615, x65614);
  nand n65617(x65617, x65313, x65554);
  nand n65618(x65618, x65593, x65530);
  nand n65619(x65619, x65618, x65617);
  nand n65620(x65620, x65313, x65557);
  nand n65621(x65621, x65593, x65533);
  nand n65622(x65622, x65621, x65620);
  nand n65623(x65623, x65313, x65560);
  nand n65624(x65624, x65593, x65536);
  nand n65625(x65625, x65624, x65623);
  nand n65626(x65626, x65313, x65563);
  nand n65627(x65627, x65593, x65539);
  nand n65628(x65628, x65627, x65626);
  nand n65629(x65629, x65313, x65566);
  nand n65630(x65630, x65593, x65542);
  nand n65631(x65631, x65630, x65629);
  nand n65632(x65632, x65313, x65569);
  nand n65633(x65633, x65593, x65545);
  nand n65634(x65634, x65633, x65632);
  nand n65635(x65635, x65313, x65572);
  nand n65636(x65636, x65593, x65548);
  nand n65637(x65637, x65636, x65635);
  nand n65638(x65638, x65313, x65575);
  nand n65639(x65639, x65593, x65551);
  nand n65640(x65640, x65639, x65638);
  nand n65641(x65641, x65313, x65578);
  nand n65642(x65642, x65593, x65554);
  nand n65643(x65643, x65642, x65641);
  nand n65644(x65644, x65313, x65581);
  nand n65645(x65645, x65593, x65557);
  nand n65646(x65646, x65645, x65644);
  nand n65647(x65647, x65313, x65584);
  nand n65648(x65648, x65593, x65560);
  nand n65649(x65649, x65648, x65647);
  nand n65650(x65650, x65313, x65587);
  nand n65651(x65651, x65593, x65563);
  nand n65652(x65652, x65651, x65650);
  nand n65653(x65653, x65313, x86335);
  nand n65654(x65654, x65593, x65566);
  nand n65655(x65655, x65654, x65653);
  nand n65656(x65656, x65313, x86336);
  nand n65657(x65657, x65593, x65569);
  nand n65658(x65658, x65657, x65656);
  nand n65659(x65659, x65313, x86337);
  nand n65660(x65660, x65593, x65572);
  nand n65661(x65661, x65660, x65659);
  nand n65662(x65662, x65313, x86338);
  nand n65663(x65663, x65593, x65575);
  nand n65664(x65664, x65663, x65662);
  nand n65665(x65665, x65593, x65578);
  nand n65666(x65666, x65593, x65581);
  nand n65667(x65667, x65593, x65584);
  nand n65668(x65668, x65593, x65587);
  nand n65669(x65669, x65593, x86335);
  nand n65670(x65670, x65593, x86336);
  nand n65671(x65671, x65593, x86337);
  nand n65672(x65672, x65593, x86338);
  nand n65673(x65673, x65314, x65643);
  nand n65675(x65675, x65674, x65595);
  nand n65676(x65676, x65675, x65673);
  nand n65677(x65677, x65314, x65646);
  nand n65678(x65678, x65674, x65598);
  nand n65679(x65679, x65678, x65677);
  nand n65680(x65680, x65314, x65649);
  nand n65681(x65681, x65674, x65601);
  nand n65682(x65682, x65681, x65680);
  nand n65683(x65683, x65314, x65652);
  nand n65684(x65684, x65674, x65604);
  nand n65685(x65685, x65684, x65683);
  nand n65686(x65686, x65314, x65655);
  nand n65687(x65687, x65674, x65607);
  nand n65688(x65688, x65687, x65686);
  nand n65689(x65689, x65314, x65658);
  nand n65690(x65690, x65674, x65610);
  nand n65691(x65691, x65690, x65689);
  nand n65692(x65692, x65314, x65661);
  nand n65693(x65693, x65674, x65613);
  nand n65694(x65694, x65693, x65692);
  nand n65695(x65695, x65314, x65664);
  nand n65696(x65696, x65674, x65616);
  nand n65697(x65697, x65696, x65695);
  nand n65698(x65698, x65314, x86339);
  nand n65699(x65699, x65674, x65619);
  nand n65700(x65700, x65699, x65698);
  nand n65701(x65701, x65314, x86340);
  nand n65702(x65702, x65674, x65622);
  nand n65703(x65703, x65702, x65701);
  nand n65704(x65704, x65314, x86341);
  nand n65705(x65705, x65674, x65625);
  nand n65706(x65706, x65705, x65704);
  nand n65707(x65707, x65314, x86342);
  nand n65708(x65708, x65674, x65628);
  nand n65709(x65709, x65708, x65707);
  nand n65710(x65710, x65314, x86343);
  nand n65711(x65711, x65674, x65631);
  nand n65712(x65712, x65711, x65710);
  nand n65713(x65713, x65314, x86344);
  nand n65714(x65714, x65674, x65634);
  nand n65715(x65715, x65714, x65713);
  nand n65716(x65716, x65314, x86345);
  nand n65717(x65717, x65674, x65637);
  nand n65718(x65718, x65717, x65716);
  nand n65719(x65719, x65314, x86346);
  nand n65720(x65720, x65674, x65640);
  nand n65721(x65721, x65720, x65719);
  nand n65722(x65722, x65674, x65643);
  nand n65723(x65723, x65674, x65646);
  nand n65724(x65724, x65674, x65649);
  nand n65725(x65725, x65674, x65652);
  nand n65726(x65726, x65674, x65655);
  nand n65727(x65727, x65674, x65658);
  nand n65728(x65728, x65674, x65661);
  nand n65729(x65729, x65674, x65664);
  nand n65730(x65730, x65674, x86339);
  nand n65731(x65731, x65674, x86340);
  nand n65732(x65732, x65674, x86341);
  nand n65733(x65733, x65674, x86342);
  nand n65734(x65734, x65674, x86343);
  nand n65735(x65735, x65674, x86344);
  nand n65736(x65736, x65674, x86345);
  nand n65737(x65737, x65674, x86346);
  nand n65738(x65738, x76792, x77716);
  nand n65739(x65739, x62933, x77812);
  nand n65740(x65740, x65739, x65738);
  nand n65741(x65741, x76792, x77719);
  nand n65742(x65742, x62933, x77815);
  nand n65743(x65743, x65742, x65741);
  nand n65744(x65744, x76792, x77722);
  nand n65745(x65745, x62933, x77818);
  nand n65746(x65746, x65745, x65744);
  nand n65747(x65747, x76792, x77725);
  nand n65748(x65748, x62933, x77821);
  nand n65749(x65749, x65748, x65747);
  nand n65750(x65750, x76792, x77728);
  nand n65751(x65751, x62933, x77824);
  nand n65752(x65752, x65751, x65750);
  nand n65753(x65753, x76792, x77731);
  nand n65754(x65754, x62933, x77827);
  nand n65755(x65755, x65754, x65753);
  nand n65756(x65756, x76792, x77734);
  nand n65757(x65757, x62933, x77830);
  nand n65758(x65758, x65757, x65756);
  nand n65759(x65759, x76792, x77737);
  nand n65760(x65760, x62933, x77833);
  nand n65761(x65761, x65760, x65759);
  nand n65762(x65762, x76792, x77740);
  nand n65763(x65763, x62933, x77836);
  nand n65764(x65764, x65763, x65762);
  nand n65765(x65765, x76792, x77743);
  nand n65766(x65766, x62933, x77839);
  nand n65767(x65767, x65766, x65765);
  nand n65768(x65768, x76675, x65740);
  nand n65770(x65770, x63028, x65769);
  nand n65771(x65771, x65770, x65768);
  nand n65772(x65772, x76678, x65743);
  nand n65774(x65774, x63033, x65773);
  nand n65775(x65775, x65774, x65772);
  nand n65777(x65777, x76681, x65746);
  nand n65779(x65779, x63039, x65778);
  nand n65780(x65780, x65779, x65777);
  nand n65782(x65782, x76684, x65749);
  nand n65784(x65784, x63045, x65783);
  nand n65785(x65785, x65784, x65782);
  nand n65787(x65787, x76687, x65752);
  nand n65789(x65789, x63051, x65788);
  nand n65790(x65790, x65789, x65787);
  nand n65792(x65792, x76690, x65755);
  nand n65794(x65794, x63057, x65793);
  nand n65795(x65795, x65794, x65792);
  nand n65797(x65797, x76693, x65758);
  nand n65799(x65799, x63063, x65798);
  nand n65800(x65800, x65799, x65797);
  nand n65802(x65802, x76696, x65761);
  nand n65804(x65804, x63069, x65803);
  nand n65805(x65805, x65804, x65802);
  nand n65807(x65807, x76699, x65764);
  nand n65809(x65809, x63075, x65808);
  nand n65810(x65810, x65809, x65807);
  nand n65812(x65812, x76702, x65767);
  nand n65814(x65814, x63081, x65813);
  nand n65815(x65815, x65814, x65812);
  nand n65825(x65825, x65776, x65817);
  nand n65826(x65826, x65825, x65772);
  nand n65827(x65827, x65781, x65818);
  nand n65828(x65828, x65827, x65777);
  nand n65829(x65829, x65781, x65776);
  nand n65831(x65831, x65786, x65819);
  nand n65832(x65832, x65831, x65782);
  nand n65833(x65833, x65786, x65781);
  nand n65835(x65835, x65791, x65820);
  nand n65836(x65836, x65835, x65787);
  nand n65837(x65837, x65791, x65786);
  nand n65839(x65839, x65796, x65821);
  nand n65840(x65840, x65839, x65792);
  nand n65841(x65841, x65796, x65791);
  nand n65843(x65843, x65801, x65822);
  nand n65844(x65844, x65843, x65797);
  nand n65845(x65845, x65801, x65796);
  nand n65847(x65847, x65806, x65823);
  nand n65848(x65848, x65847, x65802);
  nand n65849(x65849, x65806, x65801);
  nand n65851(x65851, x65811, x65824);
  nand n65852(x65852, x65851, x65807);
  nand n65853(x65853, x65811, x65806);
  nand n65856(x65856, x65830, x65817);
  nand n65858(x65858, x65856, x65857);
  nand n65859(x65859, x65834, x65826);
  nand n65861(x65861, x65859, x65860);
  nand n65862(x65862, x65838, x65828);
  nand n65864(x65864, x65862, x65863);
  nand n65865(x65865, x65838, x65830);
  nand n65867(x65867, x65842, x65832);
  nand n65869(x65869, x65867, x65868);
  nand n65870(x65870, x65842, x65834);
  nand n65872(x65872, x65846, x65836);
  nand n65874(x65874, x65872, x65873);
  nand n65875(x65875, x65846, x65838);
  nand n65877(x65877, x65850, x65840);
  nand n65879(x65879, x65877, x65878);
  nand n65880(x65880, x65850, x65842);
  nand n65882(x65882, x65854, x65844);
  nand n65884(x65884, x65882, x65883);
  nand n65885(x65885, x65854, x65846);
  nand n65888(x65888, x65866, x65817);
  nand n65890(x65890, x65888, x65889);
  nand n65891(x65891, x65871, x65826);
  nand n65893(x65893, x65891, x65892);
  nand n65894(x65894, x65876, x65858);
  nand n65896(x65896, x65894, x65895);
  nand n65897(x65897, x65881, x65861);
  nand n65899(x65899, x65897, x65898);
  nand n65900(x65900, x65886, x65864);
  nand n65902(x65902, x65900, x65901);
  nand n65903(x65903, x65886, x65866);
  nand n65906(x65906, x65904, x65817);
  nand n65908(x65908, x65906, x65907);
  nand n65909(x65909, x65775, x65768);
  nand n65910(x65910, x65909, x65825);
  nand n65911(x65911, x65781, x65826);
  nand n65912(x65912, x65780, x65855);
  nand n65913(x65913, x65912, x65911);
  nand n65915(x65915, x65786, x65858);
  nand n65917(x65917, x65785, x65916);
  nand n65918(x65918, x65917, x65915);
  nand n65920(x65920, x65791, x65861);
  nand n65921(x65921, x65790, x65887);
  nand n65922(x65922, x65921, x65920);
  nand n65924(x65924, x65796, x65890);
  nand n65926(x65926, x65795, x65925);
  nand n65927(x65927, x65926, x65924);
  nand n65929(x65929, x65801, x65893);
  nand n65931(x65931, x65800, x65930);
  nand n65932(x65932, x65931, x65929);
  nand n65934(x65934, x65806, x65896);
  nand n65936(x65936, x65805, x65935);
  nand n65937(x65937, x65936, x65934);
  nand n65939(x65939, x65811, x65899);
  nand n65940(x65940, x65810, x65905);
  nand n65941(x65941, x65940, x65939);
  nand n65943(x65943, x65816, x65908);
  nand n65945(x65945, x65815, x65944);
  nand n65946(x65946, x65945, x65943);
  nand n65985(x65985, x65980, x65949);
  nand n65987(x65987, x65986, x65948);
  nand n65988(x65988, x65987, x65985);
  nand n65989(x65989, x65980, x65950);
  nand n65990(x65990, x65986, x65949);
  nand n65991(x65991, x65990, x65989);
  nand n65992(x65992, x65980, x65951);
  nand n65993(x65993, x65986, x65950);
  nand n65994(x65994, x65993, x65992);
  nand n65995(x65995, x65980, x65952);
  nand n65996(x65996, x65986, x65951);
  nand n65997(x65997, x65996, x65995);
  nand n65998(x65998, x65980, x65953);
  nand n65999(x65999, x65986, x65952);
  nand n66000(x66000, x65999, x65998);
  nand n66001(x66001, x65980, x65954);
  nand n66002(x66002, x65986, x65953);
  nand n66003(x66003, x66002, x66001);
  nand n66004(x66004, x65980, x65955);
  nand n66005(x66005, x65986, x65954);
  nand n66006(x66006, x66005, x66004);
  nand n66007(x66007, x65980, x65956);
  nand n66008(x66008, x65986, x65955);
  nand n66009(x66009, x66008, x66007);
  nand n66010(x66010, x65980, x65957);
  nand n66011(x66011, x65986, x65956);
  nand n66012(x66012, x66011, x66010);
  nand n66013(x66013, x65980, x65958);
  nand n66014(x66014, x65986, x65957);
  nand n66015(x66015, x66014, x66013);
  nand n66016(x66016, x65980, x65959);
  nand n66017(x66017, x65986, x65958);
  nand n66018(x66018, x66017, x66016);
  nand n66019(x66019, x65980, x65960);
  nand n66020(x66020, x65986, x65959);
  nand n66021(x66021, x66020, x66019);
  nand n66022(x66022, x65980, x65961);
  nand n66023(x66023, x65986, x65960);
  nand n66024(x66024, x66023, x66022);
  nand n66025(x66025, x65980, x65962);
  nand n66026(x66026, x65986, x65961);
  nand n66027(x66027, x66026, x66025);
  nand n66028(x66028, x65980, x65963);
  nand n66029(x66029, x65986, x65962);
  nand n66030(x66030, x66029, x66028);
  nand n66031(x66031, x65980, x65964);
  nand n66032(x66032, x65986, x65963);
  nand n66033(x66033, x66032, x66031);
  nand n66034(x66034, x65980, x65965);
  nand n66035(x66035, x65986, x65964);
  nand n66036(x66036, x66035, x66034);
  nand n66037(x66037, x65980, x65966);
  nand n66038(x66038, x65986, x65965);
  nand n66039(x66039, x66038, x66037);
  nand n66040(x66040, x65980, x65967);
  nand n66041(x66041, x65986, x65966);
  nand n66042(x66042, x66041, x66040);
  nand n66043(x66043, x65980, x65968);
  nand n66044(x66044, x65986, x65967);
  nand n66045(x66045, x66044, x66043);
  nand n66046(x66046, x65980, x65969);
  nand n66047(x66047, x65986, x65968);
  nand n66048(x66048, x66047, x66046);
  nand n66049(x66049, x65980, x65970);
  nand n66050(x66050, x65986, x65969);
  nand n66051(x66051, x66050, x66049);
  nand n66052(x66052, x65980, x65971);
  nand n66053(x66053, x65986, x65970);
  nand n66054(x66054, x66053, x66052);
  nand n66055(x66055, x65980, x65972);
  nand n66056(x66056, x65986, x65971);
  nand n66057(x66057, x66056, x66055);
  nand n66058(x66058, x65980, x65973);
  nand n66059(x66059, x65986, x65972);
  nand n66060(x66060, x66059, x66058);
  nand n66061(x66061, x65980, x65974);
  nand n66062(x66062, x65986, x65973);
  nand n66063(x66063, x66062, x66061);
  nand n66064(x66064, x65980, x65975);
  nand n66065(x66065, x65986, x65974);
  nand n66066(x66066, x66065, x66064);
  nand n66067(x66067, x65980, x65976);
  nand n66068(x66068, x65986, x65975);
  nand n66069(x66069, x66068, x66067);
  nand n66070(x66070, x65980, x65977);
  nand n66071(x66071, x65986, x65976);
  nand n66072(x66072, x66071, x66070);
  nand n66073(x66073, x65980, x65978);
  nand n66074(x66074, x65986, x65977);
  nand n66075(x66075, x66074, x66073);
  nand n66076(x66076, x65980, x65979);
  nand n66077(x66077, x65986, x65978);
  nand n66078(x66078, x66077, x66076);
  nand n66079(x66079, x65986, x65979);
  nand n66080(x66080, x65981, x65994);
  nand n66082(x66082, x66081, x65988);
  nand n66083(x66083, x66082, x66080);
  nand n66084(x66084, x65981, x65997);
  nand n66085(x66085, x66081, x65991);
  nand n66086(x66086, x66085, x66084);
  nand n66087(x66087, x65981, x66000);
  nand n66088(x66088, x66081, x65994);
  nand n66089(x66089, x66088, x66087);
  nand n66090(x66090, x65981, x66003);
  nand n66091(x66091, x66081, x65997);
  nand n66092(x66092, x66091, x66090);
  nand n66093(x66093, x65981, x66006);
  nand n66094(x66094, x66081, x66000);
  nand n66095(x66095, x66094, x66093);
  nand n66096(x66096, x65981, x66009);
  nand n66097(x66097, x66081, x66003);
  nand n66098(x66098, x66097, x66096);
  nand n66099(x66099, x65981, x66012);
  nand n66100(x66100, x66081, x66006);
  nand n66101(x66101, x66100, x66099);
  nand n66102(x66102, x65981, x66015);
  nand n66103(x66103, x66081, x66009);
  nand n66104(x66104, x66103, x66102);
  nand n66105(x66105, x65981, x66018);
  nand n66106(x66106, x66081, x66012);
  nand n66107(x66107, x66106, x66105);
  nand n66108(x66108, x65981, x66021);
  nand n66109(x66109, x66081, x66015);
  nand n66110(x66110, x66109, x66108);
  nand n66111(x66111, x65981, x66024);
  nand n66112(x66112, x66081, x66018);
  nand n66113(x66113, x66112, x66111);
  nand n66114(x66114, x65981, x66027);
  nand n66115(x66115, x66081, x66021);
  nand n66116(x66116, x66115, x66114);
  nand n66117(x66117, x65981, x66030);
  nand n66118(x66118, x66081, x66024);
  nand n66119(x66119, x66118, x66117);
  nand n66120(x66120, x65981, x66033);
  nand n66121(x66121, x66081, x66027);
  nand n66122(x66122, x66121, x66120);
  nand n66123(x66123, x65981, x66036);
  nand n66124(x66124, x66081, x66030);
  nand n66125(x66125, x66124, x66123);
  nand n66126(x66126, x65981, x66039);
  nand n66127(x66127, x66081, x66033);
  nand n66128(x66128, x66127, x66126);
  nand n66129(x66129, x65981, x66042);
  nand n66130(x66130, x66081, x66036);
  nand n66131(x66131, x66130, x66129);
  nand n66132(x66132, x65981, x66045);
  nand n66133(x66133, x66081, x66039);
  nand n66134(x66134, x66133, x66132);
  nand n66135(x66135, x65981, x66048);
  nand n66136(x66136, x66081, x66042);
  nand n66137(x66137, x66136, x66135);
  nand n66138(x66138, x65981, x66051);
  nand n66139(x66139, x66081, x66045);
  nand n66140(x66140, x66139, x66138);
  nand n66141(x66141, x65981, x66054);
  nand n66142(x66142, x66081, x66048);
  nand n66143(x66143, x66142, x66141);
  nand n66144(x66144, x65981, x66057);
  nand n66145(x66145, x66081, x66051);
  nand n66146(x66146, x66145, x66144);
  nand n66147(x66147, x65981, x66060);
  nand n66148(x66148, x66081, x66054);
  nand n66149(x66149, x66148, x66147);
  nand n66150(x66150, x65981, x66063);
  nand n66151(x66151, x66081, x66057);
  nand n66152(x66152, x66151, x66150);
  nand n66153(x66153, x65981, x66066);
  nand n66154(x66154, x66081, x66060);
  nand n66155(x66155, x66154, x66153);
  nand n66156(x66156, x65981, x66069);
  nand n66157(x66157, x66081, x66063);
  nand n66158(x66158, x66157, x66156);
  nand n66159(x66159, x65981, x66072);
  nand n66160(x66160, x66081, x66066);
  nand n66161(x66161, x66160, x66159);
  nand n66162(x66162, x65981, x66075);
  nand n66163(x66163, x66081, x66069);
  nand n66164(x66164, x66163, x66162);
  nand n66165(x66165, x65981, x66078);
  nand n66166(x66166, x66081, x66072);
  nand n66167(x66167, x66166, x66165);
  nand n66168(x66168, x65981, x86365);
  nand n66169(x66169, x66081, x66075);
  nand n66170(x66170, x66169, x66168);
  nand n66171(x66171, x66081, x66078);
  nand n66172(x66172, x66081, x86365);
  nand n66173(x66173, x65982, x66095);
  nand n66175(x66175, x66174, x66083);
  nand n66176(x66176, x66175, x66173);
  nand n66177(x66177, x65982, x66098);
  nand n66178(x66178, x66174, x66086);
  nand n66179(x66179, x66178, x66177);
  nand n66180(x66180, x65982, x66101);
  nand n66181(x66181, x66174, x66089);
  nand n66182(x66182, x66181, x66180);
  nand n66183(x66183, x65982, x66104);
  nand n66184(x66184, x66174, x66092);
  nand n66185(x66185, x66184, x66183);
  nand n66186(x66186, x65982, x66107);
  nand n66187(x66187, x66174, x66095);
  nand n66188(x66188, x66187, x66186);
  nand n66189(x66189, x65982, x66110);
  nand n66190(x66190, x66174, x66098);
  nand n66191(x66191, x66190, x66189);
  nand n66192(x66192, x65982, x66113);
  nand n66193(x66193, x66174, x66101);
  nand n66194(x66194, x66193, x66192);
  nand n66195(x66195, x65982, x66116);
  nand n66196(x66196, x66174, x66104);
  nand n66197(x66197, x66196, x66195);
  nand n66198(x66198, x65982, x66119);
  nand n66199(x66199, x66174, x66107);
  nand n66200(x66200, x66199, x66198);
  nand n66201(x66201, x65982, x66122);
  nand n66202(x66202, x66174, x66110);
  nand n66203(x66203, x66202, x66201);
  nand n66204(x66204, x65982, x66125);
  nand n66205(x66205, x66174, x66113);
  nand n66206(x66206, x66205, x66204);
  nand n66207(x66207, x65982, x66128);
  nand n66208(x66208, x66174, x66116);
  nand n66209(x66209, x66208, x66207);
  nand n66210(x66210, x65982, x66131);
  nand n66211(x66211, x66174, x66119);
  nand n66212(x66212, x66211, x66210);
  nand n66213(x66213, x65982, x66134);
  nand n66214(x66214, x66174, x66122);
  nand n66215(x66215, x66214, x66213);
  nand n66216(x66216, x65982, x66137);
  nand n66217(x66217, x66174, x66125);
  nand n66218(x66218, x66217, x66216);
  nand n66219(x66219, x65982, x66140);
  nand n66220(x66220, x66174, x66128);
  nand n66221(x66221, x66220, x66219);
  nand n66222(x66222, x65982, x66143);
  nand n66223(x66223, x66174, x66131);
  nand n66224(x66224, x66223, x66222);
  nand n66225(x66225, x65982, x66146);
  nand n66226(x66226, x66174, x66134);
  nand n66227(x66227, x66226, x66225);
  nand n66228(x66228, x65982, x66149);
  nand n66229(x66229, x66174, x66137);
  nand n66230(x66230, x66229, x66228);
  nand n66231(x66231, x65982, x66152);
  nand n66232(x66232, x66174, x66140);
  nand n66233(x66233, x66232, x66231);
  nand n66234(x66234, x65982, x66155);
  nand n66235(x66235, x66174, x66143);
  nand n66236(x66236, x66235, x66234);
  nand n66237(x66237, x65982, x66158);
  nand n66238(x66238, x66174, x66146);
  nand n66239(x66239, x66238, x66237);
  nand n66240(x66240, x65982, x66161);
  nand n66241(x66241, x66174, x66149);
  nand n66242(x66242, x66241, x66240);
  nand n66243(x66243, x65982, x66164);
  nand n66244(x66244, x66174, x66152);
  nand n66245(x66245, x66244, x66243);
  nand n66246(x66246, x65982, x66167);
  nand n66247(x66247, x66174, x66155);
  nand n66248(x66248, x66247, x66246);
  nand n66249(x66249, x65982, x66170);
  nand n66250(x66250, x66174, x66158);
  nand n66251(x66251, x66250, x66249);
  nand n66252(x66252, x65982, x86366);
  nand n66253(x66253, x66174, x66161);
  nand n66254(x66254, x66253, x66252);
  nand n66255(x66255, x65982, x86367);
  nand n66256(x66256, x66174, x66164);
  nand n66257(x66257, x66256, x66255);
  nand n66258(x66258, x66174, x66167);
  nand n66259(x66259, x66174, x66170);
  nand n66260(x66260, x66174, x86366);
  nand n66261(x66261, x66174, x86367);
  nand n66262(x66262, x65983, x66200);
  nand n66264(x66264, x66263, x66176);
  nand n66265(x66265, x66264, x66262);
  nand n66266(x66266, x65983, x66203);
  nand n66267(x66267, x66263, x66179);
  nand n66268(x66268, x66267, x66266);
  nand n66269(x66269, x65983, x66206);
  nand n66270(x66270, x66263, x66182);
  nand n66271(x66271, x66270, x66269);
  nand n66272(x66272, x65983, x66209);
  nand n66273(x66273, x66263, x66185);
  nand n66274(x66274, x66273, x66272);
  nand n66275(x66275, x65983, x66212);
  nand n66276(x66276, x66263, x66188);
  nand n66277(x66277, x66276, x66275);
  nand n66278(x66278, x65983, x66215);
  nand n66279(x66279, x66263, x66191);
  nand n66280(x66280, x66279, x66278);
  nand n66281(x66281, x65983, x66218);
  nand n66282(x66282, x66263, x66194);
  nand n66283(x66283, x66282, x66281);
  nand n66284(x66284, x65983, x66221);
  nand n66285(x66285, x66263, x66197);
  nand n66286(x66286, x66285, x66284);
  nand n66287(x66287, x65983, x66224);
  nand n66288(x66288, x66263, x66200);
  nand n66289(x66289, x66288, x66287);
  nand n66290(x66290, x65983, x66227);
  nand n66291(x66291, x66263, x66203);
  nand n66292(x66292, x66291, x66290);
  nand n66293(x66293, x65983, x66230);
  nand n66294(x66294, x66263, x66206);
  nand n66295(x66295, x66294, x66293);
  nand n66296(x66296, x65983, x66233);
  nand n66297(x66297, x66263, x66209);
  nand n66298(x66298, x66297, x66296);
  nand n66299(x66299, x65983, x66236);
  nand n66300(x66300, x66263, x66212);
  nand n66301(x66301, x66300, x66299);
  nand n66302(x66302, x65983, x66239);
  nand n66303(x66303, x66263, x66215);
  nand n66304(x66304, x66303, x66302);
  nand n66305(x66305, x65983, x66242);
  nand n66306(x66306, x66263, x66218);
  nand n66307(x66307, x66306, x66305);
  nand n66308(x66308, x65983, x66245);
  nand n66309(x66309, x66263, x66221);
  nand n66310(x66310, x66309, x66308);
  nand n66311(x66311, x65983, x66248);
  nand n66312(x66312, x66263, x66224);
  nand n66313(x66313, x66312, x66311);
  nand n66314(x66314, x65983, x66251);
  nand n66315(x66315, x66263, x66227);
  nand n66316(x66316, x66315, x66314);
  nand n66317(x66317, x65983, x66254);
  nand n66318(x66318, x66263, x66230);
  nand n66319(x66319, x66318, x66317);
  nand n66320(x66320, x65983, x66257);
  nand n66321(x66321, x66263, x66233);
  nand n66322(x66322, x66321, x66320);
  nand n66323(x66323, x65983, x86368);
  nand n66324(x66324, x66263, x66236);
  nand n66325(x66325, x66324, x66323);
  nand n66326(x66326, x65983, x86369);
  nand n66327(x66327, x66263, x66239);
  nand n66328(x66328, x66327, x66326);
  nand n66329(x66329, x65983, x86370);
  nand n66330(x66330, x66263, x66242);
  nand n66331(x66331, x66330, x66329);
  nand n66332(x66332, x65983, x86371);
  nand n66333(x66333, x66263, x66245);
  nand n66334(x66334, x66333, x66332);
  nand n66335(x66335, x66263, x66248);
  nand n66336(x66336, x66263, x66251);
  nand n66337(x66337, x66263, x66254);
  nand n66338(x66338, x66263, x66257);
  nand n66339(x66339, x66263, x86368);
  nand n66340(x66340, x66263, x86369);
  nand n66341(x66341, x66263, x86370);
  nand n66342(x66342, x66263, x86371);
  nand n66343(x66343, x65984, x66313);
  nand n66345(x66345, x66344, x66265);
  nand n66346(x66346, x66345, x66343);
  nand n66347(x66347, x65984, x66316);
  nand n66348(x66348, x66344, x66268);
  nand n66349(x66349, x66348, x66347);
  nand n66350(x66350, x65984, x66319);
  nand n66351(x66351, x66344, x66271);
  nand n66352(x66352, x66351, x66350);
  nand n66353(x66353, x65984, x66322);
  nand n66354(x66354, x66344, x66274);
  nand n66355(x66355, x66354, x66353);
  nand n66356(x66356, x65984, x66325);
  nand n66357(x66357, x66344, x66277);
  nand n66358(x66358, x66357, x66356);
  nand n66359(x66359, x65984, x66328);
  nand n66360(x66360, x66344, x66280);
  nand n66361(x66361, x66360, x66359);
  nand n66362(x66362, x65984, x66331);
  nand n66363(x66363, x66344, x66283);
  nand n66364(x66364, x66363, x66362);
  nand n66365(x66365, x65984, x66334);
  nand n66366(x66366, x66344, x66286);
  nand n66367(x66367, x66366, x66365);
  nand n66368(x66368, x65984, x86372);
  nand n66369(x66369, x66344, x66289);
  nand n66370(x66370, x66369, x66368);
  nand n66371(x66371, x65984, x86373);
  nand n66372(x66372, x66344, x66292);
  nand n66373(x66373, x66372, x66371);
  nand n66374(x66374, x65984, x86374);
  nand n66375(x66375, x66344, x66295);
  nand n66376(x66376, x66375, x66374);
  nand n66377(x66377, x65984, x86375);
  nand n66378(x66378, x66344, x66298);
  nand n66379(x66379, x66378, x66377);
  nand n66380(x66380, x65984, x86376);
  nand n66381(x66381, x66344, x66301);
  nand n66382(x66382, x66381, x66380);
  nand n66383(x66383, x65984, x86377);
  nand n66384(x66384, x66344, x66304);
  nand n66385(x66385, x66384, x66383);
  nand n66386(x66386, x65984, x86378);
  nand n66387(x66387, x66344, x66307);
  nand n66388(x66388, x66387, x66386);
  nand n66389(x66389, x65984, x86379);
  nand n66390(x66390, x66344, x66310);
  nand n66391(x66391, x66390, x66389);
  nand n66392(x66392, x66344, x66313);
  nand n66393(x66393, x66344, x66316);
  nand n66394(x66394, x66344, x66319);
  nand n66395(x66395, x66344, x66322);
  nand n66396(x66396, x66344, x66325);
  nand n66397(x66397, x66344, x66328);
  nand n66398(x66398, x66344, x66331);
  nand n66399(x66399, x66344, x66334);
  nand n66400(x66400, x66344, x86372);
  nand n66401(x66401, x66344, x86373);
  nand n66402(x66402, x66344, x86374);
  nand n66403(x66403, x66344, x86375);
  nand n66404(x66404, x66344, x86376);
  nand n66405(x66405, x66344, x86377);
  nand n66406(x66406, x66344, x86378);
  nand n66407(x66407, x66344, x86379);
  nand n66408(x66408, x83367, x76792);
  nand n66410(x66410, x62931, x66409);
  nand n66411(x66411, x68741, x66413);
  nand n66412(x66412, x66411, x66410);
  nand n66414(x66414, x62931, x76774);
  nand n66415(x66415, x68741, x66417);
  nand n66416(x66416, x66415, x66414);
  nand n66418(x66418, x62931, x76777);
  nand n66419(x66419, x68741, x66421);
  nand n66420(x66420, x66419, x66418);
  nand n66422(x66422, x62931, x76780);
  nand n66423(x66423, x68741, x66425);
  nand n66424(x66424, x66423, x66422);
  nand n66426(x66426, x62931, x76783);
  nand n66427(x66427, x68741, x66429);
  nand n66428(x66428, x66427, x66426);
  nand n66430(x66430, x62931, x76786);
  nand n66431(x66431, x68741, x66433);
  nand n66432(x66432, x66431, x66430);
  nand n66434(x66434, x62931, x76789);
  nand n66435(x66435, x68741, x66437);
  nand n66436(x66436, x66435, x66434);
  nand n66438(x66438, x62931, x76810);
  nand n66439(x66439, x68741, x66441);
  nand n66440(x66440, x66439, x66438);
  nand n66442(x66442, x62931, x76813);
  nand n66443(x66443, x68741, x66445);
  nand n66444(x66444, x66443, x66442);
  nand n66446(x66446, x62931, x76816);
  nand n66447(x66447, x68741, x66449);
  nand n66448(x66448, x66447, x66446);
  nand n66450(x66450, x62931, x76819);
  nand n66451(x66451, x68741, x66453);
  nand n66452(x66452, x66451, x66450);
  nand n66454(x66454, x62931, x76822);
  nand n66455(x66455, x68741, x66457);
  nand n66456(x66456, x66455, x66454);
  nand n66458(x66458, x62931, x76825);
  nand n66459(x66459, x68741, x66461);
  nand n66460(x66460, x66459, x66458);
  nand n66462(x66462, x62931, x76828);
  nand n66463(x66463, x68741, x66465);
  nand n66464(x66464, x66463, x66462);
  nand n66466(x66466, x62931, x76831);
  nand n66467(x66467, x68741, x66469);
  nand n66468(x66468, x66467, x66466);
  nand n66471(x66471, x66601, x66470);
  nand n66602(x66602, x78106, x78010);
  nand n66604(x66604, x66603, x78265);
  nand n66605(x66605, x66604, x66602);
  nand n66606(x66606, x78106, x78013);
  nand n66607(x66607, x66603, x78268);
  nand n66608(x66608, x66607, x66606);
  nand n66609(x66609, x78106, x78016);
  nand n66610(x66610, x66603, x78271);
  nand n66611(x66611, x66610, x66609);
  nand n66612(x66612, x78106, x78019);
  nand n66613(x66613, x66603, x78274);
  nand n66614(x66614, x66613, x66612);
  nand n66615(x66615, x78106, x78022);
  nand n66616(x66616, x66603, x78277);
  nand n66617(x66617, x66616, x66615);
  nand n66618(x66618, x78106, x78025);
  nand n66619(x66619, x66603, x78280);
  nand n66620(x66620, x66619, x66618);
  nand n66621(x66621, x78106, x78028);
  nand n66622(x66622, x66603, x78283);
  nand n66623(x66623, x66622, x66621);
  nand n66624(x66624, x78106, x78031);
  nand n66625(x66625, x66603, x78286);
  nand n66626(x66626, x66625, x66624);
  nand n66627(x66627, x78106, x78034);
  nand n66628(x66628, x66603, x78289);
  nand n66629(x66629, x66628, x66627);
  nand n66630(x66630, x78106, x78037);
  nand n66631(x66631, x66603, x78292);
  nand n66632(x66632, x66631, x66630);
  nand n66633(x66633, x78106, x78040);
  nand n66634(x66634, x66603, x78295);
  nand n66635(x66635, x66634, x66633);
  nand n66636(x66636, x78106, x78043);
  nand n66637(x66637, x66603, x78298);
  nand n66638(x66638, x66637, x66636);
  nand n66639(x66639, x78106, x78046);
  nand n66640(x66640, x66603, x78301);
  nand n66641(x66641, x66640, x66639);
  nand n66642(x66642, x78106, x78049);
  nand n66643(x66643, x66603, x78304);
  nand n66644(x66644, x66643, x66642);
  nand n66645(x66645, x78106, x78052);
  nand n66646(x66646, x66603, x78307);
  nand n66647(x66647, x66646, x66645);
  nand n66648(x66648, x78106, x78055);
  nand n66649(x66649, x66603, x78310);
  nand n66650(x66650, x66649, x66648);
  nand n66651(x66651, x78106, x78058);
  nand n66652(x66652, x66603, x78313);
  nand n66653(x66653, x66652, x66651);
  nand n66654(x66654, x78106, x78061);
  nand n66655(x66655, x66603, x78316);
  nand n66656(x66656, x66655, x66654);
  nand n66657(x66657, x78106, x78064);
  nand n66658(x66658, x66603, x78319);
  nand n66659(x66659, x66658, x66657);
  nand n66660(x66660, x78106, x78067);
  nand n66661(x66661, x66603, x78322);
  nand n66662(x66662, x66661, x66660);
  nand n66663(x66663, x78106, x78070);
  nand n66664(x66664, x66603, x78325);
  nand n66665(x66665, x66664, x66663);
  nand n66666(x66666, x78106, x78073);
  nand n66667(x66667, x66603, x78328);
  nand n66668(x66668, x66667, x66666);
  nand n66669(x66669, x78106, x78076);
  nand n66670(x66670, x66603, x78331);
  nand n66671(x66671, x66670, x66669);
  nand n66672(x66672, x78106, x78079);
  nand n66673(x66673, x66603, x78334);
  nand n66674(x66674, x66673, x66672);
  nand n66675(x66675, x78106, x78082);
  nand n66676(x66676, x66603, x78337);
  nand n66677(x66677, x66676, x66675);
  nand n66678(x66678, x78106, x78085);
  nand n66679(x66679, x66603, x78340);
  nand n66680(x66680, x66679, x66678);
  nand n66681(x66681, x78106, x78088);
  nand n66682(x66682, x66603, x78343);
  nand n66683(x66683, x66682, x66681);
  nand n66684(x66684, x78106, x78091);
  nand n66685(x66685, x66603, x78346);
  nand n66686(x66686, x66685, x66684);
  nand n66687(x66687, x78106, x78094);
  nand n66688(x66688, x66603, x78349);
  nand n66689(x66689, x66688, x66687);
  nand n66690(x66690, x78106, x78097);
  nand n66691(x66691, x66603, x78352);
  nand n66692(x66692, x66691, x66690);
  nand n66693(x66693, x78106, x78100);
  nand n66694(x66694, x66603, x78355);
  nand n66695(x66695, x66694, x66693);
  nand n66696(x66696, x78106, x78103);
  nand n66697(x66697, x66603, x78358);
  nand n66698(x66698, x66697, x66696);
  nand n66699(x66699, x66603, x78559);
  nand n66700(x66700, x66699, x66602);
  nand n66701(x66701, x66603, x78562);
  nand n66702(x66702, x66701, x66606);
  nand n66703(x66703, x66603, x78565);
  nand n66704(x66704, x66703, x66609);
  nand n66705(x66705, x66603, x78568);
  nand n66706(x66706, x66705, x66612);
  nand n66707(x66707, x66603, x78571);
  nand n66708(x66708, x66707, x66615);
  nand n66709(x66709, x66603, x78574);
  nand n66710(x66710, x66709, x66618);
  nand n66711(x66711, x66603, x78577);
  nand n66712(x66712, x66711, x66621);
  nand n66713(x66713, x66603, x78580);
  nand n66714(x66714, x66713, x66624);
  nand n66715(x66715, x66603, x78583);
  nand n66716(x66716, x66715, x66627);
  nand n66717(x66717, x66603, x78586);
  nand n66718(x66718, x66717, x66630);
  nand n66719(x66719, x66603, x78589);
  nand n66720(x66720, x66719, x66633);
  nand n66721(x66721, x66603, x78592);
  nand n66722(x66722, x66721, x66636);
  nand n66723(x66723, x66603, x78595);
  nand n66724(x66724, x66723, x66639);
  nand n66725(x66725, x66603, x78598);
  nand n66726(x66726, x66725, x66642);
  nand n66727(x66727, x66603, x78601);
  nand n66728(x66728, x66727, x66645);
  nand n66729(x66729, x66603, x78604);
  nand n66730(x66730, x66729, x66648);
  nand n66731(x66731, x66603, x78607);
  nand n66732(x66732, x66731, x66651);
  nand n66733(x66733, x66603, x78610);
  nand n66734(x66734, x66733, x66654);
  nand n66735(x66735, x66603, x78613);
  nand n66736(x66736, x66735, x66657);
  nand n66737(x66737, x66603, x78616);
  nand n66738(x66738, x66737, x66660);
  nand n66739(x66739, x66603, x78619);
  nand n66740(x66740, x66739, x66663);
  nand n66741(x66741, x66603, x78622);
  nand n66742(x66742, x66741, x66666);
  nand n66743(x66743, x66603, x78625);
  nand n66744(x66744, x66743, x66669);
  nand n66745(x66745, x66603, x78628);
  nand n66746(x66746, x66745, x66672);
  nand n66747(x66747, x66603, x78631);
  nand n66748(x66748, x66747, x66675);
  nand n66749(x66749, x66603, x78634);
  nand n66750(x66750, x66749, x66678);
  nand n66751(x66751, x66603, x78637);
  nand n66752(x66752, x66751, x66681);
  nand n66753(x66753, x66603, x78640);
  nand n66754(x66754, x66753, x66684);
  nand n66755(x66755, x66603, x78643);
  nand n66756(x66756, x66755, x66687);
  nand n66757(x66757, x66603, x78646);
  nand n66758(x66758, x66757, x66690);
  nand n66759(x66759, x66603, x78649);
  nand n66760(x66760, x66759, x66693);
  nand n66761(x66761, x66603, x78652);
  nand n66762(x66762, x66761, x66696);
  nand n66763(x66763, x66603, x78853);
  nand n66764(x66764, x66763, x66602);
  nand n66765(x66765, x66603, x78856);
  nand n66766(x66766, x66765, x66606);
  nand n66767(x66767, x66603, x78859);
  nand n66768(x66768, x66767, x66609);
  nand n66769(x66769, x66603, x78862);
  nand n66770(x66770, x66769, x66612);
  nand n66771(x66771, x66603, x78865);
  nand n66772(x66772, x66771, x66615);
  nand n66773(x66773, x66603, x78868);
  nand n66774(x66774, x66773, x66618);
  nand n66775(x66775, x66603, x78871);
  nand n66776(x66776, x66775, x66621);
  nand n66777(x66777, x66603, x78874);
  nand n66778(x66778, x66777, x66624);
  nand n66779(x66779, x66603, x78877);
  nand n66780(x66780, x66779, x66627);
  nand n66781(x66781, x66603, x78880);
  nand n66782(x66782, x66781, x66630);
  nand n66783(x66783, x66603, x78883);
  nand n66784(x66784, x66783, x66633);
  nand n66785(x66785, x66603, x78886);
  nand n66786(x66786, x66785, x66636);
  nand n66787(x66787, x66603, x78889);
  nand n66788(x66788, x66787, x66639);
  nand n66789(x66789, x66603, x78892);
  nand n66790(x66790, x66789, x66642);
  nand n66791(x66791, x66603, x78895);
  nand n66792(x66792, x66791, x66645);
  nand n66793(x66793, x66603, x78898);
  nand n66794(x66794, x66793, x66648);
  nand n66795(x66795, x66603, x78901);
  nand n66796(x66796, x66795, x66651);
  nand n66797(x66797, x66603, x78904);
  nand n66798(x66798, x66797, x66654);
  nand n66799(x66799, x66603, x78907);
  nand n66800(x66800, x66799, x66657);
  nand n66801(x66801, x66603, x78910);
  nand n66802(x66802, x66801, x66660);
  nand n66803(x66803, x66603, x78913);
  nand n66804(x66804, x66803, x66663);
  nand n66805(x66805, x66603, x78916);
  nand n66806(x66806, x66805, x66666);
  nand n66807(x66807, x66603, x78919);
  nand n66808(x66808, x66807, x66669);
  nand n66809(x66809, x66603, x78922);
  nand n66810(x66810, x66809, x66672);
  nand n66811(x66811, x66603, x78925);
  nand n66812(x66812, x66811, x66675);
  nand n66813(x66813, x66603, x78928);
  nand n66814(x66814, x66813, x66678);
  nand n66815(x66815, x66603, x78931);
  nand n66816(x66816, x66815, x66681);
  nand n66817(x66817, x66603, x78934);
  nand n66818(x66818, x66817, x66684);
  nand n66819(x66819, x66603, x78937);
  nand n66820(x66820, x66819, x66687);
  nand n66821(x66821, x66603, x78940);
  nand n66822(x66822, x66821, x66690);
  nand n66823(x66823, x66603, x78943);
  nand n66824(x66824, x66823, x66693);
  nand n66825(x66825, x66603, x78946);
  nand n66826(x66826, x66825, x66696);
  nand n66827(x66827, x66603, x79147);
  nand n66828(x66828, x66827, x66602);
  nand n66829(x66829, x66603, x79150);
  nand n66830(x66830, x66829, x66606);
  nand n66831(x66831, x66603, x79153);
  nand n66832(x66832, x66831, x66609);
  nand n66833(x66833, x66603, x79156);
  nand n66834(x66834, x66833, x66612);
  nand n66835(x66835, x66603, x79159);
  nand n66836(x66836, x66835, x66615);
  nand n66837(x66837, x66603, x79162);
  nand n66838(x66838, x66837, x66618);
  nand n66839(x66839, x66603, x79165);
  nand n66840(x66840, x66839, x66621);
  nand n66841(x66841, x66603, x79168);
  nand n66842(x66842, x66841, x66624);
  nand n66843(x66843, x66603, x79171);
  nand n66844(x66844, x66843, x66627);
  nand n66845(x66845, x66603, x79174);
  nand n66846(x66846, x66845, x66630);
  nand n66847(x66847, x66603, x79177);
  nand n66848(x66848, x66847, x66633);
  nand n66849(x66849, x66603, x79180);
  nand n66850(x66850, x66849, x66636);
  nand n66851(x66851, x66603, x79183);
  nand n66852(x66852, x66851, x66639);
  nand n66853(x66853, x66603, x79186);
  nand n66854(x66854, x66853, x66642);
  nand n66855(x66855, x66603, x79189);
  nand n66856(x66856, x66855, x66645);
  nand n66857(x66857, x66603, x79192);
  nand n66858(x66858, x66857, x66648);
  nand n66859(x66859, x66603, x79195);
  nand n66860(x66860, x66859, x66651);
  nand n66861(x66861, x66603, x79198);
  nand n66862(x66862, x66861, x66654);
  nand n66863(x66863, x66603, x79201);
  nand n66864(x66864, x66863, x66657);
  nand n66865(x66865, x66603, x79204);
  nand n66866(x66866, x66865, x66660);
  nand n66867(x66867, x66603, x79207);
  nand n66868(x66868, x66867, x66663);
  nand n66869(x66869, x66603, x79210);
  nand n66870(x66870, x66869, x66666);
  nand n66871(x66871, x66603, x79213);
  nand n66872(x66872, x66871, x66669);
  nand n66873(x66873, x66603, x79216);
  nand n66874(x66874, x66873, x66672);
  nand n66875(x66875, x66603, x79219);
  nand n66876(x66876, x66875, x66675);
  nand n66877(x66877, x66603, x79222);
  nand n66878(x66878, x66877, x66678);
  nand n66879(x66879, x66603, x79225);
  nand n66880(x66880, x66879, x66681);
  nand n66881(x66881, x66603, x79228);
  nand n66882(x66882, x66881, x66684);
  nand n66883(x66883, x66603, x79231);
  nand n66884(x66884, x66883, x66687);
  nand n66885(x66885, x66603, x79234);
  nand n66886(x66886, x66885, x66690);
  nand n66887(x66887, x66603, x79237);
  nand n66888(x66888, x66887, x66693);
  nand n66889(x66889, x66603, x79240);
  nand n66890(x66890, x66889, x66696);
  nand n66891(x66891, x66472, x66473);
  nand n66892(x66892, x66471, x66894);
  nand n66893(x66893, x66892, x66891);
  nand n66895(x66895, x66472, x66474);
  nand n66896(x66896, x66471, x66898);
  nand n66897(x66897, x66896, x66895);
  nand n66899(x66899, x66472, x66475);
  nand n66900(x66900, x66471, x66902);
  nand n66901(x66901, x66900, x66899);
  nand n66903(x66903, x66472, x66476);
  nand n66904(x66904, x66471, x66906);
  nand n66905(x66905, x66904, x66903);
  nand n66907(x66907, x66472, x66477);
  nand n66908(x66908, x66471, x66910);
  nand n66909(x66909, x66908, x66907);
  nand n66911(x66911, x66472, x66478);
  nand n66912(x66912, x66471, x66914);
  nand n66913(x66913, x66912, x66911);
  nand n66915(x66915, x66472, x66479);
  nand n66916(x66916, x66471, x66918);
  nand n66917(x66917, x66916, x66915);
  nand n66919(x66919, x66472, x66480);
  nand n66920(x66920, x66471, x66922);
  nand n66921(x66921, x66920, x66919);
  nand n66923(x66923, x66472, x66481);
  nand n66924(x66924, x66471, x66926);
  nand n66925(x66925, x66924, x66923);
  nand n66927(x66927, x66472, x66482);
  nand n66928(x66928, x66471, x66930);
  nand n66929(x66929, x66928, x66927);
  nand n66931(x66931, x66472, x66483);
  nand n66932(x66932, x66471, x66934);
  nand n66933(x66933, x66932, x66931);
  nand n66935(x66935, x66472, x66484);
  nand n66936(x66936, x66471, x66938);
  nand n66937(x66937, x66936, x66935);
  nand n66939(x66939, x66472, x66485);
  nand n66940(x66940, x66471, x66942);
  nand n66941(x66941, x66940, x66939);
  nand n66943(x66943, x66472, x66486);
  nand n66944(x66944, x66471, x66946);
  nand n66945(x66945, x66944, x66943);
  nand n66947(x66947, x66472, x66487);
  nand n66948(x66948, x66471, x66950);
  nand n66949(x66949, x66948, x66947);
  nand n66951(x66951, x66472, x66488);
  nand n66952(x66952, x66471, x66954);
  nand n66953(x66953, x66952, x66951);
  nand n66955(x66955, x66472, x66489);
  nand n66956(x66956, x66471, x66958);
  nand n66957(x66957, x66956, x66955);
  nand n66959(x66959, x66472, x66490);
  nand n66960(x66960, x66471, x66962);
  nand n66961(x66961, x66960, x66959);
  nand n66963(x66963, x66472, x66491);
  nand n66964(x66964, x66471, x66966);
  nand n66965(x66965, x66964, x66963);
  nand n66967(x66967, x66472, x66492);
  nand n66968(x66968, x66471, x66970);
  nand n66969(x66969, x66968, x66967);
  nand n66971(x66971, x66472, x66493);
  nand n66972(x66972, x66471, x66974);
  nand n66973(x66973, x66972, x66971);
  nand n66975(x66975, x66472, x66494);
  nand n66976(x66976, x66471, x66978);
  nand n66977(x66977, x66976, x66975);
  nand n66979(x66979, x66472, x66495);
  nand n66980(x66980, x66471, x66982);
  nand n66981(x66981, x66980, x66979);
  nand n66983(x66983, x66472, x66496);
  nand n66984(x66984, x66471, x66986);
  nand n66985(x66985, x66984, x66983);
  nand n66987(x66987, x66472, x66497);
  nand n66988(x66988, x66471, x66990);
  nand n66989(x66989, x66988, x66987);
  nand n66991(x66991, x66472, x66498);
  nand n66992(x66992, x66471, x66994);
  nand n66993(x66993, x66992, x66991);
  nand n66995(x66995, x66472, x66499);
  nand n66996(x66996, x66471, x66998);
  nand n66997(x66997, x66996, x66995);
  nand n66999(x66999, x66472, x66500);
  nand n67000(x67000, x66471, x67002);
  nand n67001(x67001, x67000, x66999);
  nand n67003(x67003, x66472, x66501);
  nand n67004(x67004, x66471, x67006);
  nand n67005(x67005, x67004, x67003);
  nand n67007(x67007, x66472, x66502);
  nand n67008(x67008, x66471, x67010);
  nand n67009(x67009, x67008, x67007);
  nand n67011(x67011, x66472, x66503);
  nand n67012(x67012, x66471, x67014);
  nand n67013(x67013, x67012, x67011);
  nand n67015(x67015, x66472, x66504);
  nand n67016(x67016, x66471, x67018);
  nand n67017(x67017, x67016, x67015);
  nand n67019(x67019, x66472, x66505);
  nand n67020(x67020, x66471, x67022);
  nand n67021(x67021, x67020, x67019);
  nand n67023(x67023, x66472, x66506);
  nand n67024(x67024, x66471, x67026);
  nand n67025(x67025, x67024, x67023);
  nand n67027(x67027, x66472, x66507);
  nand n67028(x67028, x66471, x67030);
  nand n67029(x67029, x67028, x67027);
  nand n67031(x67031, x66472, x66508);
  nand n67032(x67032, x66471, x67034);
  nand n67033(x67033, x67032, x67031);
  nand n67035(x67035, x66472, x66509);
  nand n67036(x67036, x66471, x67038);
  nand n67037(x67037, x67036, x67035);
  nand n67039(x67039, x66472, x66510);
  nand n67040(x67040, x66471, x67042);
  nand n67041(x67041, x67040, x67039);
  nand n67043(x67043, x66472, x66511);
  nand n67044(x67044, x66471, x67046);
  nand n67045(x67045, x67044, x67043);
  nand n67047(x67047, x66472, x66512);
  nand n67048(x67048, x66471, x67050);
  nand n67049(x67049, x67048, x67047);
  nand n67051(x67051, x66472, x66513);
  nand n67052(x67052, x66471, x67054);
  nand n67053(x67053, x67052, x67051);
  nand n67055(x67055, x66472, x66514);
  nand n67056(x67056, x66471, x67058);
  nand n67057(x67057, x67056, x67055);
  nand n67059(x67059, x66472, x66515);
  nand n67060(x67060, x66471, x67062);
  nand n67061(x67061, x67060, x67059);
  nand n67063(x67063, x66472, x66516);
  nand n67064(x67064, x66471, x67066);
  nand n67065(x67065, x67064, x67063);
  nand n67067(x67067, x66472, x66517);
  nand n67068(x67068, x66471, x67070);
  nand n67069(x67069, x67068, x67067);
  nand n67071(x67071, x66472, x66518);
  nand n67072(x67072, x66471, x67074);
  nand n67073(x67073, x67072, x67071);
  nand n67075(x67075, x66472, x66519);
  nand n67076(x67076, x66471, x67078);
  nand n67077(x67077, x67076, x67075);
  nand n67079(x67079, x66472, x66520);
  nand n67080(x67080, x66471, x67082);
  nand n67081(x67081, x67080, x67079);
  nand n67083(x67083, x66472, x66521);
  nand n67084(x67084, x66471, x67086);
  nand n67085(x67085, x67084, x67083);
  nand n67087(x67087, x66472, x66522);
  nand n67088(x67088, x66471, x67090);
  nand n67089(x67089, x67088, x67087);
  nand n67091(x67091, x66472, x66523);
  nand n67092(x67092, x66471, x67094);
  nand n67093(x67093, x67092, x67091);
  nand n67095(x67095, x66472, x66524);
  nand n67096(x67096, x66471, x67098);
  nand n67097(x67097, x67096, x67095);
  nand n67099(x67099, x66472, x66525);
  nand n67100(x67100, x66471, x67102);
  nand n67101(x67101, x67100, x67099);
  nand n67103(x67103, x66472, x66526);
  nand n67104(x67104, x66471, x67106);
  nand n67105(x67105, x67104, x67103);
  nand n67107(x67107, x66472, x66527);
  nand n67108(x67108, x66471, x67110);
  nand n67109(x67109, x67108, x67107);
  nand n67111(x67111, x66472, x66528);
  nand n67112(x67112, x66471, x67114);
  nand n67113(x67113, x67112, x67111);
  nand n67115(x67115, x66472, x66529);
  nand n67116(x67116, x66471, x67118);
  nand n67117(x67117, x67116, x67115);
  nand n67119(x67119, x66472, x66530);
  nand n67120(x67120, x66471, x67122);
  nand n67121(x67121, x67120, x67119);
  nand n67123(x67123, x66472, x66531);
  nand n67124(x67124, x66471, x67126);
  nand n67125(x67125, x67124, x67123);
  nand n67127(x67127, x66472, x66532);
  nand n67128(x67128, x66471, x67130);
  nand n67129(x67129, x67128, x67127);
  nand n67131(x67131, x66472, x66533);
  nand n67132(x67132, x66471, x67134);
  nand n67133(x67133, x67132, x67131);
  nand n67135(x67135, x66472, x66534);
  nand n67136(x67136, x66471, x67138);
  nand n67137(x67137, x67136, x67135);
  nand n67139(x67139, x66472, x66535);
  nand n67140(x67140, x66471, x67142);
  nand n67141(x67141, x67140, x67139);
  nand n67143(x67143, x66472, x66536);
  nand n67144(x67144, x66471, x67146);
  nand n67145(x67145, x67144, x67143);
  nand n67147(x67147, x66472, x66537);
  nand n67148(x67148, x66471, x67150);
  nand n67149(x67149, x67148, x67147);
  nand n67151(x67151, x66472, x66538);
  nand n67152(x67152, x66471, x67154);
  nand n67153(x67153, x67152, x67151);
  nand n67155(x67155, x66472, x66539);
  nand n67156(x67156, x66471, x67158);
  nand n67157(x67157, x67156, x67155);
  nand n67159(x67159, x66472, x66540);
  nand n67160(x67160, x66471, x67162);
  nand n67161(x67161, x67160, x67159);
  nand n67163(x67163, x66472, x66541);
  nand n67164(x67164, x66471, x67166);
  nand n67165(x67165, x67164, x67163);
  nand n67167(x67167, x66472, x66542);
  nand n67168(x67168, x66471, x67170);
  nand n67169(x67169, x67168, x67167);
  nand n67171(x67171, x66472, x66543);
  nand n67172(x67172, x66471, x67174);
  nand n67173(x67173, x67172, x67171);
  nand n67175(x67175, x66472, x66544);
  nand n67176(x67176, x66471, x67178);
  nand n67177(x67177, x67176, x67175);
  nand n67179(x67179, x66472, x66545);
  nand n67180(x67180, x66471, x67182);
  nand n67181(x67181, x67180, x67179);
  nand n67183(x67183, x66472, x66546);
  nand n67184(x67184, x66471, x67186);
  nand n67185(x67185, x67184, x67183);
  nand n67187(x67187, x66472, x66547);
  nand n67188(x67188, x66471, x67190);
  nand n67189(x67189, x67188, x67187);
  nand n67191(x67191, x66472, x66548);
  nand n67192(x67192, x66471, x67194);
  nand n67193(x67193, x67192, x67191);
  nand n67195(x67195, x66472, x66549);
  nand n67196(x67196, x66471, x67198);
  nand n67197(x67197, x67196, x67195);
  nand n67199(x67199, x66472, x66550);
  nand n67200(x67200, x66471, x67202);
  nand n67201(x67201, x67200, x67199);
  nand n67203(x67203, x66472, x66551);
  nand n67204(x67204, x66471, x67206);
  nand n67205(x67205, x67204, x67203);
  nand n67207(x67207, x66472, x66552);
  nand n67208(x67208, x66471, x67210);
  nand n67209(x67209, x67208, x67207);
  nand n67211(x67211, x66472, x66553);
  nand n67212(x67212, x66471, x67214);
  nand n67213(x67213, x67212, x67211);
  nand n67215(x67215, x66472, x66554);
  nand n67216(x67216, x66471, x67218);
  nand n67217(x67217, x67216, x67215);
  nand n67219(x67219, x66472, x66555);
  nand n67220(x67220, x66471, x67222);
  nand n67221(x67221, x67220, x67219);
  nand n67223(x67223, x66472, x66556);
  nand n67224(x67224, x66471, x67226);
  nand n67225(x67225, x67224, x67223);
  nand n67227(x67227, x66472, x66557);
  nand n67228(x67228, x66471, x67230);
  nand n67229(x67229, x67228, x67227);
  nand n67231(x67231, x66472, x66558);
  nand n67232(x67232, x66471, x67234);
  nand n67233(x67233, x67232, x67231);
  nand n67235(x67235, x66472, x66559);
  nand n67236(x67236, x66471, x67238);
  nand n67237(x67237, x67236, x67235);
  nand n67239(x67239, x66472, x66560);
  nand n67240(x67240, x66471, x67242);
  nand n67241(x67241, x67240, x67239);
  nand n67243(x67243, x66472, x66561);
  nand n67244(x67244, x66471, x67246);
  nand n67245(x67245, x67244, x67243);
  nand n67247(x67247, x66472, x66562);
  nand n67248(x67248, x66471, x67250);
  nand n67249(x67249, x67248, x67247);
  nand n67251(x67251, x66472, x66563);
  nand n67252(x67252, x66471, x67254);
  nand n67253(x67253, x67252, x67251);
  nand n67255(x67255, x66472, x66564);
  nand n67256(x67256, x66471, x67258);
  nand n67257(x67257, x67256, x67255);
  nand n67259(x67259, x66472, x66565);
  nand n67260(x67260, x66471, x67262);
  nand n67261(x67261, x67260, x67259);
  nand n67263(x67263, x66472, x66566);
  nand n67264(x67264, x66471, x67266);
  nand n67265(x67265, x67264, x67263);
  nand n67267(x67267, x66472, x66567);
  nand n67268(x67268, x66471, x67270);
  nand n67269(x67269, x67268, x67267);
  nand n67271(x67271, x66472, x66568);
  nand n67272(x67272, x66471, x67274);
  nand n67273(x67273, x67272, x67271);
  nand n67275(x67275, x66472, x66569);
  nand n67276(x67276, x66471, x67278);
  nand n67277(x67277, x67276, x67275);
  nand n67279(x67279, x66472, x66570);
  nand n67280(x67280, x66471, x67282);
  nand n67281(x67281, x67280, x67279);
  nand n67283(x67283, x66472, x66571);
  nand n67284(x67284, x66471, x67286);
  nand n67285(x67285, x67284, x67283);
  nand n67287(x67287, x66472, x66572);
  nand n67288(x67288, x66471, x67290);
  nand n67289(x67289, x67288, x67287);
  nand n67291(x67291, x66472, x66573);
  nand n67292(x67292, x66471, x67294);
  nand n67293(x67293, x67292, x67291);
  nand n67295(x67295, x66472, x66574);
  nand n67296(x67296, x66471, x67298);
  nand n67297(x67297, x67296, x67295);
  nand n67299(x67299, x66472, x66575);
  nand n67300(x67300, x66471, x67302);
  nand n67301(x67301, x67300, x67299);
  nand n67303(x67303, x66472, x66576);
  nand n67304(x67304, x66471, x67306);
  nand n67305(x67305, x67304, x67303);
  nand n67307(x67307, x66472, x66577);
  nand n67308(x67308, x66471, x67310);
  nand n67309(x67309, x67308, x67307);
  nand n67311(x67311, x66472, x66578);
  nand n67312(x67312, x66471, x67314);
  nand n67313(x67313, x67312, x67311);
  nand n67315(x67315, x66472, x66579);
  nand n67316(x67316, x66471, x67318);
  nand n67317(x67317, x67316, x67315);
  nand n67319(x67319, x66472, x66580);
  nand n67320(x67320, x66471, x67322);
  nand n67321(x67321, x67320, x67319);
  nand n67323(x67323, x66472, x66581);
  nand n67324(x67324, x66471, x67326);
  nand n67325(x67325, x67324, x67323);
  nand n67327(x67327, x66472, x66582);
  nand n67328(x67328, x66471, x67330);
  nand n67329(x67329, x67328, x67327);
  nand n67331(x67331, x66472, x66583);
  nand n67332(x67332, x66471, x67334);
  nand n67333(x67333, x67332, x67331);
  nand n67335(x67335, x66472, x66584);
  nand n67336(x67336, x66471, x67338);
  nand n67337(x67337, x67336, x67335);
  nand n67339(x67339, x66472, x66585);
  nand n67340(x67340, x66471, x67342);
  nand n67341(x67341, x67340, x67339);
  nand n67343(x67343, x66472, x66586);
  nand n67344(x67344, x66471, x67346);
  nand n67345(x67345, x67344, x67343);
  nand n67347(x67347, x66472, x66587);
  nand n67348(x67348, x66471, x67350);
  nand n67349(x67349, x67348, x67347);
  nand n67351(x67351, x66472, x66588);
  nand n67352(x67352, x66471, x67354);
  nand n67353(x67353, x67352, x67351);
  nand n67355(x67355, x66472, x66589);
  nand n67356(x67356, x66471, x67358);
  nand n67357(x67357, x67356, x67355);
  nand n67359(x67359, x66472, x66590);
  nand n67360(x67360, x66471, x67362);
  nand n67361(x67361, x67360, x67359);
  nand n67363(x67363, x66472, x66591);
  nand n67364(x67364, x66471, x67366);
  nand n67365(x67365, x67364, x67363);
  nand n67367(x67367, x66472, x66592);
  nand n67368(x67368, x66471, x67370);
  nand n67369(x67369, x67368, x67367);
  nand n67371(x67371, x66472, x66593);
  nand n67372(x67372, x66471, x67374);
  nand n67373(x67373, x67372, x67371);
  nand n67375(x67375, x66472, x66594);
  nand n67376(x67376, x66471, x67378);
  nand n67377(x67377, x67376, x67375);
  nand n67379(x67379, x66472, x66595);
  nand n67380(x67380, x66471, x67382);
  nand n67381(x67381, x67380, x67379);
  nand n67383(x67383, x66472, x66596);
  nand n67384(x67384, x66471, x67386);
  nand n67385(x67385, x67384, x67383);
  nand n67387(x67387, x66472, x66597);
  nand n67388(x67388, x66471, x67390);
  nand n67389(x67389, x67388, x67387);
  nand n67391(x67391, x66472, x66598);
  nand n67392(x67392, x66471, x67394);
  nand n67393(x67393, x67392, x67391);
  nand n67395(x67395, x66472, x66599);
  nand n67396(x67396, x66471, x67398);
  nand n67397(x67397, x67396, x67395);
  nand n67399(x67399, x66472, x66600);
  nand n67400(x67400, x66471, x67402);
  nand n67401(x67401, x67400, x67399);
  nand n67403(x67403, x83372, x66601);
  nand n67404(x67404, x66472, x83372);
  nand n67406(x67406, x66472, x78109);
  nand n67407(x67407, x66471, x67409);
  nand n67408(x67408, x67407, x67406);
  nand n67410(x67410, x66472, x78112);
  nand n67411(x67411, x66471, x67413);
  nand n67412(x67412, x67411, x67410);
  nand n67414(x67414, x66472, x78115);
  nand n67415(x67415, x66471, x67417);
  nand n67416(x67416, x67415, x67414);
  nand n67418(x67418, x66472, x78118);
  nand n67419(x67419, x66471, x67421);
  nand n67420(x67420, x67419, x67418);
  nand n67422(x67422, x66472, x78121);
  nand n67423(x67423, x66471, x67425);
  nand n67424(x67424, x67423, x67422);
  nand n67426(x67426, x66472, x78124);
  nand n67427(x67427, x66471, x67429);
  nand n67428(x67428, x67427, x67426);
  nand n67430(x67430, x66472, x78145);
  nand n67431(x67431, x66471, x67433);
  nand n67432(x67432, x67431, x67430);
  nand n67434(x67434, x66472, x78148);
  nand n67435(x67435, x66471, x67437);
  nand n67436(x67436, x67435, x67434);
  nand n67438(x67438, x66472, x78151);
  nand n67439(x67439, x66471, x67441);
  nand n67440(x67440, x67439, x67438);
  nand n67442(x67442, x66472, x78154);
  nand n67443(x67443, x66471, x67445);
  nand n67444(x67444, x67443, x67442);
  nand n67446(x67446, x66472, x78157);
  nand n67447(x67447, x66471, x67449);
  nand n67448(x67448, x67447, x67446);
  nand n67450(x67450, x66472, x78160);
  nand n67451(x67451, x66471, x67453);
  nand n67452(x67452, x67451, x67450);
  nand n67454(x67454, x66472, x78163);
  nand n67455(x67455, x66471, x67457);
  nand n67456(x67456, x67455, x67454);
  nand n67458(x67458, x66472, x78166);
  nand n67459(x67459, x66471, x67461);
  nand n67460(x67460, x67459, x67458);
  nand n67462(x67462, x67403, x83372);
  nand n67464(x67464, x67594, x67463);
  nand n67595(x67595, x79441, x79345);
  nand n67597(x67597, x67596, x79600);
  nand n67598(x67598, x67597, x67595);
  nand n67599(x67599, x79441, x79348);
  nand n67600(x67600, x67596, x79603);
  nand n67601(x67601, x67600, x67599);
  nand n67602(x67602, x79441, x79351);
  nand n67603(x67603, x67596, x79606);
  nand n67604(x67604, x67603, x67602);
  nand n67605(x67605, x79441, x79354);
  nand n67606(x67606, x67596, x79609);
  nand n67607(x67607, x67606, x67605);
  nand n67608(x67608, x79441, x79357);
  nand n67609(x67609, x67596, x79612);
  nand n67610(x67610, x67609, x67608);
  nand n67611(x67611, x79441, x79360);
  nand n67612(x67612, x67596, x79615);
  nand n67613(x67613, x67612, x67611);
  nand n67614(x67614, x79441, x79363);
  nand n67615(x67615, x67596, x79618);
  nand n67616(x67616, x67615, x67614);
  nand n67617(x67617, x79441, x79366);
  nand n67618(x67618, x67596, x79621);
  nand n67619(x67619, x67618, x67617);
  nand n67620(x67620, x79441, x79369);
  nand n67621(x67621, x67596, x79624);
  nand n67622(x67622, x67621, x67620);
  nand n67623(x67623, x79441, x79372);
  nand n67624(x67624, x67596, x79627);
  nand n67625(x67625, x67624, x67623);
  nand n67626(x67626, x79441, x79375);
  nand n67627(x67627, x67596, x79630);
  nand n67628(x67628, x67627, x67626);
  nand n67629(x67629, x79441, x79378);
  nand n67630(x67630, x67596, x79633);
  nand n67631(x67631, x67630, x67629);
  nand n67632(x67632, x79441, x79381);
  nand n67633(x67633, x67596, x79636);
  nand n67634(x67634, x67633, x67632);
  nand n67635(x67635, x79441, x79384);
  nand n67636(x67636, x67596, x79639);
  nand n67637(x67637, x67636, x67635);
  nand n67638(x67638, x79441, x79387);
  nand n67639(x67639, x67596, x79642);
  nand n67640(x67640, x67639, x67638);
  nand n67641(x67641, x79441, x79390);
  nand n67642(x67642, x67596, x79645);
  nand n67643(x67643, x67642, x67641);
  nand n67644(x67644, x79441, x79393);
  nand n67645(x67645, x67596, x79648);
  nand n67646(x67646, x67645, x67644);
  nand n67647(x67647, x79441, x79396);
  nand n67648(x67648, x67596, x79651);
  nand n67649(x67649, x67648, x67647);
  nand n67650(x67650, x79441, x79399);
  nand n67651(x67651, x67596, x79654);
  nand n67652(x67652, x67651, x67650);
  nand n67653(x67653, x79441, x79402);
  nand n67654(x67654, x67596, x79657);
  nand n67655(x67655, x67654, x67653);
  nand n67656(x67656, x79441, x79405);
  nand n67657(x67657, x67596, x79660);
  nand n67658(x67658, x67657, x67656);
  nand n67659(x67659, x79441, x79408);
  nand n67660(x67660, x67596, x79663);
  nand n67661(x67661, x67660, x67659);
  nand n67662(x67662, x79441, x79411);
  nand n67663(x67663, x67596, x79666);
  nand n67664(x67664, x67663, x67662);
  nand n67665(x67665, x79441, x79414);
  nand n67666(x67666, x67596, x79669);
  nand n67667(x67667, x67666, x67665);
  nand n67668(x67668, x79441, x79417);
  nand n67669(x67669, x67596, x79672);
  nand n67670(x67670, x67669, x67668);
  nand n67671(x67671, x79441, x79420);
  nand n67672(x67672, x67596, x79675);
  nand n67673(x67673, x67672, x67671);
  nand n67674(x67674, x79441, x79423);
  nand n67675(x67675, x67596, x79678);
  nand n67676(x67676, x67675, x67674);
  nand n67677(x67677, x79441, x79426);
  nand n67678(x67678, x67596, x79681);
  nand n67679(x67679, x67678, x67677);
  nand n67680(x67680, x79441, x79429);
  nand n67681(x67681, x67596, x79684);
  nand n67682(x67682, x67681, x67680);
  nand n67683(x67683, x79441, x79432);
  nand n67684(x67684, x67596, x79687);
  nand n67685(x67685, x67684, x67683);
  nand n67686(x67686, x79441, x79435);
  nand n67687(x67687, x67596, x79690);
  nand n67688(x67688, x67687, x67686);
  nand n67689(x67689, x79441, x79438);
  nand n67690(x67690, x67596, x79693);
  nand n67691(x67691, x67690, x67689);
  nand n67692(x67692, x67596, x79894);
  nand n67693(x67693, x67692, x67595);
  nand n67694(x67694, x67596, x79897);
  nand n67695(x67695, x67694, x67599);
  nand n67696(x67696, x67596, x79900);
  nand n67697(x67697, x67696, x67602);
  nand n67698(x67698, x67596, x79903);
  nand n67699(x67699, x67698, x67605);
  nand n67700(x67700, x67596, x79906);
  nand n67701(x67701, x67700, x67608);
  nand n67702(x67702, x67596, x79909);
  nand n67703(x67703, x67702, x67611);
  nand n67704(x67704, x67596, x79912);
  nand n67705(x67705, x67704, x67614);
  nand n67706(x67706, x67596, x79915);
  nand n67707(x67707, x67706, x67617);
  nand n67708(x67708, x67596, x79918);
  nand n67709(x67709, x67708, x67620);
  nand n67710(x67710, x67596, x79921);
  nand n67711(x67711, x67710, x67623);
  nand n67712(x67712, x67596, x79924);
  nand n67713(x67713, x67712, x67626);
  nand n67714(x67714, x67596, x79927);
  nand n67715(x67715, x67714, x67629);
  nand n67716(x67716, x67596, x79930);
  nand n67717(x67717, x67716, x67632);
  nand n67718(x67718, x67596, x79933);
  nand n67719(x67719, x67718, x67635);
  nand n67720(x67720, x67596, x79936);
  nand n67721(x67721, x67720, x67638);
  nand n67722(x67722, x67596, x79939);
  nand n67723(x67723, x67722, x67641);
  nand n67724(x67724, x67596, x79942);
  nand n67725(x67725, x67724, x67644);
  nand n67726(x67726, x67596, x79945);
  nand n67727(x67727, x67726, x67647);
  nand n67728(x67728, x67596, x79948);
  nand n67729(x67729, x67728, x67650);
  nand n67730(x67730, x67596, x79951);
  nand n67731(x67731, x67730, x67653);
  nand n67732(x67732, x67596, x79954);
  nand n67733(x67733, x67732, x67656);
  nand n67734(x67734, x67596, x79957);
  nand n67735(x67735, x67734, x67659);
  nand n67736(x67736, x67596, x79960);
  nand n67737(x67737, x67736, x67662);
  nand n67738(x67738, x67596, x79963);
  nand n67739(x67739, x67738, x67665);
  nand n67740(x67740, x67596, x79966);
  nand n67741(x67741, x67740, x67668);
  nand n67742(x67742, x67596, x79969);
  nand n67743(x67743, x67742, x67671);
  nand n67744(x67744, x67596, x79972);
  nand n67745(x67745, x67744, x67674);
  nand n67746(x67746, x67596, x79975);
  nand n67747(x67747, x67746, x67677);
  nand n67748(x67748, x67596, x79978);
  nand n67749(x67749, x67748, x67680);
  nand n67750(x67750, x67596, x79981);
  nand n67751(x67751, x67750, x67683);
  nand n67752(x67752, x67596, x79984);
  nand n67753(x67753, x67752, x67686);
  nand n67754(x67754, x67596, x79987);
  nand n67755(x67755, x67754, x67689);
  nand n67756(x67756, x67596, x80188);
  nand n67757(x67757, x67756, x67595);
  nand n67758(x67758, x67596, x80191);
  nand n67759(x67759, x67758, x67599);
  nand n67760(x67760, x67596, x80194);
  nand n67761(x67761, x67760, x67602);
  nand n67762(x67762, x67596, x80197);
  nand n67763(x67763, x67762, x67605);
  nand n67764(x67764, x67596, x80200);
  nand n67765(x67765, x67764, x67608);
  nand n67766(x67766, x67596, x80203);
  nand n67767(x67767, x67766, x67611);
  nand n67768(x67768, x67596, x80206);
  nand n67769(x67769, x67768, x67614);
  nand n67770(x67770, x67596, x80209);
  nand n67771(x67771, x67770, x67617);
  nand n67772(x67772, x67596, x80212);
  nand n67773(x67773, x67772, x67620);
  nand n67774(x67774, x67596, x80215);
  nand n67775(x67775, x67774, x67623);
  nand n67776(x67776, x67596, x80218);
  nand n67777(x67777, x67776, x67626);
  nand n67778(x67778, x67596, x80221);
  nand n67779(x67779, x67778, x67629);
  nand n67780(x67780, x67596, x80224);
  nand n67781(x67781, x67780, x67632);
  nand n67782(x67782, x67596, x80227);
  nand n67783(x67783, x67782, x67635);
  nand n67784(x67784, x67596, x80230);
  nand n67785(x67785, x67784, x67638);
  nand n67786(x67786, x67596, x80233);
  nand n67787(x67787, x67786, x67641);
  nand n67788(x67788, x67596, x80236);
  nand n67789(x67789, x67788, x67644);
  nand n67790(x67790, x67596, x80239);
  nand n67791(x67791, x67790, x67647);
  nand n67792(x67792, x67596, x80242);
  nand n67793(x67793, x67792, x67650);
  nand n67794(x67794, x67596, x80245);
  nand n67795(x67795, x67794, x67653);
  nand n67796(x67796, x67596, x80248);
  nand n67797(x67797, x67796, x67656);
  nand n67798(x67798, x67596, x80251);
  nand n67799(x67799, x67798, x67659);
  nand n67800(x67800, x67596, x80254);
  nand n67801(x67801, x67800, x67662);
  nand n67802(x67802, x67596, x80257);
  nand n67803(x67803, x67802, x67665);
  nand n67804(x67804, x67596, x80260);
  nand n67805(x67805, x67804, x67668);
  nand n67806(x67806, x67596, x80263);
  nand n67807(x67807, x67806, x67671);
  nand n67808(x67808, x67596, x80266);
  nand n67809(x67809, x67808, x67674);
  nand n67810(x67810, x67596, x80269);
  nand n67811(x67811, x67810, x67677);
  nand n67812(x67812, x67596, x80272);
  nand n67813(x67813, x67812, x67680);
  nand n67814(x67814, x67596, x80275);
  nand n67815(x67815, x67814, x67683);
  nand n67816(x67816, x67596, x80278);
  nand n67817(x67817, x67816, x67686);
  nand n67818(x67818, x67596, x80281);
  nand n67819(x67819, x67818, x67689);
  nand n67820(x67820, x67596, x80482);
  nand n67821(x67821, x67820, x67595);
  nand n67822(x67822, x67596, x80485);
  nand n67823(x67823, x67822, x67599);
  nand n67824(x67824, x67596, x80488);
  nand n67825(x67825, x67824, x67602);
  nand n67826(x67826, x67596, x80491);
  nand n67827(x67827, x67826, x67605);
  nand n67828(x67828, x67596, x80494);
  nand n67829(x67829, x67828, x67608);
  nand n67830(x67830, x67596, x80497);
  nand n67831(x67831, x67830, x67611);
  nand n67832(x67832, x67596, x80500);
  nand n67833(x67833, x67832, x67614);
  nand n67834(x67834, x67596, x80503);
  nand n67835(x67835, x67834, x67617);
  nand n67836(x67836, x67596, x80506);
  nand n67837(x67837, x67836, x67620);
  nand n67838(x67838, x67596, x80509);
  nand n67839(x67839, x67838, x67623);
  nand n67840(x67840, x67596, x80512);
  nand n67841(x67841, x67840, x67626);
  nand n67842(x67842, x67596, x80515);
  nand n67843(x67843, x67842, x67629);
  nand n67844(x67844, x67596, x80518);
  nand n67845(x67845, x67844, x67632);
  nand n67846(x67846, x67596, x80521);
  nand n67847(x67847, x67846, x67635);
  nand n67848(x67848, x67596, x80524);
  nand n67849(x67849, x67848, x67638);
  nand n67850(x67850, x67596, x80527);
  nand n67851(x67851, x67850, x67641);
  nand n67852(x67852, x67596, x80530);
  nand n67853(x67853, x67852, x67644);
  nand n67854(x67854, x67596, x80533);
  nand n67855(x67855, x67854, x67647);
  nand n67856(x67856, x67596, x80536);
  nand n67857(x67857, x67856, x67650);
  nand n67858(x67858, x67596, x80539);
  nand n67859(x67859, x67858, x67653);
  nand n67860(x67860, x67596, x80542);
  nand n67861(x67861, x67860, x67656);
  nand n67862(x67862, x67596, x80545);
  nand n67863(x67863, x67862, x67659);
  nand n67864(x67864, x67596, x80548);
  nand n67865(x67865, x67864, x67662);
  nand n67866(x67866, x67596, x80551);
  nand n67867(x67867, x67866, x67665);
  nand n67868(x67868, x67596, x80554);
  nand n67869(x67869, x67868, x67668);
  nand n67870(x67870, x67596, x80557);
  nand n67871(x67871, x67870, x67671);
  nand n67872(x67872, x67596, x80560);
  nand n67873(x67873, x67872, x67674);
  nand n67874(x67874, x67596, x80563);
  nand n67875(x67875, x67874, x67677);
  nand n67876(x67876, x67596, x80566);
  nand n67877(x67877, x67876, x67680);
  nand n67878(x67878, x67596, x80569);
  nand n67879(x67879, x67878, x67683);
  nand n67880(x67880, x67596, x80572);
  nand n67881(x67881, x67880, x67686);
  nand n67882(x67882, x67596, x80575);
  nand n67883(x67883, x67882, x67689);
  nand n67884(x67884, x67465, x67466);
  nand n67885(x67885, x67464, x67887);
  nand n67886(x67886, x67885, x67884);
  nand n67888(x67888, x67465, x67467);
  nand n67889(x67889, x67464, x67891);
  nand n67890(x67890, x67889, x67888);
  nand n67892(x67892, x67465, x67468);
  nand n67893(x67893, x67464, x67895);
  nand n67894(x67894, x67893, x67892);
  nand n67896(x67896, x67465, x67469);
  nand n67897(x67897, x67464, x67899);
  nand n67898(x67898, x67897, x67896);
  nand n67900(x67900, x67465, x67470);
  nand n67901(x67901, x67464, x67903);
  nand n67902(x67902, x67901, x67900);
  nand n67904(x67904, x67465, x67471);
  nand n67905(x67905, x67464, x67907);
  nand n67906(x67906, x67905, x67904);
  nand n67908(x67908, x67465, x67472);
  nand n67909(x67909, x67464, x67911);
  nand n67910(x67910, x67909, x67908);
  nand n67912(x67912, x67465, x67473);
  nand n67913(x67913, x67464, x67915);
  nand n67914(x67914, x67913, x67912);
  nand n67916(x67916, x67465, x67474);
  nand n67917(x67917, x67464, x67919);
  nand n67918(x67918, x67917, x67916);
  nand n67920(x67920, x67465, x67475);
  nand n67921(x67921, x67464, x67923);
  nand n67922(x67922, x67921, x67920);
  nand n67924(x67924, x67465, x67476);
  nand n67925(x67925, x67464, x67927);
  nand n67926(x67926, x67925, x67924);
  nand n67928(x67928, x67465, x67477);
  nand n67929(x67929, x67464, x67931);
  nand n67930(x67930, x67929, x67928);
  nand n67932(x67932, x67465, x67478);
  nand n67933(x67933, x67464, x67935);
  nand n67934(x67934, x67933, x67932);
  nand n67936(x67936, x67465, x67479);
  nand n67937(x67937, x67464, x67939);
  nand n67938(x67938, x67937, x67936);
  nand n67940(x67940, x67465, x67480);
  nand n67941(x67941, x67464, x67943);
  nand n67942(x67942, x67941, x67940);
  nand n67944(x67944, x67465, x67481);
  nand n67945(x67945, x67464, x67947);
  nand n67946(x67946, x67945, x67944);
  nand n67948(x67948, x67465, x67482);
  nand n67949(x67949, x67464, x67951);
  nand n67950(x67950, x67949, x67948);
  nand n67952(x67952, x67465, x67483);
  nand n67953(x67953, x67464, x67955);
  nand n67954(x67954, x67953, x67952);
  nand n67956(x67956, x67465, x67484);
  nand n67957(x67957, x67464, x67959);
  nand n67958(x67958, x67957, x67956);
  nand n67960(x67960, x67465, x67485);
  nand n67961(x67961, x67464, x67963);
  nand n67962(x67962, x67961, x67960);
  nand n67964(x67964, x67465, x67486);
  nand n67965(x67965, x67464, x67967);
  nand n67966(x67966, x67965, x67964);
  nand n67968(x67968, x67465, x67487);
  nand n67969(x67969, x67464, x67971);
  nand n67970(x67970, x67969, x67968);
  nand n67972(x67972, x67465, x67488);
  nand n67973(x67973, x67464, x67975);
  nand n67974(x67974, x67973, x67972);
  nand n67976(x67976, x67465, x67489);
  nand n67977(x67977, x67464, x67979);
  nand n67978(x67978, x67977, x67976);
  nand n67980(x67980, x67465, x67490);
  nand n67981(x67981, x67464, x67983);
  nand n67982(x67982, x67981, x67980);
  nand n67984(x67984, x67465, x67491);
  nand n67985(x67985, x67464, x67987);
  nand n67986(x67986, x67985, x67984);
  nand n67988(x67988, x67465, x67492);
  nand n67989(x67989, x67464, x67991);
  nand n67990(x67990, x67989, x67988);
  nand n67992(x67992, x67465, x67493);
  nand n67993(x67993, x67464, x67995);
  nand n67994(x67994, x67993, x67992);
  nand n67996(x67996, x67465, x67494);
  nand n67997(x67997, x67464, x67999);
  nand n67998(x67998, x67997, x67996);
  nand n68000(x68000, x67465, x67495);
  nand n68001(x68001, x67464, x68003);
  nand n68002(x68002, x68001, x68000);
  nand n68004(x68004, x67465, x67496);
  nand n68005(x68005, x67464, x68007);
  nand n68006(x68006, x68005, x68004);
  nand n68008(x68008, x67465, x67497);
  nand n68009(x68009, x67464, x68011);
  nand n68010(x68010, x68009, x68008);
  nand n68012(x68012, x67465, x67498);
  nand n68013(x68013, x67464, x68015);
  nand n68014(x68014, x68013, x68012);
  nand n68016(x68016, x67465, x67499);
  nand n68017(x68017, x67464, x68019);
  nand n68018(x68018, x68017, x68016);
  nand n68020(x68020, x67465, x67500);
  nand n68021(x68021, x67464, x68023);
  nand n68022(x68022, x68021, x68020);
  nand n68024(x68024, x67465, x67501);
  nand n68025(x68025, x67464, x68027);
  nand n68026(x68026, x68025, x68024);
  nand n68028(x68028, x67465, x67502);
  nand n68029(x68029, x67464, x68031);
  nand n68030(x68030, x68029, x68028);
  nand n68032(x68032, x67465, x67503);
  nand n68033(x68033, x67464, x68035);
  nand n68034(x68034, x68033, x68032);
  nand n68036(x68036, x67465, x67504);
  nand n68037(x68037, x67464, x68039);
  nand n68038(x68038, x68037, x68036);
  nand n68040(x68040, x67465, x67505);
  nand n68041(x68041, x67464, x68043);
  nand n68042(x68042, x68041, x68040);
  nand n68044(x68044, x67465, x67506);
  nand n68045(x68045, x67464, x68047);
  nand n68046(x68046, x68045, x68044);
  nand n68048(x68048, x67465, x67507);
  nand n68049(x68049, x67464, x68051);
  nand n68050(x68050, x68049, x68048);
  nand n68052(x68052, x67465, x67508);
  nand n68053(x68053, x67464, x68055);
  nand n68054(x68054, x68053, x68052);
  nand n68056(x68056, x67465, x67509);
  nand n68057(x68057, x67464, x68059);
  nand n68058(x68058, x68057, x68056);
  nand n68060(x68060, x67465, x67510);
  nand n68061(x68061, x67464, x68063);
  nand n68062(x68062, x68061, x68060);
  nand n68064(x68064, x67465, x67511);
  nand n68065(x68065, x67464, x68067);
  nand n68066(x68066, x68065, x68064);
  nand n68068(x68068, x67465, x67512);
  nand n68069(x68069, x67464, x68071);
  nand n68070(x68070, x68069, x68068);
  nand n68072(x68072, x67465, x67513);
  nand n68073(x68073, x67464, x68075);
  nand n68074(x68074, x68073, x68072);
  nand n68076(x68076, x67465, x67514);
  nand n68077(x68077, x67464, x68079);
  nand n68078(x68078, x68077, x68076);
  nand n68080(x68080, x67465, x67515);
  nand n68081(x68081, x67464, x68083);
  nand n68082(x68082, x68081, x68080);
  nand n68084(x68084, x67465, x67516);
  nand n68085(x68085, x67464, x68087);
  nand n68086(x68086, x68085, x68084);
  nand n68088(x68088, x67465, x67517);
  nand n68089(x68089, x67464, x68091);
  nand n68090(x68090, x68089, x68088);
  nand n68092(x68092, x67465, x67518);
  nand n68093(x68093, x67464, x68095);
  nand n68094(x68094, x68093, x68092);
  nand n68096(x68096, x67465, x67519);
  nand n68097(x68097, x67464, x68099);
  nand n68098(x68098, x68097, x68096);
  nand n68100(x68100, x67465, x67520);
  nand n68101(x68101, x67464, x68103);
  nand n68102(x68102, x68101, x68100);
  nand n68104(x68104, x67465, x67521);
  nand n68105(x68105, x67464, x68107);
  nand n68106(x68106, x68105, x68104);
  nand n68108(x68108, x67465, x67522);
  nand n68109(x68109, x67464, x68111);
  nand n68110(x68110, x68109, x68108);
  nand n68112(x68112, x67465, x67523);
  nand n68113(x68113, x67464, x68115);
  nand n68114(x68114, x68113, x68112);
  nand n68116(x68116, x67465, x67524);
  nand n68117(x68117, x67464, x68119);
  nand n68118(x68118, x68117, x68116);
  nand n68120(x68120, x67465, x67525);
  nand n68121(x68121, x67464, x68123);
  nand n68122(x68122, x68121, x68120);
  nand n68124(x68124, x67465, x67526);
  nand n68125(x68125, x67464, x68127);
  nand n68126(x68126, x68125, x68124);
  nand n68128(x68128, x67465, x67527);
  nand n68129(x68129, x67464, x68131);
  nand n68130(x68130, x68129, x68128);
  nand n68132(x68132, x67465, x67528);
  nand n68133(x68133, x67464, x68135);
  nand n68134(x68134, x68133, x68132);
  nand n68136(x68136, x67465, x67529);
  nand n68137(x68137, x67464, x68139);
  nand n68138(x68138, x68137, x68136);
  nand n68140(x68140, x67465, x67530);
  nand n68141(x68141, x67464, x68143);
  nand n68142(x68142, x68141, x68140);
  nand n68144(x68144, x67465, x67531);
  nand n68145(x68145, x67464, x68147);
  nand n68146(x68146, x68145, x68144);
  nand n68148(x68148, x67465, x67532);
  nand n68149(x68149, x67464, x68151);
  nand n68150(x68150, x68149, x68148);
  nand n68152(x68152, x67465, x67533);
  nand n68153(x68153, x67464, x68155);
  nand n68154(x68154, x68153, x68152);
  nand n68156(x68156, x67465, x67534);
  nand n68157(x68157, x67464, x68159);
  nand n68158(x68158, x68157, x68156);
  nand n68160(x68160, x67465, x67535);
  nand n68161(x68161, x67464, x68163);
  nand n68162(x68162, x68161, x68160);
  nand n68164(x68164, x67465, x67536);
  nand n68165(x68165, x67464, x68167);
  nand n68166(x68166, x68165, x68164);
  nand n68168(x68168, x67465, x67537);
  nand n68169(x68169, x67464, x68171);
  nand n68170(x68170, x68169, x68168);
  nand n68172(x68172, x67465, x67538);
  nand n68173(x68173, x67464, x68175);
  nand n68174(x68174, x68173, x68172);
  nand n68176(x68176, x67465, x67539);
  nand n68177(x68177, x67464, x68179);
  nand n68178(x68178, x68177, x68176);
  nand n68180(x68180, x67465, x67540);
  nand n68181(x68181, x67464, x68183);
  nand n68182(x68182, x68181, x68180);
  nand n68184(x68184, x67465, x67541);
  nand n68185(x68185, x67464, x68187);
  nand n68186(x68186, x68185, x68184);
  nand n68188(x68188, x67465, x67542);
  nand n68189(x68189, x67464, x68191);
  nand n68190(x68190, x68189, x68188);
  nand n68192(x68192, x67465, x67543);
  nand n68193(x68193, x67464, x68195);
  nand n68194(x68194, x68193, x68192);
  nand n68196(x68196, x67465, x67544);
  nand n68197(x68197, x67464, x68199);
  nand n68198(x68198, x68197, x68196);
  nand n68200(x68200, x67465, x67545);
  nand n68201(x68201, x67464, x68203);
  nand n68202(x68202, x68201, x68200);
  nand n68204(x68204, x67465, x67546);
  nand n68205(x68205, x67464, x68207);
  nand n68206(x68206, x68205, x68204);
  nand n68208(x68208, x67465, x67547);
  nand n68209(x68209, x67464, x68211);
  nand n68210(x68210, x68209, x68208);
  nand n68212(x68212, x67465, x67548);
  nand n68213(x68213, x67464, x68215);
  nand n68214(x68214, x68213, x68212);
  nand n68216(x68216, x67465, x67549);
  nand n68217(x68217, x67464, x68219);
  nand n68218(x68218, x68217, x68216);
  nand n68220(x68220, x67465, x67550);
  nand n68221(x68221, x67464, x68223);
  nand n68222(x68222, x68221, x68220);
  nand n68224(x68224, x67465, x67551);
  nand n68225(x68225, x67464, x68227);
  nand n68226(x68226, x68225, x68224);
  nand n68228(x68228, x67465, x67552);
  nand n68229(x68229, x67464, x68231);
  nand n68230(x68230, x68229, x68228);
  nand n68232(x68232, x67465, x67553);
  nand n68233(x68233, x67464, x68235);
  nand n68234(x68234, x68233, x68232);
  nand n68236(x68236, x67465, x67554);
  nand n68237(x68237, x67464, x68239);
  nand n68238(x68238, x68237, x68236);
  nand n68240(x68240, x67465, x67555);
  nand n68241(x68241, x67464, x68243);
  nand n68242(x68242, x68241, x68240);
  nand n68244(x68244, x67465, x67556);
  nand n68245(x68245, x67464, x68247);
  nand n68246(x68246, x68245, x68244);
  nand n68248(x68248, x67465, x67557);
  nand n68249(x68249, x67464, x68251);
  nand n68250(x68250, x68249, x68248);
  nand n68252(x68252, x67465, x67558);
  nand n68253(x68253, x67464, x68255);
  nand n68254(x68254, x68253, x68252);
  nand n68256(x68256, x67465, x67559);
  nand n68257(x68257, x67464, x68259);
  nand n68258(x68258, x68257, x68256);
  nand n68260(x68260, x67465, x67560);
  nand n68261(x68261, x67464, x68263);
  nand n68262(x68262, x68261, x68260);
  nand n68264(x68264, x67465, x67561);
  nand n68265(x68265, x67464, x68267);
  nand n68266(x68266, x68265, x68264);
  nand n68268(x68268, x67465, x67562);
  nand n68269(x68269, x67464, x68271);
  nand n68270(x68270, x68269, x68268);
  nand n68272(x68272, x67465, x67563);
  nand n68273(x68273, x67464, x68275);
  nand n68274(x68274, x68273, x68272);
  nand n68276(x68276, x67465, x67564);
  nand n68277(x68277, x67464, x68279);
  nand n68278(x68278, x68277, x68276);
  nand n68280(x68280, x67465, x67565);
  nand n68281(x68281, x67464, x68283);
  nand n68282(x68282, x68281, x68280);
  nand n68284(x68284, x67465, x67566);
  nand n68285(x68285, x67464, x68287);
  nand n68286(x68286, x68285, x68284);
  nand n68288(x68288, x67465, x67567);
  nand n68289(x68289, x67464, x68291);
  nand n68290(x68290, x68289, x68288);
  nand n68292(x68292, x67465, x67568);
  nand n68293(x68293, x67464, x68295);
  nand n68294(x68294, x68293, x68292);
  nand n68296(x68296, x67465, x67569);
  nand n68297(x68297, x67464, x68299);
  nand n68298(x68298, x68297, x68296);
  nand n68300(x68300, x67465, x67570);
  nand n68301(x68301, x67464, x68303);
  nand n68302(x68302, x68301, x68300);
  nand n68304(x68304, x67465, x67571);
  nand n68305(x68305, x67464, x68307);
  nand n68306(x68306, x68305, x68304);
  nand n68308(x68308, x67465, x67572);
  nand n68309(x68309, x67464, x68311);
  nand n68310(x68310, x68309, x68308);
  nand n68312(x68312, x67465, x67573);
  nand n68313(x68313, x67464, x68315);
  nand n68314(x68314, x68313, x68312);
  nand n68316(x68316, x67465, x67574);
  nand n68317(x68317, x67464, x68319);
  nand n68318(x68318, x68317, x68316);
  nand n68320(x68320, x67465, x67575);
  nand n68321(x68321, x67464, x68323);
  nand n68322(x68322, x68321, x68320);
  nand n68324(x68324, x67465, x67576);
  nand n68325(x68325, x67464, x68327);
  nand n68326(x68326, x68325, x68324);
  nand n68328(x68328, x67465, x67577);
  nand n68329(x68329, x67464, x68331);
  nand n68330(x68330, x68329, x68328);
  nand n68332(x68332, x67465, x67578);
  nand n68333(x68333, x67464, x68335);
  nand n68334(x68334, x68333, x68332);
  nand n68336(x68336, x67465, x67579);
  nand n68337(x68337, x67464, x68339);
  nand n68338(x68338, x68337, x68336);
  nand n68340(x68340, x67465, x67580);
  nand n68341(x68341, x67464, x68343);
  nand n68342(x68342, x68341, x68340);
  nand n68344(x68344, x67465, x67581);
  nand n68345(x68345, x67464, x68347);
  nand n68346(x68346, x68345, x68344);
  nand n68348(x68348, x67465, x67582);
  nand n68349(x68349, x67464, x68351);
  nand n68350(x68350, x68349, x68348);
  nand n68352(x68352, x67465, x67583);
  nand n68353(x68353, x67464, x68355);
  nand n68354(x68354, x68353, x68352);
  nand n68356(x68356, x67465, x67584);
  nand n68357(x68357, x67464, x68359);
  nand n68358(x68358, x68357, x68356);
  nand n68360(x68360, x67465, x67585);
  nand n68361(x68361, x67464, x68363);
  nand n68362(x68362, x68361, x68360);
  nand n68364(x68364, x67465, x67586);
  nand n68365(x68365, x67464, x68367);
  nand n68366(x68366, x68365, x68364);
  nand n68368(x68368, x67465, x67587);
  nand n68369(x68369, x67464, x68371);
  nand n68370(x68370, x68369, x68368);
  nand n68372(x68372, x67465, x67588);
  nand n68373(x68373, x67464, x68375);
  nand n68374(x68374, x68373, x68372);
  nand n68376(x68376, x67465, x67589);
  nand n68377(x68377, x67464, x68379);
  nand n68378(x68378, x68377, x68376);
  nand n68380(x68380, x67465, x67590);
  nand n68381(x68381, x67464, x68383);
  nand n68382(x68382, x68381, x68380);
  nand n68384(x68384, x67465, x67591);
  nand n68385(x68385, x67464, x68387);
  nand n68386(x68386, x68385, x68384);
  nand n68388(x68388, x67465, x67592);
  nand n68389(x68389, x67464, x68391);
  nand n68390(x68390, x68389, x68388);
  nand n68392(x68392, x67465, x67593);
  nand n68393(x68393, x67464, x68395);
  nand n68394(x68394, x68393, x68392);
  nand n68396(x68396, x83377, x67594);
  nand n68397(x68397, x67465, x83377);
  nand n68399(x68399, x67465, x79444);
  nand n68400(x68400, x67464, x68402);
  nand n68401(x68401, x68400, x68399);
  nand n68403(x68403, x67465, x79447);
  nand n68404(x68404, x67464, x68406);
  nand n68405(x68405, x68404, x68403);
  nand n68407(x68407, x67465, x79450);
  nand n68408(x68408, x67464, x68410);
  nand n68409(x68409, x68408, x68407);
  nand n68411(x68411, x67465, x79453);
  nand n68412(x68412, x67464, x68414);
  nand n68413(x68413, x68412, x68411);
  nand n68415(x68415, x67465, x79456);
  nand n68416(x68416, x67464, x68418);
  nand n68417(x68417, x68416, x68415);
  nand n68419(x68419, x67465, x79459);
  nand n68420(x68420, x67464, x68422);
  nand n68421(x68421, x68420, x68419);
  nand n68423(x68423, x67465, x79480);
  nand n68424(x68424, x67464, x68426);
  nand n68425(x68425, x68424, x68423);
  nand n68427(x68427, x67465, x79483);
  nand n68428(x68428, x67464, x68430);
  nand n68429(x68429, x68428, x68427);
  nand n68431(x68431, x67465, x79486);
  nand n68432(x68432, x67464, x68434);
  nand n68433(x68433, x68432, x68431);
  nand n68435(x68435, x67465, x79489);
  nand n68436(x68436, x67464, x68438);
  nand n68437(x68437, x68436, x68435);
  nand n68439(x68439, x67465, x79492);
  nand n68440(x68440, x67464, x68442);
  nand n68441(x68441, x68440, x68439);
  nand n68443(x68443, x67465, x79495);
  nand n68444(x68444, x67464, x68446);
  nand n68445(x68445, x68444, x68443);
  nand n68447(x68447, x67465, x79498);
  nand n68448(x68448, x67464, x68450);
  nand n68449(x68449, x68448, x68447);
  nand n68451(x68451, x67465, x79501);
  nand n68452(x68452, x67464, x68454);
  nand n68453(x68453, x68452, x68451);
  nand n68455(x68455, x68396, x83377);
  nand n68456(x68456, x67462, x68455);
  nand n68457(x68457, x60841, x61424);
  nand n68460(x68460, x68459, x62930);
  nand n68462(x68462, x68461, x68458);
  nand n68463(x68463, x15225, x1107);
  nand n68465(x68465, x68464, x1037);
  nand n68466(x68466, x71449, x1143);
  nand n68468(x68468, x68467, x68465);
  nand n68472(x68472, x68471, x68618);
  nand n68474(x68474, x68475, x68619);
  nand n68476(x68476, x68474, x68475);
  nand n68477(x68477, x68475, x68471);
  nand n68479(x68479, x68480, x68620);
  nand n68481(x68481, x68479, x68480);
  nand n68482(x68482, x68480, x68475);
  nand n68484(x68484, x68485, x68621);
  nand n68486(x68486, x68484, x68485);
  nand n68487(x68487, x68485, x68480);
  nand n68489(x68489, x68472, x68471);
  nand n68490(x68490, x68478, x68618);
  nand n68492(x68492, x68490, x68491);
  nand n68493(x68493, x68483, x68619);
  nand n68495(x68495, x68493, x68494);
  nand n68496(x68496, x68483, x68473);
  nand n68497(x68497, x68488, x68476);
  nand n68499(x68499, x68497, x68498);
  nand n68500(x68500, x68488, x68478);
  nand n68503(x68503, x68496, x68502);
  nand n68504(x68504, x68501, x68618);
  nand n68506(x68506, x68504, x68505);
  nand n68507(x68507, x68619, x68470);
  nand n68508(x68508, x68507, x68472);
  nand n68510(x68510, x68475, x68489);
  nand n68512(x68512, x68620, x68511);
  nand n68513(x68513, x68512, x68510);
  nand n68515(x68515, x68480, x68492);
  nand n68517(x68517, x68621, x68516);
  nand n68518(x68518, x68517, x68515);
  nand n68520(x68520, x68485, x68503);
  nand n68522(x68522, x68622, x68521);
  nand n68523(x68523, x68522, x68520);
  nand n68525(x68525, x68530, x68506);
  nand n68527(x68527, x68623, x68526);
  nand n68528(x68528, x68527, x68525);
  nand n68531(x68531, x68619, x68618);
  nand n68532(x68532, x68620, x68619);
  nand n68534(x68534, x68621, x68620);
  nand n68536(x68536, x68622, x68621);
  nand n68538(x68538, x68533, x68618);
  nand n68539(x68539, x68535, x86398);
  nand n68540(x68540, x68537, x68533);
  nand n68542(x68542, x68541, x68618);
  nand n68543(x68543, x68471, x68470);
  nand n68544(x68544, x68543, x68531);
  nand n68546(x68546, x68620, x86398);
  nand n68547(x68547, x68475, x68531);
  nand n68548(x68548, x68547, x68546);
  nand n68550(x68550, x68621, x86399);
  nand n68551(x68551, x68480, x68538);
  nand n68552(x68552, x68551, x68550);
  nand n68554(x68554, x68622, x86400);
  nand n68555(x68555, x68485, x68539);
  nand n68556(x68556, x68555, x68554);
  nand n68558(x68558, x68623, x86401);
  nand n68559(x68559, x68530, x68542);
  nand n68560(x68560, x68559, x68558);
  nand n68562(x68562, x71128, x68618);
  nand n68564(x68564, x68563, x68470);
  nand n68565(x68565, x68564, x68562);
  nand n68566(x68566, x71128, x68470);
  nand n68567(x68567, x68563, x68618);
  nand n68568(x68568, x68567, x68566);
  nand n68569(x68569, x83382, x68565);
  nand n68571(x68571, x68570, x68568);
  nand n68572(x68572, x68571, x68569);
  nand n68573(x68573, x71128, x68619);
  nand n68574(x68574, x68563, x68545);
  nand n68575(x68575, x68574, x68573);
  nand n68576(x68576, x71128, x68509);
  nand n68577(x68577, x68563, x68619);
  nand n68578(x68578, x68577, x68576);
  nand n68579(x68579, x83382, x68575);
  nand n68580(x68580, x68570, x68578);
  nand n68581(x68581, x68580, x68579);
  nand n68582(x68582, x71128, x68620);
  nand n68583(x68583, x68563, x68549);
  nand n68584(x68584, x68583, x68582);
  nand n68585(x68585, x71128, x68514);
  nand n68586(x68586, x68563, x68620);
  nand n68587(x68587, x68586, x68585);
  nand n68588(x68588, x83382, x68584);
  nand n68589(x68589, x68570, x68587);
  nand n68590(x68590, x68589, x68588);
  nand n68591(x68591, x71128, x68621);
  nand n68592(x68592, x68563, x68553);
  nand n68593(x68593, x68592, x68591);
  nand n68594(x68594, x71128, x68519);
  nand n68595(x68595, x68563, x68621);
  nand n68596(x68596, x68595, x68594);
  nand n68597(x68597, x83382, x68593);
  nand n68598(x68598, x68570, x68596);
  nand n68599(x68599, x68598, x68597);
  nand n68600(x68600, x71128, x68622);
  nand n68601(x68601, x68563, x68557);
  nand n68602(x68602, x68601, x68600);
  nand n68603(x68603, x71128, x68524);
  nand n68604(x68604, x68563, x68622);
  nand n68605(x68605, x68604, x68603);
  nand n68606(x68606, x83382, x68602);
  nand n68607(x68607, x68570, x68605);
  nand n68608(x68608, x68607, x68606);
  nand n68609(x68609, x71128, x68623);
  nand n68610(x68610, x68563, x68561);
  nand n68611(x68611, x68610, x68609);
  nand n68612(x68612, x71128, x68529);
  nand n68613(x68613, x68563, x68623);
  nand n68614(x68614, x68613, x68612);
  nand n68615(x68615, x83382, x68611);
  nand n68616(x68616, x68570, x68614);
  nand n68617(x68617, x68616, x68615);
  nand n68630(x68630, x60784, x68624);
  nand n68631(x68631, x61367, x68625);
  nand n68632(x68632, x62873, x68626);
  nand n68633(x68633, x66413, x68627);
  nand n68634(x68634, x67405, x68628);
  nand n68635(x68635, x68398, x68629);
  nand n68636(x68636, x68634, x68635);
  nand n68637(x68637, x68632, x68633);
  nand n68638(x68638, x68630, x68631);
  nand n68642(x68642, x68641, x68640);
  nand n68644(x68644, x68643, x68639);
  nand n68645(x68645, x60784, x60824);
  nand n68646(x68646, x61367, x61407);
  nand n68647(x68647, x62873, x62913);
  nand n68648(x68648, x66413, x66453);
  nand n68649(x68649, x67405, x67445);
  nand n68650(x68650, x68398, x68438);
  nand n68651(x68651, x68649, x68650);
  nand n68652(x68652, x68647, x68648);
  nand n68653(x68653, x68645, x68646);
  nand n68657(x68657, x68656, x68655);
  nand n68659(x68659, x68658, x68654);
  nand n68664(x68664, x68639, x68660);
  nand n68665(x68665, x68639, x68661);
  nand n68666(x68666, x68639, x68662);
  nand n68667(x68667, x68636, x68663);
  nand n68668(x68668, x68639, x68663);
  nand n68669(x68669, x68668, x68667);
  nand n68670(x68670, x68665, x68666);
  nand n68672(x68672, x68671, x86402);
  nand n68673(x68673, x68670, x86403);
  nand n68674(x68674, x68671, x86403);
  nand n68675(x68675, x68674, x68673);
  nand n68676(x68676, x68671, x68669);
  nand n68678(x68678, x68672, x68677);
  nand n68680(x68680, x68679, x68676);
  nand n68685(x68685, x68654, x68681);
  nand n68686(x68686, x68654, x68682);
  nand n68687(x68687, x68654, x68683);
  nand n68688(x68688, x68651, x68684);
  nand n68689(x68689, x68654, x68684);
  nand n68690(x68690, x68689, x68688);
  nand n68691(x68691, x68686, x68687);
  nand n68693(x68693, x68692, x86404);
  nand n68694(x68694, x68691, x86405);
  nand n68695(x68695, x68692, x86405);
  nand n68696(x68696, x68695, x68694);
  nand n68697(x68697, x68692, x68690);
  nand n68699(x68699, x68693, x68698);
  nand n68701(x68701, x68700, x68697);
  nand n68704(x68704, x68671, x68745);
  nand n68705(x68705, x68671, x68680);
  nand n68706(x68706, x68670, x68745);
  nand n68707(x68707, x68670, x68680);
  nand n68708(x68708, x68639, x86406);
  nand n68709(x68709, x68639, x86407);
  nand n68710(x68710, x68639, x86408);
  nand n68711(x68711, x68639, x86409);
  nand n68712(x68712, x68636, x86406);
  nand n68713(x68713, x68636, x86407);
  nand n68714(x68714, x68708, x68702);
  nand n68715(x68715, x68709, x68660);
  nand n68716(x68716, x68710, x68661);
  nand n68717(x68717, x68711, x68662);
  nand n68718(x68718, x68712, x68703);
  nand n68719(x68719, x68713, x68663);
  nand n68722(x68722, x68692, x68810);
  nand n68723(x68723, x68692, x68701);
  nand n68724(x68724, x68691, x68810);
  nand n68725(x68725, x68691, x68701);
  nand n68726(x68726, x68654, x86410);
  nand n68727(x68727, x68654, x86411);
  nand n68728(x68728, x68654, x86412);
  nand n68729(x68729, x68654, x86413);
  nand n68730(x68730, x68651, x86410);
  nand n68731(x68731, x68651, x86411);
  nand n68732(x68732, x68726, x68720);
  nand n68733(x68733, x68727, x68681);
  nand n68734(x68734, x68728, x68682);
  nand n68735(x68735, x68729, x68683);
  nand n68736(x68736, x68730, x68721);
  nand n68737(x68737, x68731, x68684);
  nand n68738(x68738, x68714, x68732);
  nand n68739(x68739, x68715, x68733);
  nand n68740(x68740, x68716, x68734);
  nand n68741(x68741, x68717, x68735);
  nand n68742(x68742, x68718, x68736);
  nand n68743(x68743, x68719, x68737);
  nand n68744(x68744, x68680, x68442);
  nand n68746(x68746, x68745, x67449);
  nand n68747(x68747, x68746, x68744);
  nand n68748(x68748, x68680, x66457);
  nand n68749(x68749, x68745, x62917);
  nand n68750(x68750, x68749, x68748);
  nand n68751(x68751, x68680, x61411);
  nand n68752(x68752, x68745, x60828);
  nand n68753(x68753, x68752, x68751);
  nand n68754(x68754, x68671, x68747);
  nand n68755(x68755, x68670, x68750);
  nand n68756(x68756, x68671, x68753);
  nand n68757(x68757, x68756, x68755);
  nand n68758(x68758, x68636, x86414);
  nand n68759(x68759, x68639, x68757);
  nand n68760(x68760, x68759, x68758);
  nand n68761(x68761, x68680, x68446);
  nand n68762(x68762, x68745, x67453);
  nand n68763(x68763, x68762, x68761);
  nand n68764(x68764, x68680, x66461);
  nand n68765(x68765, x68745, x62921);
  nand n68766(x68766, x68765, x68764);
  nand n68767(x68767, x68680, x61415);
  nand n68768(x68768, x68745, x60832);
  nand n68769(x68769, x68768, x68767);
  nand n68770(x68770, x68671, x68763);
  nand n68771(x68771, x68670, x68766);
  nand n68772(x68772, x68671, x68769);
  nand n68773(x68773, x68772, x68771);
  nand n68774(x68774, x68636, x86415);
  nand n68775(x68775, x68639, x68773);
  nand n68776(x68776, x68775, x68774);
  nand n68777(x68777, x68680, x68450);
  nand n68778(x68778, x68745, x67457);
  nand n68779(x68779, x68778, x68777);
  nand n68780(x68780, x68680, x66465);
  nand n68781(x68781, x68745, x62925);
  nand n68782(x68782, x68781, x68780);
  nand n68783(x68783, x68680, x61419);
  nand n68784(x68784, x68745, x60836);
  nand n68785(x68785, x68784, x68783);
  nand n68786(x68786, x68671, x68779);
  nand n68787(x68787, x68670, x68782);
  nand n68788(x68788, x68671, x68785);
  nand n68789(x68789, x68788, x68787);
  nand n68790(x68790, x68636, x86416);
  nand n68791(x68791, x68639, x68789);
  nand n68792(x68792, x68791, x68790);
  nand n68793(x68793, x68680, x68454);
  nand n68794(x68794, x68745, x67461);
  nand n68795(x68795, x68794, x68793);
  nand n68796(x68796, x68680, x66469);
  nand n68797(x68797, x68745, x62929);
  nand n68798(x68798, x68797, x68796);
  nand n68799(x68799, x68680, x61423);
  nand n68800(x68800, x68745, x60840);
  nand n68801(x68801, x68800, x68799);
  nand n68802(x68802, x68671, x68795);
  nand n68803(x68803, x68670, x68798);
  nand n68804(x68804, x68671, x68801);
  nand n68805(x68805, x68804, x68803);
  nand n68806(x68806, x68636, x86417);
  nand n68807(x68807, x68639, x68805);
  nand n68808(x68808, x68807, x68806);
  nand n68809(x68809, x68701, x68442);
  nand n68811(x68811, x68810, x67449);
  nand n68812(x68812, x68811, x68809);
  nand n68813(x68813, x68701, x66457);
  nand n68814(x68814, x68810, x62917);
  nand n68815(x68815, x68814, x68813);
  nand n68816(x68816, x68701, x61411);
  nand n68817(x68817, x68810, x60828);
  nand n68818(x68818, x68817, x68816);
  nand n68819(x68819, x68692, x68812);
  nand n68820(x68820, x68691, x68815);
  nand n68821(x68821, x68692, x68818);
  nand n68822(x68822, x68821, x68820);
  nand n68823(x68823, x68651, x86418);
  nand n68824(x68824, x68654, x68822);
  nand n68825(x68825, x68824, x68823);
  nand n68826(x68826, x68701, x68446);
  nand n68827(x68827, x68810, x67453);
  nand n68828(x68828, x68827, x68826);
  nand n68829(x68829, x68701, x66461);
  nand n68830(x68830, x68810, x62921);
  nand n68831(x68831, x68830, x68829);
  nand n68832(x68832, x68701, x61415);
  nand n68833(x68833, x68810, x60832);
  nand n68834(x68834, x68833, x68832);
  nand n68835(x68835, x68692, x68828);
  nand n68836(x68836, x68691, x68831);
  nand n68837(x68837, x68692, x68834);
  nand n68838(x68838, x68837, x68836);
  nand n68839(x68839, x68651, x86419);
  nand n68840(x68840, x68654, x68838);
  nand n68841(x68841, x68840, x68839);
  nand n68842(x68842, x68701, x68450);
  nand n68843(x68843, x68810, x67457);
  nand n68844(x68844, x68843, x68842);
  nand n68845(x68845, x68701, x66465);
  nand n68846(x68846, x68810, x62925);
  nand n68847(x68847, x68846, x68845);
  nand n68848(x68848, x68701, x61419);
  nand n68849(x68849, x68810, x60836);
  nand n68850(x68850, x68849, x68848);
  nand n68851(x68851, x68692, x68844);
  nand n68852(x68852, x68691, x68847);
  nand n68853(x68853, x68692, x68850);
  nand n68854(x68854, x68853, x68852);
  nand n68855(x68855, x68651, x86420);
  nand n68856(x68856, x68654, x68854);
  nand n68857(x68857, x68856, x68855);
  nand n68858(x68858, x68701, x68454);
  nand n68859(x68859, x68810, x67461);
  nand n68860(x68860, x68859, x68858);
  nand n68861(x68861, x68701, x66469);
  nand n68862(x68862, x68810, x62929);
  nand n68863(x68863, x68862, x68861);
  nand n68864(x68864, x68701, x61423);
  nand n68865(x68865, x68810, x60840);
  nand n68866(x68866, x68865, x68864);
  nand n68867(x68867, x68692, x68860);
  nand n68868(x68868, x68691, x68863);
  nand n68869(x68869, x68692, x68866);
  nand n68870(x68870, x68869, x68868);
  nand n68871(x68871, x68651, x86421);
  nand n68872(x68872, x68654, x68870);
  nand n68873(x68873, x68872, x68871);
  nand n68874(x68874, x68680, x67887);
  nand n68875(x68875, x68745, x66894);
  nand n68876(x68876, x68875, x68874);
  nand n68877(x68877, x68680, x64274);
  nand n68878(x68878, x68745, x61981);
  nand n68879(x68879, x68878, x68877);
  nand n68880(x68880, x68680, x60976);
  nand n68881(x68881, x68745, x27755);
  nand n68882(x68882, x68881, x68880);
  nand n68883(x68883, x68671, x68876);
  nand n68884(x68884, x68670, x68879);
  nand n68885(x68885, x68671, x68882);
  nand n68886(x68886, x68885, x68884);
  nand n68887(x68887, x68636, x86422);
  nand n68888(x68888, x68639, x68886);
  nand n68889(x68889, x68888, x68887);
  nand n68890(x68890, x68680, x67891);
  nand n68891(x68891, x68745, x66898);
  nand n68892(x68892, x68891, x68890);
  nand n68893(x68893, x68680, x64277);
  nand n68894(x68894, x68745, x61988);
  nand n68895(x68895, x68894, x68893);
  nand n68896(x68896, x68745, x27759);
  nand n68897(x68897, x68671, x68892);
  nand n68898(x68898, x68670, x68895);
  nand n68899(x68899, x68671, x86423);
  nand n68900(x68900, x68899, x68898);
  nand n68901(x68901, x68636, x86424);
  nand n68902(x68902, x68639, x68900);
  nand n68903(x68903, x68902, x68901);
  nand n68904(x68904, x68680, x67895);
  nand n68905(x68905, x68745, x66902);
  nand n68906(x68906, x68905, x68904);
  nand n68907(x68907, x68680, x64280);
  nand n68908(x68908, x68745, x61995);
  nand n68909(x68909, x68908, x68907);
  nand n68910(x68910, x68745, x27763);
  nand n68911(x68911, x68671, x68906);
  nand n68912(x68912, x68670, x68909);
  nand n68913(x68913, x68671, x86425);
  nand n68914(x68914, x68913, x68912);
  nand n68915(x68915, x68636, x86426);
  nand n68916(x68916, x68639, x68914);
  nand n68917(x68917, x68916, x68915);
  nand n68918(x68918, x68680, x67899);
  nand n68919(x68919, x68745, x66906);
  nand n68920(x68920, x68919, x68918);
  nand n68921(x68921, x68680, x64283);
  nand n68922(x68922, x68745, x62002);
  nand n68923(x68923, x68922, x68921);
  nand n68924(x68924, x68745, x27767);
  nand n68925(x68925, x68671, x68920);
  nand n68926(x68926, x68670, x68923);
  nand n68927(x68927, x68671, x86427);
  nand n68928(x68928, x68927, x68926);
  nand n68929(x68929, x68636, x86428);
  nand n68930(x68930, x68639, x68928);
  nand n68931(x68931, x68930, x68929);
  nand n68932(x68932, x68680, x67903);
  nand n68933(x68933, x68745, x66910);
  nand n68934(x68934, x68933, x68932);
  nand n68935(x68935, x68680, x64286);
  nand n68936(x68936, x68745, x62009);
  nand n68937(x68937, x68936, x68935);
  nand n68938(x68938, x68745, x27771);
  nand n68939(x68939, x68671, x68934);
  nand n68940(x68940, x68670, x68937);
  nand n68941(x68941, x68671, x86429);
  nand n68942(x68942, x68941, x68940);
  nand n68943(x68943, x68636, x86430);
  nand n68944(x68944, x68639, x68942);
  nand n68945(x68945, x68944, x68943);
  nand n68946(x68946, x68680, x67907);
  nand n68947(x68947, x68745, x66914);
  nand n68948(x68948, x68947, x68946);
  nand n68949(x68949, x68680, x64289);
  nand n68950(x68950, x68745, x62016);
  nand n68951(x68951, x68950, x68949);
  nand n68952(x68952, x68745, x27775);
  nand n68953(x68953, x68671, x68948);
  nand n68954(x68954, x68670, x68951);
  nand n68955(x68955, x68671, x86431);
  nand n68956(x68956, x68955, x68954);
  nand n68957(x68957, x68636, x86432);
  nand n68958(x68958, x68639, x68956);
  nand n68959(x68959, x68958, x68957);
  nand n68960(x68960, x68680, x67911);
  nand n68961(x68961, x68745, x66918);
  nand n68962(x68962, x68961, x68960);
  nand n68963(x68963, x68680, x64292);
  nand n68964(x68964, x68745, x62023);
  nand n68965(x68965, x68964, x68963);
  nand n68966(x68966, x68745, x27779);
  nand n68967(x68967, x68671, x68962);
  nand n68968(x68968, x68670, x68965);
  nand n68969(x68969, x68671, x86433);
  nand n68970(x68970, x68969, x68968);
  nand n68971(x68971, x68636, x86434);
  nand n68972(x68972, x68639, x68970);
  nand n68973(x68973, x68972, x68971);
  nand n68974(x68974, x68680, x67915);
  nand n68975(x68975, x68745, x66922);
  nand n68976(x68976, x68975, x68974);
  nand n68977(x68977, x68680, x64295);
  nand n68978(x68978, x68745, x62030);
  nand n68979(x68979, x68978, x68977);
  nand n68980(x68980, x68745, x27783);
  nand n68981(x68981, x68671, x68976);
  nand n68982(x68982, x68670, x68979);
  nand n68983(x68983, x68671, x86435);
  nand n68984(x68984, x68983, x68982);
  nand n68985(x68985, x68636, x86436);
  nand n68986(x68986, x68639, x68984);
  nand n68987(x68987, x68986, x68985);
  nand n68988(x68988, x68680, x67919);
  nand n68989(x68989, x68745, x66926);
  nand n68990(x68990, x68989, x68988);
  nand n68991(x68991, x68680, x64298);
  nand n68992(x68992, x68745, x62037);
  nand n68993(x68993, x68992, x68991);
  nand n68994(x68994, x68745, x27787);
  nand n68995(x68995, x68671, x68990);
  nand n68996(x68996, x68670, x68993);
  nand n68997(x68997, x68671, x86437);
  nand n68998(x68998, x68997, x68996);
  nand n68999(x68999, x68636, x86438);
  nand n69000(x69000, x68639, x68998);
  nand n69001(x69001, x69000, x68999);
  nand n69002(x69002, x68680, x67923);
  nand n69003(x69003, x68745, x66930);
  nand n69004(x69004, x69003, x69002);
  nand n69005(x69005, x68680, x64301);
  nand n69006(x69006, x68745, x62044);
  nand n69007(x69007, x69006, x69005);
  nand n69008(x69008, x68745, x27791);
  nand n69009(x69009, x68671, x69004);
  nand n69010(x69010, x68670, x69007);
  nand n69011(x69011, x68671, x86439);
  nand n69012(x69012, x69011, x69010);
  nand n69013(x69013, x68636, x86440);
  nand n69014(x69014, x68639, x69012);
  nand n69015(x69015, x69014, x69013);
  nand n69016(x69016, x68680, x67927);
  nand n69017(x69017, x68745, x66934);
  nand n69018(x69018, x69017, x69016);
  nand n69019(x69019, x68680, x64304);
  nand n69020(x69020, x68745, x62051);
  nand n69021(x69021, x69020, x69019);
  nand n69022(x69022, x68745, x27795);
  nand n69023(x69023, x68671, x69018);
  nand n69024(x69024, x68670, x69021);
  nand n69025(x69025, x68671, x86441);
  nand n69026(x69026, x69025, x69024);
  nand n69027(x69027, x68636, x86442);
  nand n69028(x69028, x68639, x69026);
  nand n69029(x69029, x69028, x69027);
  nand n69030(x69030, x68680, x67931);
  nand n69031(x69031, x68745, x66938);
  nand n69032(x69032, x69031, x69030);
  nand n69033(x69033, x68680, x64307);
  nand n69034(x69034, x68745, x62058);
  nand n69035(x69035, x69034, x69033);
  nand n69036(x69036, x68745, x27799);
  nand n69037(x69037, x68671, x69032);
  nand n69038(x69038, x68670, x69035);
  nand n69039(x69039, x68671, x86443);
  nand n69040(x69040, x69039, x69038);
  nand n69041(x69041, x68636, x86444);
  nand n69042(x69042, x68639, x69040);
  nand n69043(x69043, x69042, x69041);
  nand n69044(x69044, x68680, x67935);
  nand n69045(x69045, x68745, x66942);
  nand n69046(x69046, x69045, x69044);
  nand n69047(x69047, x68680, x64310);
  nand n69048(x69048, x68745, x62065);
  nand n69049(x69049, x69048, x69047);
  nand n69050(x69050, x68745, x27803);
  nand n69051(x69051, x68671, x69046);
  nand n69052(x69052, x68670, x69049);
  nand n69053(x69053, x68671, x86445);
  nand n69054(x69054, x69053, x69052);
  nand n69055(x69055, x68636, x86446);
  nand n69056(x69056, x68639, x69054);
  nand n69057(x69057, x69056, x69055);
  nand n69058(x69058, x68680, x67939);
  nand n69059(x69059, x68745, x66946);
  nand n69060(x69060, x69059, x69058);
  nand n69061(x69061, x68680, x64313);
  nand n69062(x69062, x68745, x62072);
  nand n69063(x69063, x69062, x69061);
  nand n69064(x69064, x68745, x27807);
  nand n69065(x69065, x68671, x69060);
  nand n69066(x69066, x68670, x69063);
  nand n69067(x69067, x68671, x86447);
  nand n69068(x69068, x69067, x69066);
  nand n69069(x69069, x68636, x86448);
  nand n69070(x69070, x68639, x69068);
  nand n69071(x69071, x69070, x69069);
  nand n69072(x69072, x68680, x67943);
  nand n69073(x69073, x68745, x66950);
  nand n69074(x69074, x69073, x69072);
  nand n69075(x69075, x68680, x64316);
  nand n69076(x69076, x68745, x62079);
  nand n69077(x69077, x69076, x69075);
  nand n69078(x69078, x68745, x27811);
  nand n69079(x69079, x68671, x69074);
  nand n69080(x69080, x68670, x69077);
  nand n69081(x69081, x68671, x86449);
  nand n69082(x69082, x69081, x69080);
  nand n69083(x69083, x68636, x86450);
  nand n69084(x69084, x68639, x69082);
  nand n69085(x69085, x69084, x69083);
  nand n69086(x69086, x68680, x67947);
  nand n69087(x69087, x68745, x66954);
  nand n69088(x69088, x69087, x69086);
  nand n69089(x69089, x68680, x64319);
  nand n69090(x69090, x68745, x62086);
  nand n69091(x69091, x69090, x69089);
  nand n69092(x69092, x68745, x27815);
  nand n69093(x69093, x68671, x69088);
  nand n69094(x69094, x68670, x69091);
  nand n69095(x69095, x68671, x86451);
  nand n69096(x69096, x69095, x69094);
  nand n69097(x69097, x68636, x86452);
  nand n69098(x69098, x68639, x69096);
  nand n69099(x69099, x69098, x69097);
  nand n69100(x69100, x68680, x67951);
  nand n69101(x69101, x68745, x66958);
  nand n69102(x69102, x69101, x69100);
  nand n69103(x69103, x68680, x86281);
  nand n69104(x69104, x68745, x62093);
  nand n69105(x69105, x69104, x69103);
  nand n69106(x69106, x68745, x27819);
  nand n69107(x69107, x68671, x69102);
  nand n69108(x69108, x68670, x69105);
  nand n69109(x69109, x68671, x86453);
  nand n69110(x69110, x69109, x69108);
  nand n69111(x69111, x68636, x86454);
  nand n69112(x69112, x68639, x69110);
  nand n69113(x69113, x69112, x69111);
  nand n69114(x69114, x68680, x67955);
  nand n69115(x69115, x68745, x66962);
  nand n69116(x69116, x69115, x69114);
  nand n69117(x69117, x68680, x86282);
  nand n69118(x69118, x68745, x62100);
  nand n69119(x69119, x69118, x69117);
  nand n69120(x69120, x68745, x27823);
  nand n69121(x69121, x68671, x69116);
  nand n69122(x69122, x68670, x69119);
  nand n69123(x69123, x68671, x86455);
  nand n69124(x69124, x69123, x69122);
  nand n69125(x69125, x68636, x86456);
  nand n69126(x69126, x68639, x69124);
  nand n69127(x69127, x69126, x69125);
  nand n69128(x69128, x68680, x67959);
  nand n69129(x69129, x68745, x66966);
  nand n69130(x69130, x69129, x69128);
  nand n69131(x69131, x68680, x86283);
  nand n69132(x69132, x68745, x62107);
  nand n69133(x69133, x69132, x69131);
  nand n69134(x69134, x68745, x27827);
  nand n69135(x69135, x68671, x69130);
  nand n69136(x69136, x68670, x69133);
  nand n69137(x69137, x68671, x86457);
  nand n69138(x69138, x69137, x69136);
  nand n69139(x69139, x68636, x86458);
  nand n69140(x69140, x68639, x69138);
  nand n69141(x69141, x69140, x69139);
  nand n69142(x69142, x68680, x67963);
  nand n69143(x69143, x68745, x66970);
  nand n69144(x69144, x69143, x69142);
  nand n69145(x69145, x68680, x86284);
  nand n69146(x69146, x68745, x62114);
  nand n69147(x69147, x69146, x69145);
  nand n69148(x69148, x68745, x27831);
  nand n69149(x69149, x68671, x69144);
  nand n69150(x69150, x68670, x69147);
  nand n69151(x69151, x68671, x86459);
  nand n69152(x69152, x69151, x69150);
  nand n69153(x69153, x68636, x86460);
  nand n69154(x69154, x68639, x69152);
  nand n69155(x69155, x69154, x69153);
  nand n69156(x69156, x68680, x67967);
  nand n69157(x69157, x68745, x66974);
  nand n69158(x69158, x69157, x69156);
  nand n69159(x69159, x68680, x86285);
  nand n69160(x69160, x68745, x62121);
  nand n69161(x69161, x69160, x69159);
  nand n69162(x69162, x68745, x27835);
  nand n69163(x69163, x68671, x69158);
  nand n69164(x69164, x68670, x69161);
  nand n69165(x69165, x68671, x86461);
  nand n69166(x69166, x69165, x69164);
  nand n69167(x69167, x68636, x86462);
  nand n69168(x69168, x68639, x69166);
  nand n69169(x69169, x69168, x69167);
  nand n69170(x69170, x68680, x67971);
  nand n69171(x69171, x68745, x66978);
  nand n69172(x69172, x69171, x69170);
  nand n69173(x69173, x68680, x86286);
  nand n69174(x69174, x68745, x62128);
  nand n69175(x69175, x69174, x69173);
  nand n69176(x69176, x68745, x27839);
  nand n69177(x69177, x68671, x69172);
  nand n69178(x69178, x68670, x69175);
  nand n69179(x69179, x68671, x86463);
  nand n69180(x69180, x69179, x69178);
  nand n69181(x69181, x68636, x86464);
  nand n69182(x69182, x68639, x69180);
  nand n69183(x69183, x69182, x69181);
  nand n69184(x69184, x68680, x67975);
  nand n69185(x69185, x68745, x66982);
  nand n69186(x69186, x69185, x69184);
  nand n69187(x69187, x68680, x86287);
  nand n69188(x69188, x68745, x62135);
  nand n69189(x69189, x69188, x69187);
  nand n69190(x69190, x68745, x27843);
  nand n69191(x69191, x68671, x69186);
  nand n69192(x69192, x68670, x69189);
  nand n69193(x69193, x68671, x86465);
  nand n69194(x69194, x69193, x69192);
  nand n69195(x69195, x68636, x86466);
  nand n69196(x69196, x68639, x69194);
  nand n69197(x69197, x69196, x69195);
  nand n69198(x69198, x68680, x67979);
  nand n69199(x69199, x68745, x66986);
  nand n69200(x69200, x69199, x69198);
  nand n69201(x69201, x68680, x86288);
  nand n69202(x69202, x68745, x62142);
  nand n69203(x69203, x69202, x69201);
  nand n69204(x69204, x68745, x27847);
  nand n69205(x69205, x68671, x69200);
  nand n69206(x69206, x68670, x69203);
  nand n69207(x69207, x68671, x86467);
  nand n69208(x69208, x69207, x69206);
  nand n69209(x69209, x68636, x86468);
  nand n69210(x69210, x68639, x69208);
  nand n69211(x69211, x69210, x69209);
  nand n69212(x69212, x68680, x67983);
  nand n69213(x69213, x68745, x66990);
  nand n69214(x69214, x69213, x69212);
  nand n69215(x69215, x68680, x86289);
  nand n69216(x69216, x68745, x62149);
  nand n69217(x69217, x69216, x69215);
  nand n69218(x69218, x68745, x27851);
  nand n69219(x69219, x68671, x69214);
  nand n69220(x69220, x68670, x69217);
  nand n69221(x69221, x68671, x86469);
  nand n69222(x69222, x69221, x69220);
  nand n69223(x69223, x68636, x86470);
  nand n69224(x69224, x68639, x69222);
  nand n69225(x69225, x69224, x69223);
  nand n69226(x69226, x68680, x67987);
  nand n69227(x69227, x68745, x66994);
  nand n69228(x69228, x69227, x69226);
  nand n69229(x69229, x68680, x86290);
  nand n69230(x69230, x68745, x62156);
  nand n69231(x69231, x69230, x69229);
  nand n69232(x69232, x68745, x27855);
  nand n69233(x69233, x68671, x69228);
  nand n69234(x69234, x68670, x69231);
  nand n69235(x69235, x68671, x86471);
  nand n69236(x69236, x69235, x69234);
  nand n69237(x69237, x68636, x86472);
  nand n69238(x69238, x68639, x69236);
  nand n69239(x69239, x69238, x69237);
  nand n69240(x69240, x68680, x67991);
  nand n69241(x69241, x68745, x66998);
  nand n69242(x69242, x69241, x69240);
  nand n69243(x69243, x68680, x86291);
  nand n69244(x69244, x68745, x62163);
  nand n69245(x69245, x69244, x69243);
  nand n69246(x69246, x68745, x27859);
  nand n69247(x69247, x68671, x69242);
  nand n69248(x69248, x68670, x69245);
  nand n69249(x69249, x68671, x86473);
  nand n69250(x69250, x69249, x69248);
  nand n69251(x69251, x68636, x86474);
  nand n69252(x69252, x68639, x69250);
  nand n69253(x69253, x69252, x69251);
  nand n69254(x69254, x68680, x67995);
  nand n69255(x69255, x68745, x67002);
  nand n69256(x69256, x69255, x69254);
  nand n69257(x69257, x68680, x86292);
  nand n69258(x69258, x68745, x62170);
  nand n69259(x69259, x69258, x69257);
  nand n69260(x69260, x68745, x27863);
  nand n69261(x69261, x68671, x69256);
  nand n69262(x69262, x68670, x69259);
  nand n69263(x69263, x68671, x86475);
  nand n69264(x69264, x69263, x69262);
  nand n69265(x69265, x68636, x86476);
  nand n69266(x69266, x68639, x69264);
  nand n69267(x69267, x69266, x69265);
  nand n69268(x69268, x68680, x67999);
  nand n69269(x69269, x68745, x67006);
  nand n69270(x69270, x69269, x69268);
  nand n69271(x69271, x68680, x86293);
  nand n69272(x69272, x68745, x62177);
  nand n69273(x69273, x69272, x69271);
  nand n69274(x69274, x68745, x27867);
  nand n69275(x69275, x68671, x69270);
  nand n69276(x69276, x68670, x69273);
  nand n69277(x69277, x68671, x86477);
  nand n69278(x69278, x69277, x69276);
  nand n69279(x69279, x68636, x86478);
  nand n69280(x69280, x68639, x69278);
  nand n69281(x69281, x69280, x69279);
  nand n69282(x69282, x68680, x68003);
  nand n69283(x69283, x68745, x67010);
  nand n69284(x69284, x69283, x69282);
  nand n69285(x69285, x68680, x86294);
  nand n69286(x69286, x68745, x62184);
  nand n69287(x69287, x69286, x69285);
  nand n69288(x69288, x68745, x27871);
  nand n69289(x69289, x68671, x69284);
  nand n69290(x69290, x68670, x69287);
  nand n69291(x69291, x68671, x86479);
  nand n69292(x69292, x69291, x69290);
  nand n69293(x69293, x68636, x86480);
  nand n69294(x69294, x68639, x69292);
  nand n69295(x69295, x69294, x69293);
  nand n69296(x69296, x68680, x68007);
  nand n69297(x69297, x68745, x67014);
  nand n69298(x69298, x69297, x69296);
  nand n69299(x69299, x68680, x86295);
  nand n69300(x69300, x68745, x62191);
  nand n69301(x69301, x69300, x69299);
  nand n69302(x69302, x68745, x27875);
  nand n69303(x69303, x68671, x69298);
  nand n69304(x69304, x68670, x69301);
  nand n69305(x69305, x68671, x86481);
  nand n69306(x69306, x69305, x69304);
  nand n69307(x69307, x68636, x86482);
  nand n69308(x69308, x68639, x69306);
  nand n69309(x69309, x69308, x69307);
  nand n69310(x69310, x68680, x68011);
  nand n69311(x69311, x68745, x67018);
  nand n69312(x69312, x69311, x69310);
  nand n69313(x69313, x68680, x86296);
  nand n69314(x69314, x68745, x62198);
  nand n69315(x69315, x69314, x69313);
  nand n69316(x69316, x68745, x27879);
  nand n69317(x69317, x68671, x69312);
  nand n69318(x69318, x68670, x69315);
  nand n69319(x69319, x68671, x86483);
  nand n69320(x69320, x69319, x69318);
  nand n69321(x69321, x68636, x86484);
  nand n69322(x69322, x68639, x69320);
  nand n69323(x69323, x69322, x69321);
  nand n69324(x69324, x68680, x68015);
  nand n69325(x69325, x68745, x67022);
  nand n69326(x69326, x69325, x69324);
  nand n69327(x69327, x68680, x65006);
  nand n69328(x69328, x68745, x62205);
  nand n69329(x69329, x69328, x69327);
  nand n69330(x69330, x68680, x61105);
  nand n69331(x69331, x68745, x38722);
  nand n69332(x69332, x69331, x69330);
  nand n69333(x69333, x68671, x69326);
  nand n69334(x69334, x68670, x69329);
  nand n69335(x69335, x68671, x69332);
  nand n69336(x69336, x69335, x69334);
  nand n69337(x69337, x68636, x86485);
  nand n69338(x69338, x68639, x69336);
  nand n69339(x69339, x69338, x69337);
  nand n69340(x69340, x68680, x68019);
  nand n69341(x69341, x68745, x67026);
  nand n69342(x69342, x69341, x69340);
  nand n69343(x69343, x68680, x65009);
  nand n69344(x69344, x68745, x62212);
  nand n69345(x69345, x69344, x69343);
  nand n69346(x69346, x68745, x38726);
  nand n69347(x69347, x68671, x69342);
  nand n69348(x69348, x68670, x69345);
  nand n69349(x69349, x68671, x86486);
  nand n69350(x69350, x69349, x69348);
  nand n69351(x69351, x68636, x86487);
  nand n69352(x69352, x68639, x69350);
  nand n69353(x69353, x69352, x69351);
  nand n69354(x69354, x68680, x68023);
  nand n69355(x69355, x68745, x67030);
  nand n69356(x69356, x69355, x69354);
  nand n69357(x69357, x68680, x65012);
  nand n69358(x69358, x68745, x62219);
  nand n69359(x69359, x69358, x69357);
  nand n69360(x69360, x68745, x38730);
  nand n69361(x69361, x68671, x69356);
  nand n69362(x69362, x68670, x69359);
  nand n69363(x69363, x68671, x86488);
  nand n69364(x69364, x69363, x69362);
  nand n69365(x69365, x68636, x86489);
  nand n69366(x69366, x68639, x69364);
  nand n69367(x69367, x69366, x69365);
  nand n69368(x69368, x68680, x68027);
  nand n69369(x69369, x68745, x67034);
  nand n69370(x69370, x69369, x69368);
  nand n69371(x69371, x68680, x65015);
  nand n69372(x69372, x68745, x62226);
  nand n69373(x69373, x69372, x69371);
  nand n69374(x69374, x68745, x38734);
  nand n69375(x69375, x68671, x69370);
  nand n69376(x69376, x68670, x69373);
  nand n69377(x69377, x68671, x86490);
  nand n69378(x69378, x69377, x69376);
  nand n69379(x69379, x68636, x86491);
  nand n69380(x69380, x68639, x69378);
  nand n69381(x69381, x69380, x69379);
  nand n69382(x69382, x68680, x68031);
  nand n69383(x69383, x68745, x67038);
  nand n69384(x69384, x69383, x69382);
  nand n69385(x69385, x68680, x65018);
  nand n69386(x69386, x68745, x62233);
  nand n69387(x69387, x69386, x69385);
  nand n69388(x69388, x68745, x38738);
  nand n69389(x69389, x68671, x69384);
  nand n69390(x69390, x68670, x69387);
  nand n69391(x69391, x68671, x86492);
  nand n69392(x69392, x69391, x69390);
  nand n69393(x69393, x68636, x86493);
  nand n69394(x69394, x68639, x69392);
  nand n69395(x69395, x69394, x69393);
  nand n69396(x69396, x68680, x68035);
  nand n69397(x69397, x68745, x67042);
  nand n69398(x69398, x69397, x69396);
  nand n69399(x69399, x68680, x65021);
  nand n69400(x69400, x68745, x62240);
  nand n69401(x69401, x69400, x69399);
  nand n69402(x69402, x68745, x38742);
  nand n69403(x69403, x68671, x69398);
  nand n69404(x69404, x68670, x69401);
  nand n69405(x69405, x68671, x86494);
  nand n69406(x69406, x69405, x69404);
  nand n69407(x69407, x68636, x86495);
  nand n69408(x69408, x68639, x69406);
  nand n69409(x69409, x69408, x69407);
  nand n69410(x69410, x68680, x68039);
  nand n69411(x69411, x68745, x67046);
  nand n69412(x69412, x69411, x69410);
  nand n69413(x69413, x68680, x65024);
  nand n69414(x69414, x68745, x62247);
  nand n69415(x69415, x69414, x69413);
  nand n69416(x69416, x68745, x38746);
  nand n69417(x69417, x68671, x69412);
  nand n69418(x69418, x68670, x69415);
  nand n69419(x69419, x68671, x86496);
  nand n69420(x69420, x69419, x69418);
  nand n69421(x69421, x68636, x86497);
  nand n69422(x69422, x68639, x69420);
  nand n69423(x69423, x69422, x69421);
  nand n69424(x69424, x68680, x68043);
  nand n69425(x69425, x68745, x67050);
  nand n69426(x69426, x69425, x69424);
  nand n69427(x69427, x68680, x65027);
  nand n69428(x69428, x68745, x62254);
  nand n69429(x69429, x69428, x69427);
  nand n69430(x69430, x68745, x38750);
  nand n69431(x69431, x68671, x69426);
  nand n69432(x69432, x68670, x69429);
  nand n69433(x69433, x68671, x86498);
  nand n69434(x69434, x69433, x69432);
  nand n69435(x69435, x68636, x86499);
  nand n69436(x69436, x68639, x69434);
  nand n69437(x69437, x69436, x69435);
  nand n69438(x69438, x68680, x68047);
  nand n69439(x69439, x68745, x67054);
  nand n69440(x69440, x69439, x69438);
  nand n69441(x69441, x68680, x65030);
  nand n69442(x69442, x68745, x62261);
  nand n69443(x69443, x69442, x69441);
  nand n69444(x69444, x68745, x38754);
  nand n69445(x69445, x68671, x69440);
  nand n69446(x69446, x68670, x69443);
  nand n69447(x69447, x68671, x86500);
  nand n69448(x69448, x69447, x69446);
  nand n69449(x69449, x68636, x86501);
  nand n69450(x69450, x68639, x69448);
  nand n69451(x69451, x69450, x69449);
  nand n69452(x69452, x68680, x68051);
  nand n69453(x69453, x68745, x67058);
  nand n69454(x69454, x69453, x69452);
  nand n69455(x69455, x68680, x65033);
  nand n69456(x69456, x68745, x62268);
  nand n69457(x69457, x69456, x69455);
  nand n69458(x69458, x68745, x38758);
  nand n69459(x69459, x68671, x69454);
  nand n69460(x69460, x68670, x69457);
  nand n69461(x69461, x68671, x86502);
  nand n69462(x69462, x69461, x69460);
  nand n69463(x69463, x68636, x86503);
  nand n69464(x69464, x68639, x69462);
  nand n69465(x69465, x69464, x69463);
  nand n69466(x69466, x68680, x68055);
  nand n69467(x69467, x68745, x67062);
  nand n69468(x69468, x69467, x69466);
  nand n69469(x69469, x68680, x65036);
  nand n69470(x69470, x68745, x62275);
  nand n69471(x69471, x69470, x69469);
  nand n69472(x69472, x68745, x38762);
  nand n69473(x69473, x68671, x69468);
  nand n69474(x69474, x68670, x69471);
  nand n69475(x69475, x68671, x86504);
  nand n69476(x69476, x69475, x69474);
  nand n69477(x69477, x68636, x86505);
  nand n69478(x69478, x68639, x69476);
  nand n69479(x69479, x69478, x69477);
  nand n69480(x69480, x68680, x68059);
  nand n69481(x69481, x68745, x67066);
  nand n69482(x69482, x69481, x69480);
  nand n69483(x69483, x68680, x65039);
  nand n69484(x69484, x68745, x62282);
  nand n69485(x69485, x69484, x69483);
  nand n69486(x69486, x68745, x38766);
  nand n69487(x69487, x68671, x69482);
  nand n69488(x69488, x68670, x69485);
  nand n69489(x69489, x68671, x86506);
  nand n69490(x69490, x69489, x69488);
  nand n69491(x69491, x68636, x86507);
  nand n69492(x69492, x68639, x69490);
  nand n69493(x69493, x69492, x69491);
  nand n69494(x69494, x68680, x68063);
  nand n69495(x69495, x68745, x67070);
  nand n69496(x69496, x69495, x69494);
  nand n69497(x69497, x68680, x65042);
  nand n69498(x69498, x68745, x62289);
  nand n69499(x69499, x69498, x69497);
  nand n69500(x69500, x68745, x38770);
  nand n69501(x69501, x68671, x69496);
  nand n69502(x69502, x68670, x69499);
  nand n69503(x69503, x68671, x86508);
  nand n69504(x69504, x69503, x69502);
  nand n69505(x69505, x68636, x86509);
  nand n69506(x69506, x68639, x69504);
  nand n69507(x69507, x69506, x69505);
  nand n69508(x69508, x68680, x68067);
  nand n69509(x69509, x68745, x67074);
  nand n69510(x69510, x69509, x69508);
  nand n69511(x69511, x68680, x65045);
  nand n69512(x69512, x68745, x62296);
  nand n69513(x69513, x69512, x69511);
  nand n69514(x69514, x68745, x38774);
  nand n69515(x69515, x68671, x69510);
  nand n69516(x69516, x68670, x69513);
  nand n69517(x69517, x68671, x86510);
  nand n69518(x69518, x69517, x69516);
  nand n69519(x69519, x68636, x86511);
  nand n69520(x69520, x68639, x69518);
  nand n69521(x69521, x69520, x69519);
  nand n69522(x69522, x68680, x68071);
  nand n69523(x69523, x68745, x67078);
  nand n69524(x69524, x69523, x69522);
  nand n69525(x69525, x68680, x65048);
  nand n69526(x69526, x68745, x62303);
  nand n69527(x69527, x69526, x69525);
  nand n69528(x69528, x68745, x38778);
  nand n69529(x69529, x68671, x69524);
  nand n69530(x69530, x68670, x69527);
  nand n69531(x69531, x68671, x86512);
  nand n69532(x69532, x69531, x69530);
  nand n69533(x69533, x68636, x86513);
  nand n69534(x69534, x68639, x69532);
  nand n69535(x69535, x69534, x69533);
  nand n69536(x69536, x68680, x68075);
  nand n69537(x69537, x68745, x67082);
  nand n69538(x69538, x69537, x69536);
  nand n69539(x69539, x68680, x65051);
  nand n69540(x69540, x68745, x62310);
  nand n69541(x69541, x69540, x69539);
  nand n69542(x69542, x68745, x38782);
  nand n69543(x69543, x68671, x69538);
  nand n69544(x69544, x68670, x69541);
  nand n69545(x69545, x68671, x86514);
  nand n69546(x69546, x69545, x69544);
  nand n69547(x69547, x68636, x86515);
  nand n69548(x69548, x68639, x69546);
  nand n69549(x69549, x69548, x69547);
  nand n69550(x69550, x68680, x68079);
  nand n69551(x69551, x68745, x67086);
  nand n69552(x69552, x69551, x69550);
  nand n69553(x69553, x68680, x86314);
  nand n69554(x69554, x68745, x62317);
  nand n69555(x69555, x69554, x69553);
  nand n69556(x69556, x68745, x38786);
  nand n69557(x69557, x68671, x69552);
  nand n69558(x69558, x68670, x69555);
  nand n69559(x69559, x68671, x86516);
  nand n69560(x69560, x69559, x69558);
  nand n69561(x69561, x68636, x86517);
  nand n69562(x69562, x68639, x69560);
  nand n69563(x69563, x69562, x69561);
  nand n69564(x69564, x68680, x68083);
  nand n69565(x69565, x68745, x67090);
  nand n69566(x69566, x69565, x69564);
  nand n69567(x69567, x68680, x86315);
  nand n69568(x69568, x68745, x62324);
  nand n69569(x69569, x69568, x69567);
  nand n69570(x69570, x68745, x38790);
  nand n69571(x69571, x68671, x69566);
  nand n69572(x69572, x68670, x69569);
  nand n69573(x69573, x68671, x86518);
  nand n69574(x69574, x69573, x69572);
  nand n69575(x69575, x68636, x86519);
  nand n69576(x69576, x68639, x69574);
  nand n69577(x69577, x69576, x69575);
  nand n69578(x69578, x68680, x68087);
  nand n69579(x69579, x68745, x67094);
  nand n69580(x69580, x69579, x69578);
  nand n69581(x69581, x68680, x86316);
  nand n69582(x69582, x68745, x62331);
  nand n69583(x69583, x69582, x69581);
  nand n69584(x69584, x68745, x38794);
  nand n69585(x69585, x68671, x69580);
  nand n69586(x69586, x68670, x69583);
  nand n69587(x69587, x68671, x86520);
  nand n69588(x69588, x69587, x69586);
  nand n69589(x69589, x68636, x86521);
  nand n69590(x69590, x68639, x69588);
  nand n69591(x69591, x69590, x69589);
  nand n69592(x69592, x68680, x68091);
  nand n69593(x69593, x68745, x67098);
  nand n69594(x69594, x69593, x69592);
  nand n69595(x69595, x68680, x86317);
  nand n69596(x69596, x68745, x62338);
  nand n69597(x69597, x69596, x69595);
  nand n69598(x69598, x68745, x38798);
  nand n69599(x69599, x68671, x69594);
  nand n69600(x69600, x68670, x69597);
  nand n69601(x69601, x68671, x86522);
  nand n69602(x69602, x69601, x69600);
  nand n69603(x69603, x68636, x86523);
  nand n69604(x69604, x68639, x69602);
  nand n69605(x69605, x69604, x69603);
  nand n69606(x69606, x68680, x68095);
  nand n69607(x69607, x68745, x67102);
  nand n69608(x69608, x69607, x69606);
  nand n69609(x69609, x68680, x86318);
  nand n69610(x69610, x68745, x62345);
  nand n69611(x69611, x69610, x69609);
  nand n69612(x69612, x68745, x38802);
  nand n69613(x69613, x68671, x69608);
  nand n69614(x69614, x68670, x69611);
  nand n69615(x69615, x68671, x86524);
  nand n69616(x69616, x69615, x69614);
  nand n69617(x69617, x68636, x86525);
  nand n69618(x69618, x68639, x69616);
  nand n69619(x69619, x69618, x69617);
  nand n69620(x69620, x68680, x68099);
  nand n69621(x69621, x68745, x67106);
  nand n69622(x69622, x69621, x69620);
  nand n69623(x69623, x68680, x86319);
  nand n69624(x69624, x68745, x62352);
  nand n69625(x69625, x69624, x69623);
  nand n69626(x69626, x68745, x38806);
  nand n69627(x69627, x68671, x69622);
  nand n69628(x69628, x68670, x69625);
  nand n69629(x69629, x68671, x86526);
  nand n69630(x69630, x69629, x69628);
  nand n69631(x69631, x68636, x86527);
  nand n69632(x69632, x68639, x69630);
  nand n69633(x69633, x69632, x69631);
  nand n69634(x69634, x68680, x68103);
  nand n69635(x69635, x68745, x67110);
  nand n69636(x69636, x69635, x69634);
  nand n69637(x69637, x68680, x86320);
  nand n69638(x69638, x68745, x62359);
  nand n69639(x69639, x69638, x69637);
  nand n69640(x69640, x68745, x38810);
  nand n69641(x69641, x68671, x69636);
  nand n69642(x69642, x68670, x69639);
  nand n69643(x69643, x68671, x86528);
  nand n69644(x69644, x69643, x69642);
  nand n69645(x69645, x68636, x86529);
  nand n69646(x69646, x68639, x69644);
  nand n69647(x69647, x69646, x69645);
  nand n69648(x69648, x68680, x68107);
  nand n69649(x69649, x68745, x67114);
  nand n69650(x69650, x69649, x69648);
  nand n69651(x69651, x68680, x86321);
  nand n69652(x69652, x68745, x62366);
  nand n69653(x69653, x69652, x69651);
  nand n69654(x69654, x68745, x38814);
  nand n69655(x69655, x68671, x69650);
  nand n69656(x69656, x68670, x69653);
  nand n69657(x69657, x68671, x86530);
  nand n69658(x69658, x69657, x69656);
  nand n69659(x69659, x68636, x86531);
  nand n69660(x69660, x68639, x69658);
  nand n69661(x69661, x69660, x69659);
  nand n69662(x69662, x68680, x68111);
  nand n69663(x69663, x68745, x67118);
  nand n69664(x69664, x69663, x69662);
  nand n69665(x69665, x68680, x86322);
  nand n69666(x69666, x68745, x62373);
  nand n69667(x69667, x69666, x69665);
  nand n69668(x69668, x68745, x38818);
  nand n69669(x69669, x68671, x69664);
  nand n69670(x69670, x68670, x69667);
  nand n69671(x69671, x68671, x86532);
  nand n69672(x69672, x69671, x69670);
  nand n69673(x69673, x68636, x86533);
  nand n69674(x69674, x68639, x69672);
  nand n69675(x69675, x69674, x69673);
  nand n69676(x69676, x68680, x68115);
  nand n69677(x69677, x68745, x67122);
  nand n69678(x69678, x69677, x69676);
  nand n69679(x69679, x68680, x86323);
  nand n69680(x69680, x68745, x62380);
  nand n69681(x69681, x69680, x69679);
  nand n69682(x69682, x68745, x38822);
  nand n69683(x69683, x68671, x69678);
  nand n69684(x69684, x68670, x69681);
  nand n69685(x69685, x68671, x86534);
  nand n69686(x69686, x69685, x69684);
  nand n69687(x69687, x68636, x86535);
  nand n69688(x69688, x68639, x69686);
  nand n69689(x69689, x69688, x69687);
  nand n69690(x69690, x68680, x68119);
  nand n69691(x69691, x68745, x67126);
  nand n69692(x69692, x69691, x69690);
  nand n69693(x69693, x68680, x86324);
  nand n69694(x69694, x68745, x62387);
  nand n69695(x69695, x69694, x69693);
  nand n69696(x69696, x68745, x38826);
  nand n69697(x69697, x68671, x69692);
  nand n69698(x69698, x68670, x69695);
  nand n69699(x69699, x68671, x86536);
  nand n69700(x69700, x69699, x69698);
  nand n69701(x69701, x68636, x86537);
  nand n69702(x69702, x68639, x69700);
  nand n69703(x69703, x69702, x69701);
  nand n69704(x69704, x68680, x68123);
  nand n69705(x69705, x68745, x67130);
  nand n69706(x69706, x69705, x69704);
  nand n69707(x69707, x68680, x86325);
  nand n69708(x69708, x68745, x62394);
  nand n69709(x69709, x69708, x69707);
  nand n69710(x69710, x68745, x38830);
  nand n69711(x69711, x68671, x69706);
  nand n69712(x69712, x68670, x69709);
  nand n69713(x69713, x68671, x86538);
  nand n69714(x69714, x69713, x69712);
  nand n69715(x69715, x68636, x86539);
  nand n69716(x69716, x68639, x69714);
  nand n69717(x69717, x69716, x69715);
  nand n69718(x69718, x68680, x68127);
  nand n69719(x69719, x68745, x67134);
  nand n69720(x69720, x69719, x69718);
  nand n69721(x69721, x68680, x86326);
  nand n69722(x69722, x68745, x62401);
  nand n69723(x69723, x69722, x69721);
  nand n69724(x69724, x68745, x38834);
  nand n69725(x69725, x68671, x69720);
  nand n69726(x69726, x68670, x69723);
  nand n69727(x69727, x68671, x86540);
  nand n69728(x69728, x69727, x69726);
  nand n69729(x69729, x68636, x86541);
  nand n69730(x69730, x68639, x69728);
  nand n69731(x69731, x69730, x69729);
  nand n69732(x69732, x68680, x68131);
  nand n69733(x69733, x68745, x67138);
  nand n69734(x69734, x69733, x69732);
  nand n69735(x69735, x68680, x86327);
  nand n69736(x69736, x68745, x62408);
  nand n69737(x69737, x69736, x69735);
  nand n69738(x69738, x68745, x38838);
  nand n69739(x69739, x68671, x69734);
  nand n69740(x69740, x68670, x69737);
  nand n69741(x69741, x68671, x86542);
  nand n69742(x69742, x69741, x69740);
  nand n69743(x69743, x68636, x86543);
  nand n69744(x69744, x68639, x69742);
  nand n69745(x69745, x69744, x69743);
  nand n69746(x69746, x68680, x68135);
  nand n69747(x69747, x68745, x67142);
  nand n69748(x69748, x69747, x69746);
  nand n69749(x69749, x68680, x86328);
  nand n69750(x69750, x68745, x62415);
  nand n69751(x69751, x69750, x69749);
  nand n69752(x69752, x68745, x38842);
  nand n69753(x69753, x68671, x69748);
  nand n69754(x69754, x68670, x69751);
  nand n69755(x69755, x68671, x86544);
  nand n69756(x69756, x69755, x69754);
  nand n69757(x69757, x68636, x86545);
  nand n69758(x69758, x68639, x69756);
  nand n69759(x69759, x69758, x69757);
  nand n69760(x69760, x68680, x68139);
  nand n69761(x69761, x68745, x67146);
  nand n69762(x69762, x69761, x69760);
  nand n69763(x69763, x68680, x86329);
  nand n69764(x69764, x68745, x62422);
  nand n69765(x69765, x69764, x69763);
  nand n69766(x69766, x68745, x38846);
  nand n69767(x69767, x68671, x69762);
  nand n69768(x69768, x68670, x69765);
  nand n69769(x69769, x68671, x86546);
  nand n69770(x69770, x69769, x69768);
  nand n69771(x69771, x68636, x86547);
  nand n69772(x69772, x68639, x69770);
  nand n69773(x69773, x69772, x69771);
  nand n69774(x69774, x68680, x68143);
  nand n69775(x69775, x68745, x67150);
  nand n69776(x69776, x69775, x69774);
  nand n69777(x69777, x68680, x65676);
  nand n69778(x69778, x68745, x62429);
  nand n69779(x69779, x69778, x69777);
  nand n69780(x69780, x68680, x61234);
  nand n69781(x69781, x68745, x49689);
  nand n69782(x69782, x69781, x69780);
  nand n69783(x69783, x68671, x69776);
  nand n69784(x69784, x68670, x69779);
  nand n69785(x69785, x68671, x69782);
  nand n69786(x69786, x69785, x69784);
  nand n69787(x69787, x68636, x86548);
  nand n69788(x69788, x68639, x69786);
  nand n69789(x69789, x69788, x69787);
  nand n69790(x69790, x68680, x68147);
  nand n69791(x69791, x68745, x67154);
  nand n69792(x69792, x69791, x69790);
  nand n69793(x69793, x68680, x65679);
  nand n69794(x69794, x68745, x62436);
  nand n69795(x69795, x69794, x69793);
  nand n69796(x69796, x68745, x49693);
  nand n69797(x69797, x68671, x69792);
  nand n69798(x69798, x68670, x69795);
  nand n69799(x69799, x68671, x86549);
  nand n69800(x69800, x69799, x69798);
  nand n69801(x69801, x68636, x86550);
  nand n69802(x69802, x68639, x69800);
  nand n69803(x69803, x69802, x69801);
  nand n69804(x69804, x68680, x68151);
  nand n69805(x69805, x68745, x67158);
  nand n69806(x69806, x69805, x69804);
  nand n69807(x69807, x68680, x65682);
  nand n69808(x69808, x68745, x62443);
  nand n69809(x69809, x69808, x69807);
  nand n69810(x69810, x68745, x49697);
  nand n69811(x69811, x68671, x69806);
  nand n69812(x69812, x68670, x69809);
  nand n69813(x69813, x68671, x86551);
  nand n69814(x69814, x69813, x69812);
  nand n69815(x69815, x68636, x86552);
  nand n69816(x69816, x68639, x69814);
  nand n69817(x69817, x69816, x69815);
  nand n69818(x69818, x68680, x68155);
  nand n69819(x69819, x68745, x67162);
  nand n69820(x69820, x69819, x69818);
  nand n69821(x69821, x68680, x65685);
  nand n69822(x69822, x68745, x62450);
  nand n69823(x69823, x69822, x69821);
  nand n69824(x69824, x68745, x49701);
  nand n69825(x69825, x68671, x69820);
  nand n69826(x69826, x68670, x69823);
  nand n69827(x69827, x68671, x86553);
  nand n69828(x69828, x69827, x69826);
  nand n69829(x69829, x68636, x86554);
  nand n69830(x69830, x68639, x69828);
  nand n69831(x69831, x69830, x69829);
  nand n69832(x69832, x68680, x68159);
  nand n69833(x69833, x68745, x67166);
  nand n69834(x69834, x69833, x69832);
  nand n69835(x69835, x68680, x65688);
  nand n69836(x69836, x68745, x62457);
  nand n69837(x69837, x69836, x69835);
  nand n69838(x69838, x68745, x49705);
  nand n69839(x69839, x68671, x69834);
  nand n69840(x69840, x68670, x69837);
  nand n69841(x69841, x68671, x86555);
  nand n69842(x69842, x69841, x69840);
  nand n69843(x69843, x68636, x86556);
  nand n69844(x69844, x68639, x69842);
  nand n69845(x69845, x69844, x69843);
  nand n69846(x69846, x68680, x68163);
  nand n69847(x69847, x68745, x67170);
  nand n69848(x69848, x69847, x69846);
  nand n69849(x69849, x68680, x65691);
  nand n69850(x69850, x68745, x62464);
  nand n69851(x69851, x69850, x69849);
  nand n69852(x69852, x68745, x49709);
  nand n69853(x69853, x68671, x69848);
  nand n69854(x69854, x68670, x69851);
  nand n69855(x69855, x68671, x86557);
  nand n69856(x69856, x69855, x69854);
  nand n69857(x69857, x68636, x86558);
  nand n69858(x69858, x68639, x69856);
  nand n69859(x69859, x69858, x69857);
  nand n69860(x69860, x68680, x68167);
  nand n69861(x69861, x68745, x67174);
  nand n69862(x69862, x69861, x69860);
  nand n69863(x69863, x68680, x65694);
  nand n69864(x69864, x68745, x62471);
  nand n69865(x69865, x69864, x69863);
  nand n69866(x69866, x68745, x49713);
  nand n69867(x69867, x68671, x69862);
  nand n69868(x69868, x68670, x69865);
  nand n69869(x69869, x68671, x86559);
  nand n69870(x69870, x69869, x69868);
  nand n69871(x69871, x68636, x86560);
  nand n69872(x69872, x68639, x69870);
  nand n69873(x69873, x69872, x69871);
  nand n69874(x69874, x68680, x68171);
  nand n69875(x69875, x68745, x67178);
  nand n69876(x69876, x69875, x69874);
  nand n69877(x69877, x68680, x65697);
  nand n69878(x69878, x68745, x62478);
  nand n69879(x69879, x69878, x69877);
  nand n69880(x69880, x68745, x49717);
  nand n69881(x69881, x68671, x69876);
  nand n69882(x69882, x68670, x69879);
  nand n69883(x69883, x68671, x86561);
  nand n69884(x69884, x69883, x69882);
  nand n69885(x69885, x68636, x86562);
  nand n69886(x69886, x68639, x69884);
  nand n69887(x69887, x69886, x69885);
  nand n69888(x69888, x68680, x68175);
  nand n69889(x69889, x68745, x67182);
  nand n69890(x69890, x69889, x69888);
  nand n69891(x69891, x68680, x65700);
  nand n69892(x69892, x68745, x62485);
  nand n69893(x69893, x69892, x69891);
  nand n69894(x69894, x68745, x49721);
  nand n69895(x69895, x68671, x69890);
  nand n69896(x69896, x68670, x69893);
  nand n69897(x69897, x68671, x86563);
  nand n69898(x69898, x69897, x69896);
  nand n69899(x69899, x68636, x86564);
  nand n69900(x69900, x68639, x69898);
  nand n69901(x69901, x69900, x69899);
  nand n69902(x69902, x68680, x68179);
  nand n69903(x69903, x68745, x67186);
  nand n69904(x69904, x69903, x69902);
  nand n69905(x69905, x68680, x65703);
  nand n69906(x69906, x68745, x62492);
  nand n69907(x69907, x69906, x69905);
  nand n69908(x69908, x68745, x49725);
  nand n69909(x69909, x68671, x69904);
  nand n69910(x69910, x68670, x69907);
  nand n69911(x69911, x68671, x86565);
  nand n69912(x69912, x69911, x69910);
  nand n69913(x69913, x68636, x86566);
  nand n69914(x69914, x68639, x69912);
  nand n69915(x69915, x69914, x69913);
  nand n69916(x69916, x68680, x68183);
  nand n69917(x69917, x68745, x67190);
  nand n69918(x69918, x69917, x69916);
  nand n69919(x69919, x68680, x65706);
  nand n69920(x69920, x68745, x62499);
  nand n69921(x69921, x69920, x69919);
  nand n69922(x69922, x68745, x49729);
  nand n69923(x69923, x68671, x69918);
  nand n69924(x69924, x68670, x69921);
  nand n69925(x69925, x68671, x86567);
  nand n69926(x69926, x69925, x69924);
  nand n69927(x69927, x68636, x86568);
  nand n69928(x69928, x68639, x69926);
  nand n69929(x69929, x69928, x69927);
  nand n69930(x69930, x68680, x68187);
  nand n69931(x69931, x68745, x67194);
  nand n69932(x69932, x69931, x69930);
  nand n69933(x69933, x68680, x65709);
  nand n69934(x69934, x68745, x62506);
  nand n69935(x69935, x69934, x69933);
  nand n69936(x69936, x68745, x49733);
  nand n69937(x69937, x68671, x69932);
  nand n69938(x69938, x68670, x69935);
  nand n69939(x69939, x68671, x86569);
  nand n69940(x69940, x69939, x69938);
  nand n69941(x69941, x68636, x86570);
  nand n69942(x69942, x68639, x69940);
  nand n69943(x69943, x69942, x69941);
  nand n69944(x69944, x68680, x68191);
  nand n69945(x69945, x68745, x67198);
  nand n69946(x69946, x69945, x69944);
  nand n69947(x69947, x68680, x65712);
  nand n69948(x69948, x68745, x62513);
  nand n69949(x69949, x69948, x69947);
  nand n69950(x69950, x68745, x49737);
  nand n69951(x69951, x68671, x69946);
  nand n69952(x69952, x68670, x69949);
  nand n69953(x69953, x68671, x86571);
  nand n69954(x69954, x69953, x69952);
  nand n69955(x69955, x68636, x86572);
  nand n69956(x69956, x68639, x69954);
  nand n69957(x69957, x69956, x69955);
  nand n69958(x69958, x68680, x68195);
  nand n69959(x69959, x68745, x67202);
  nand n69960(x69960, x69959, x69958);
  nand n69961(x69961, x68680, x65715);
  nand n69962(x69962, x68745, x62520);
  nand n69963(x69963, x69962, x69961);
  nand n69964(x69964, x68745, x49741);
  nand n69965(x69965, x68671, x69960);
  nand n69966(x69966, x68670, x69963);
  nand n69967(x69967, x68671, x86573);
  nand n69968(x69968, x69967, x69966);
  nand n69969(x69969, x68636, x86574);
  nand n69970(x69970, x68639, x69968);
  nand n69971(x69971, x69970, x69969);
  nand n69972(x69972, x68680, x68199);
  nand n69973(x69973, x68745, x67206);
  nand n69974(x69974, x69973, x69972);
  nand n69975(x69975, x68680, x65718);
  nand n69976(x69976, x68745, x62527);
  nand n69977(x69977, x69976, x69975);
  nand n69978(x69978, x68745, x49745);
  nand n69979(x69979, x68671, x69974);
  nand n69980(x69980, x68670, x69977);
  nand n69981(x69981, x68671, x86575);
  nand n69982(x69982, x69981, x69980);
  nand n69983(x69983, x68636, x86576);
  nand n69984(x69984, x68639, x69982);
  nand n69985(x69985, x69984, x69983);
  nand n69986(x69986, x68680, x68203);
  nand n69987(x69987, x68745, x67210);
  nand n69988(x69988, x69987, x69986);
  nand n69989(x69989, x68680, x65721);
  nand n69990(x69990, x68745, x62534);
  nand n69991(x69991, x69990, x69989);
  nand n69992(x69992, x68745, x49749);
  nand n69993(x69993, x68671, x69988);
  nand n69994(x69994, x68670, x69991);
  nand n69995(x69995, x68671, x86577);
  nand n69996(x69996, x69995, x69994);
  nand n69997(x69997, x68636, x86578);
  nand n69998(x69998, x68639, x69996);
  nand n69999(x69999, x69998, x69997);
  nand n70000(x70000, x68680, x68207);
  nand n70001(x70001, x68745, x67214);
  nand n70002(x70002, x70001, x70000);
  nand n70003(x70003, x68680, x86347);
  nand n70004(x70004, x68745, x62541);
  nand n70005(x70005, x70004, x70003);
  nand n70006(x70006, x68745, x49753);
  nand n70007(x70007, x68671, x70002);
  nand n70008(x70008, x68670, x70005);
  nand n70009(x70009, x68671, x86579);
  nand n70010(x70010, x70009, x70008);
  nand n70011(x70011, x68636, x86580);
  nand n70012(x70012, x68639, x70010);
  nand n70013(x70013, x70012, x70011);
  nand n70014(x70014, x68680, x68211);
  nand n70015(x70015, x68745, x67218);
  nand n70016(x70016, x70015, x70014);
  nand n70017(x70017, x68680, x86348);
  nand n70018(x70018, x68745, x62548);
  nand n70019(x70019, x70018, x70017);
  nand n70020(x70020, x68745, x49757);
  nand n70021(x70021, x68671, x70016);
  nand n70022(x70022, x68670, x70019);
  nand n70023(x70023, x68671, x86581);
  nand n70024(x70024, x70023, x70022);
  nand n70025(x70025, x68636, x86582);
  nand n70026(x70026, x68639, x70024);
  nand n70027(x70027, x70026, x70025);
  nand n70028(x70028, x68680, x68215);
  nand n70029(x70029, x68745, x67222);
  nand n70030(x70030, x70029, x70028);
  nand n70031(x70031, x68680, x86349);
  nand n70032(x70032, x68745, x62555);
  nand n70033(x70033, x70032, x70031);
  nand n70034(x70034, x68745, x49761);
  nand n70035(x70035, x68671, x70030);
  nand n70036(x70036, x68670, x70033);
  nand n70037(x70037, x68671, x86583);
  nand n70038(x70038, x70037, x70036);
  nand n70039(x70039, x68636, x86584);
  nand n70040(x70040, x68639, x70038);
  nand n70041(x70041, x70040, x70039);
  nand n70042(x70042, x68680, x68219);
  nand n70043(x70043, x68745, x67226);
  nand n70044(x70044, x70043, x70042);
  nand n70045(x70045, x68680, x86350);
  nand n70046(x70046, x68745, x62562);
  nand n70047(x70047, x70046, x70045);
  nand n70048(x70048, x68745, x49765);
  nand n70049(x70049, x68671, x70044);
  nand n70050(x70050, x68670, x70047);
  nand n70051(x70051, x68671, x86585);
  nand n70052(x70052, x70051, x70050);
  nand n70053(x70053, x68636, x86586);
  nand n70054(x70054, x68639, x70052);
  nand n70055(x70055, x70054, x70053);
  nand n70056(x70056, x68680, x68223);
  nand n70057(x70057, x68745, x67230);
  nand n70058(x70058, x70057, x70056);
  nand n70059(x70059, x68680, x86351);
  nand n70060(x70060, x68745, x62569);
  nand n70061(x70061, x70060, x70059);
  nand n70062(x70062, x68745, x49769);
  nand n70063(x70063, x68671, x70058);
  nand n70064(x70064, x68670, x70061);
  nand n70065(x70065, x68671, x86587);
  nand n70066(x70066, x70065, x70064);
  nand n70067(x70067, x68636, x86588);
  nand n70068(x70068, x68639, x70066);
  nand n70069(x70069, x70068, x70067);
  nand n70070(x70070, x68680, x68227);
  nand n70071(x70071, x68745, x67234);
  nand n70072(x70072, x70071, x70070);
  nand n70073(x70073, x68680, x86352);
  nand n70074(x70074, x68745, x62576);
  nand n70075(x70075, x70074, x70073);
  nand n70076(x70076, x68745, x49773);
  nand n70077(x70077, x68671, x70072);
  nand n70078(x70078, x68670, x70075);
  nand n70079(x70079, x68671, x86589);
  nand n70080(x70080, x70079, x70078);
  nand n70081(x70081, x68636, x86590);
  nand n70082(x70082, x68639, x70080);
  nand n70083(x70083, x70082, x70081);
  nand n70084(x70084, x68680, x68231);
  nand n70085(x70085, x68745, x67238);
  nand n70086(x70086, x70085, x70084);
  nand n70087(x70087, x68680, x86353);
  nand n70088(x70088, x68745, x62583);
  nand n70089(x70089, x70088, x70087);
  nand n70090(x70090, x68745, x49777);
  nand n70091(x70091, x68671, x70086);
  nand n70092(x70092, x68670, x70089);
  nand n70093(x70093, x68671, x86591);
  nand n70094(x70094, x70093, x70092);
  nand n70095(x70095, x68636, x86592);
  nand n70096(x70096, x68639, x70094);
  nand n70097(x70097, x70096, x70095);
  nand n70098(x70098, x68680, x68235);
  nand n70099(x70099, x68745, x67242);
  nand n70100(x70100, x70099, x70098);
  nand n70101(x70101, x68680, x86354);
  nand n70102(x70102, x68745, x62590);
  nand n70103(x70103, x70102, x70101);
  nand n70104(x70104, x68745, x49781);
  nand n70105(x70105, x68671, x70100);
  nand n70106(x70106, x68670, x70103);
  nand n70107(x70107, x68671, x86593);
  nand n70108(x70108, x70107, x70106);
  nand n70109(x70109, x68636, x86594);
  nand n70110(x70110, x68639, x70108);
  nand n70111(x70111, x70110, x70109);
  nand n70112(x70112, x68680, x68239);
  nand n70113(x70113, x68745, x67246);
  nand n70114(x70114, x70113, x70112);
  nand n70115(x70115, x68680, x86355);
  nand n70116(x70116, x68745, x62597);
  nand n70117(x70117, x70116, x70115);
  nand n70118(x70118, x68745, x49785);
  nand n70119(x70119, x68671, x70114);
  nand n70120(x70120, x68670, x70117);
  nand n70121(x70121, x68671, x86595);
  nand n70122(x70122, x70121, x70120);
  nand n70123(x70123, x68636, x86596);
  nand n70124(x70124, x68639, x70122);
  nand n70125(x70125, x70124, x70123);
  nand n70126(x70126, x68680, x68243);
  nand n70127(x70127, x68745, x67250);
  nand n70128(x70128, x70127, x70126);
  nand n70129(x70129, x68680, x86356);
  nand n70130(x70130, x68745, x62604);
  nand n70131(x70131, x70130, x70129);
  nand n70132(x70132, x68745, x49789);
  nand n70133(x70133, x68671, x70128);
  nand n70134(x70134, x68670, x70131);
  nand n70135(x70135, x68671, x86597);
  nand n70136(x70136, x70135, x70134);
  nand n70137(x70137, x68636, x86598);
  nand n70138(x70138, x68639, x70136);
  nand n70139(x70139, x70138, x70137);
  nand n70140(x70140, x68680, x68247);
  nand n70141(x70141, x68745, x67254);
  nand n70142(x70142, x70141, x70140);
  nand n70143(x70143, x68680, x86357);
  nand n70144(x70144, x68745, x62611);
  nand n70145(x70145, x70144, x70143);
  nand n70146(x70146, x68745, x49793);
  nand n70147(x70147, x68671, x70142);
  nand n70148(x70148, x68670, x70145);
  nand n70149(x70149, x68671, x86599);
  nand n70150(x70150, x70149, x70148);
  nand n70151(x70151, x68636, x86600);
  nand n70152(x70152, x68639, x70150);
  nand n70153(x70153, x70152, x70151);
  nand n70154(x70154, x68680, x68251);
  nand n70155(x70155, x68745, x67258);
  nand n70156(x70156, x70155, x70154);
  nand n70157(x70157, x68680, x86358);
  nand n70158(x70158, x68745, x62618);
  nand n70159(x70159, x70158, x70157);
  nand n70160(x70160, x68745, x49797);
  nand n70161(x70161, x68671, x70156);
  nand n70162(x70162, x68670, x70159);
  nand n70163(x70163, x68671, x86601);
  nand n70164(x70164, x70163, x70162);
  nand n70165(x70165, x68636, x86602);
  nand n70166(x70166, x68639, x70164);
  nand n70167(x70167, x70166, x70165);
  nand n70168(x70168, x68680, x68255);
  nand n70169(x70169, x68745, x67262);
  nand n70170(x70170, x70169, x70168);
  nand n70171(x70171, x68680, x86359);
  nand n70172(x70172, x68745, x62625);
  nand n70173(x70173, x70172, x70171);
  nand n70174(x70174, x68745, x49801);
  nand n70175(x70175, x68671, x70170);
  nand n70176(x70176, x68670, x70173);
  nand n70177(x70177, x68671, x86603);
  nand n70178(x70178, x70177, x70176);
  nand n70179(x70179, x68636, x86604);
  nand n70180(x70180, x68639, x70178);
  nand n70181(x70181, x70180, x70179);
  nand n70182(x70182, x68680, x68259);
  nand n70183(x70183, x68745, x67266);
  nand n70184(x70184, x70183, x70182);
  nand n70185(x70185, x68680, x86360);
  nand n70186(x70186, x68745, x62632);
  nand n70187(x70187, x70186, x70185);
  nand n70188(x70188, x68745, x49805);
  nand n70189(x70189, x68671, x70184);
  nand n70190(x70190, x68670, x70187);
  nand n70191(x70191, x68671, x86605);
  nand n70192(x70192, x70191, x70190);
  nand n70193(x70193, x68636, x86606);
  nand n70194(x70194, x68639, x70192);
  nand n70195(x70195, x70194, x70193);
  nand n70196(x70196, x68680, x68263);
  nand n70197(x70197, x68745, x67270);
  nand n70198(x70198, x70197, x70196);
  nand n70199(x70199, x68680, x86361);
  nand n70200(x70200, x68745, x62639);
  nand n70201(x70201, x70200, x70199);
  nand n70202(x70202, x68745, x49809);
  nand n70203(x70203, x68671, x70198);
  nand n70204(x70204, x68670, x70201);
  nand n70205(x70205, x68671, x86607);
  nand n70206(x70206, x70205, x70204);
  nand n70207(x70207, x68636, x86608);
  nand n70208(x70208, x68639, x70206);
  nand n70209(x70209, x70208, x70207);
  nand n70210(x70210, x68680, x68267);
  nand n70211(x70211, x68745, x67274);
  nand n70212(x70212, x70211, x70210);
  nand n70213(x70213, x68680, x86362);
  nand n70214(x70214, x68745, x62646);
  nand n70215(x70215, x70214, x70213);
  nand n70216(x70216, x68745, x49813);
  nand n70217(x70217, x68671, x70212);
  nand n70218(x70218, x68670, x70215);
  nand n70219(x70219, x68671, x86609);
  nand n70220(x70220, x70219, x70218);
  nand n70221(x70221, x68636, x86610);
  nand n70222(x70222, x68639, x70220);
  nand n70223(x70223, x70222, x70221);
  nand n70224(x70224, x68680, x68271);
  nand n70225(x70225, x68745, x67278);
  nand n70226(x70226, x70225, x70224);
  nand n70227(x70227, x68680, x66346);
  nand n70228(x70228, x68745, x62653);
  nand n70229(x70229, x70228, x70227);
  nand n70230(x70230, x68680, x61363);
  nand n70231(x70231, x68745, x60656);
  nand n70232(x70232, x70231, x70230);
  nand n70233(x70233, x68671, x70226);
  nand n70234(x70234, x68670, x70229);
  nand n70235(x70235, x68671, x70232);
  nand n70236(x70236, x70235, x70234);
  nand n70237(x70237, x68636, x86611);
  nand n70238(x70238, x68639, x70236);
  nand n70239(x70239, x70238, x70237);
  nand n70240(x70240, x68680, x68275);
  nand n70241(x70241, x68745, x67282);
  nand n70242(x70242, x70241, x70240);
  nand n70243(x70243, x68680, x66349);
  nand n70244(x70244, x68745, x62660);
  nand n70245(x70245, x70244, x70243);
  nand n70246(x70246, x68745, x60660);
  nand n70247(x70247, x68671, x70242);
  nand n70248(x70248, x68670, x70245);
  nand n70249(x70249, x68671, x86612);
  nand n70250(x70250, x70249, x70248);
  nand n70251(x70251, x68636, x86613);
  nand n70252(x70252, x68639, x70250);
  nand n70253(x70253, x70252, x70251);
  nand n70254(x70254, x68680, x68279);
  nand n70255(x70255, x68745, x67286);
  nand n70256(x70256, x70255, x70254);
  nand n70257(x70257, x68680, x66352);
  nand n70258(x70258, x68745, x62667);
  nand n70259(x70259, x70258, x70257);
  nand n70260(x70260, x68745, x60664);
  nand n70261(x70261, x68671, x70256);
  nand n70262(x70262, x68670, x70259);
  nand n70263(x70263, x68671, x86614);
  nand n70264(x70264, x70263, x70262);
  nand n70265(x70265, x68636, x86615);
  nand n70266(x70266, x68639, x70264);
  nand n70267(x70267, x70266, x70265);
  nand n70268(x70268, x68680, x68283);
  nand n70269(x70269, x68745, x67290);
  nand n70270(x70270, x70269, x70268);
  nand n70271(x70271, x68680, x66355);
  nand n70272(x70272, x68745, x62674);
  nand n70273(x70273, x70272, x70271);
  nand n70274(x70274, x68745, x60668);
  nand n70275(x70275, x68671, x70270);
  nand n70276(x70276, x68670, x70273);
  nand n70277(x70277, x68671, x86616);
  nand n70278(x70278, x70277, x70276);
  nand n70279(x70279, x68636, x86617);
  nand n70280(x70280, x68639, x70278);
  nand n70281(x70281, x70280, x70279);
  nand n70282(x70282, x68680, x68287);
  nand n70283(x70283, x68745, x67294);
  nand n70284(x70284, x70283, x70282);
  nand n70285(x70285, x68680, x66358);
  nand n70286(x70286, x68745, x62681);
  nand n70287(x70287, x70286, x70285);
  nand n70288(x70288, x68745, x60672);
  nand n70289(x70289, x68671, x70284);
  nand n70290(x70290, x68670, x70287);
  nand n70291(x70291, x68671, x86618);
  nand n70292(x70292, x70291, x70290);
  nand n70293(x70293, x68636, x86619);
  nand n70294(x70294, x68639, x70292);
  nand n70295(x70295, x70294, x70293);
  nand n70296(x70296, x68680, x68291);
  nand n70297(x70297, x68745, x67298);
  nand n70298(x70298, x70297, x70296);
  nand n70299(x70299, x68680, x66361);
  nand n70300(x70300, x68745, x62688);
  nand n70301(x70301, x70300, x70299);
  nand n70302(x70302, x68745, x60676);
  nand n70303(x70303, x68671, x70298);
  nand n70304(x70304, x68670, x70301);
  nand n70305(x70305, x68671, x86620);
  nand n70306(x70306, x70305, x70304);
  nand n70307(x70307, x68636, x86621);
  nand n70308(x70308, x68639, x70306);
  nand n70309(x70309, x70308, x70307);
  nand n70310(x70310, x68680, x68295);
  nand n70311(x70311, x68745, x67302);
  nand n70312(x70312, x70311, x70310);
  nand n70313(x70313, x68680, x66364);
  nand n70314(x70314, x68745, x62695);
  nand n70315(x70315, x70314, x70313);
  nand n70316(x70316, x68745, x60680);
  nand n70317(x70317, x68671, x70312);
  nand n70318(x70318, x68670, x70315);
  nand n70319(x70319, x68671, x86622);
  nand n70320(x70320, x70319, x70318);
  nand n70321(x70321, x68636, x86623);
  nand n70322(x70322, x68639, x70320);
  nand n70323(x70323, x70322, x70321);
  nand n70324(x70324, x68680, x68299);
  nand n70325(x70325, x68745, x67306);
  nand n70326(x70326, x70325, x70324);
  nand n70327(x70327, x68680, x66367);
  nand n70328(x70328, x68745, x62702);
  nand n70329(x70329, x70328, x70327);
  nand n70330(x70330, x68745, x60684);
  nand n70331(x70331, x68671, x70326);
  nand n70332(x70332, x68670, x70329);
  nand n70333(x70333, x68671, x86624);
  nand n70334(x70334, x70333, x70332);
  nand n70335(x70335, x68636, x86625);
  nand n70336(x70336, x68639, x70334);
  nand n70337(x70337, x70336, x70335);
  nand n70338(x70338, x68680, x68303);
  nand n70339(x70339, x68745, x67310);
  nand n70340(x70340, x70339, x70338);
  nand n70341(x70341, x68680, x66370);
  nand n70342(x70342, x68745, x62709);
  nand n70343(x70343, x70342, x70341);
  nand n70344(x70344, x68745, x60688);
  nand n70345(x70345, x68671, x70340);
  nand n70346(x70346, x68670, x70343);
  nand n70347(x70347, x68671, x86626);
  nand n70348(x70348, x70347, x70346);
  nand n70349(x70349, x68636, x86627);
  nand n70350(x70350, x68639, x70348);
  nand n70351(x70351, x70350, x70349);
  nand n70352(x70352, x68680, x68307);
  nand n70353(x70353, x68745, x67314);
  nand n70354(x70354, x70353, x70352);
  nand n70355(x70355, x68680, x66373);
  nand n70356(x70356, x68745, x62716);
  nand n70357(x70357, x70356, x70355);
  nand n70358(x70358, x68745, x60692);
  nand n70359(x70359, x68671, x70354);
  nand n70360(x70360, x68670, x70357);
  nand n70361(x70361, x68671, x86628);
  nand n70362(x70362, x70361, x70360);
  nand n70363(x70363, x68636, x86629);
  nand n70364(x70364, x68639, x70362);
  nand n70365(x70365, x70364, x70363);
  nand n70366(x70366, x68680, x68311);
  nand n70367(x70367, x68745, x67318);
  nand n70368(x70368, x70367, x70366);
  nand n70369(x70369, x68680, x66376);
  nand n70370(x70370, x68745, x62723);
  nand n70371(x70371, x70370, x70369);
  nand n70372(x70372, x68745, x60696);
  nand n70373(x70373, x68671, x70368);
  nand n70374(x70374, x68670, x70371);
  nand n70375(x70375, x68671, x86630);
  nand n70376(x70376, x70375, x70374);
  nand n70377(x70377, x68636, x86631);
  nand n70378(x70378, x68639, x70376);
  nand n70379(x70379, x70378, x70377);
  nand n70380(x70380, x68680, x68315);
  nand n70381(x70381, x68745, x67322);
  nand n70382(x70382, x70381, x70380);
  nand n70383(x70383, x68680, x66379);
  nand n70384(x70384, x68745, x62730);
  nand n70385(x70385, x70384, x70383);
  nand n70386(x70386, x68745, x60700);
  nand n70387(x70387, x68671, x70382);
  nand n70388(x70388, x68670, x70385);
  nand n70389(x70389, x68671, x86632);
  nand n70390(x70390, x70389, x70388);
  nand n70391(x70391, x68636, x86633);
  nand n70392(x70392, x68639, x70390);
  nand n70393(x70393, x70392, x70391);
  nand n70394(x70394, x68680, x68319);
  nand n70395(x70395, x68745, x67326);
  nand n70396(x70396, x70395, x70394);
  nand n70397(x70397, x68680, x66382);
  nand n70398(x70398, x68745, x62737);
  nand n70399(x70399, x70398, x70397);
  nand n70400(x70400, x68745, x60704);
  nand n70401(x70401, x68671, x70396);
  nand n70402(x70402, x68670, x70399);
  nand n70403(x70403, x68671, x86634);
  nand n70404(x70404, x70403, x70402);
  nand n70405(x70405, x68636, x86635);
  nand n70406(x70406, x68639, x70404);
  nand n70407(x70407, x70406, x70405);
  nand n70408(x70408, x68680, x68323);
  nand n70409(x70409, x68745, x67330);
  nand n70410(x70410, x70409, x70408);
  nand n70411(x70411, x68680, x66385);
  nand n70412(x70412, x68745, x62744);
  nand n70413(x70413, x70412, x70411);
  nand n70414(x70414, x68745, x60708);
  nand n70415(x70415, x68671, x70410);
  nand n70416(x70416, x68670, x70413);
  nand n70417(x70417, x68671, x86636);
  nand n70418(x70418, x70417, x70416);
  nand n70419(x70419, x68636, x86637);
  nand n70420(x70420, x68639, x70418);
  nand n70421(x70421, x70420, x70419);
  nand n70422(x70422, x68680, x68327);
  nand n70423(x70423, x68745, x67334);
  nand n70424(x70424, x70423, x70422);
  nand n70425(x70425, x68680, x66388);
  nand n70426(x70426, x68745, x62751);
  nand n70427(x70427, x70426, x70425);
  nand n70428(x70428, x68745, x60712);
  nand n70429(x70429, x68671, x70424);
  nand n70430(x70430, x68670, x70427);
  nand n70431(x70431, x68671, x86638);
  nand n70432(x70432, x70431, x70430);
  nand n70433(x70433, x68636, x86639);
  nand n70434(x70434, x68639, x70432);
  nand n70435(x70435, x70434, x70433);
  nand n70436(x70436, x68680, x68331);
  nand n70437(x70437, x68745, x67338);
  nand n70438(x70438, x70437, x70436);
  nand n70439(x70439, x68680, x66391);
  nand n70440(x70440, x68745, x62758);
  nand n70441(x70441, x70440, x70439);
  nand n70442(x70442, x68745, x60716);
  nand n70443(x70443, x68671, x70438);
  nand n70444(x70444, x68670, x70441);
  nand n70445(x70445, x68671, x86640);
  nand n70446(x70446, x70445, x70444);
  nand n70447(x70447, x68636, x86641);
  nand n70448(x70448, x68639, x70446);
  nand n70449(x70449, x70448, x70447);
  nand n70450(x70450, x68680, x68335);
  nand n70451(x70451, x68745, x67342);
  nand n70452(x70452, x70451, x70450);
  nand n70453(x70453, x68680, x86380);
  nand n70454(x70454, x68745, x62765);
  nand n70455(x70455, x70454, x70453);
  nand n70456(x70456, x68745, x60720);
  nand n70457(x70457, x68671, x70452);
  nand n70458(x70458, x68670, x70455);
  nand n70459(x70459, x68671, x86642);
  nand n70460(x70460, x70459, x70458);
  nand n70461(x70461, x68636, x86643);
  nand n70462(x70462, x68639, x70460);
  nand n70463(x70463, x70462, x70461);
  nand n70464(x70464, x68680, x68339);
  nand n70465(x70465, x68745, x67346);
  nand n70466(x70466, x70465, x70464);
  nand n70467(x70467, x68680, x86381);
  nand n70468(x70468, x68745, x62772);
  nand n70469(x70469, x70468, x70467);
  nand n70470(x70470, x68745, x60724);
  nand n70471(x70471, x68671, x70466);
  nand n70472(x70472, x68670, x70469);
  nand n70473(x70473, x68671, x86644);
  nand n70474(x70474, x70473, x70472);
  nand n70475(x70475, x68636, x86645);
  nand n70476(x70476, x68639, x70474);
  nand n70477(x70477, x70476, x70475);
  nand n70478(x70478, x68680, x68343);
  nand n70479(x70479, x68745, x67350);
  nand n70480(x70480, x70479, x70478);
  nand n70481(x70481, x68680, x86382);
  nand n70482(x70482, x68745, x62779);
  nand n70483(x70483, x70482, x70481);
  nand n70484(x70484, x68745, x60728);
  nand n70485(x70485, x68671, x70480);
  nand n70486(x70486, x68670, x70483);
  nand n70487(x70487, x68671, x86646);
  nand n70488(x70488, x70487, x70486);
  nand n70489(x70489, x68636, x86647);
  nand n70490(x70490, x68639, x70488);
  nand n70491(x70491, x70490, x70489);
  nand n70492(x70492, x68680, x68347);
  nand n70493(x70493, x68745, x67354);
  nand n70494(x70494, x70493, x70492);
  nand n70495(x70495, x68680, x86383);
  nand n70496(x70496, x68745, x62786);
  nand n70497(x70497, x70496, x70495);
  nand n70498(x70498, x68745, x60732);
  nand n70499(x70499, x68671, x70494);
  nand n70500(x70500, x68670, x70497);
  nand n70501(x70501, x68671, x86648);
  nand n70502(x70502, x70501, x70500);
  nand n70503(x70503, x68636, x86649);
  nand n70504(x70504, x68639, x70502);
  nand n70505(x70505, x70504, x70503);
  nand n70506(x70506, x68680, x68351);
  nand n70507(x70507, x68745, x67358);
  nand n70508(x70508, x70507, x70506);
  nand n70509(x70509, x68680, x86384);
  nand n70510(x70510, x68745, x62793);
  nand n70511(x70511, x70510, x70509);
  nand n70512(x70512, x68745, x60736);
  nand n70513(x70513, x68671, x70508);
  nand n70514(x70514, x68670, x70511);
  nand n70515(x70515, x68671, x86650);
  nand n70516(x70516, x70515, x70514);
  nand n70517(x70517, x68636, x86651);
  nand n70518(x70518, x68639, x70516);
  nand n70519(x70519, x70518, x70517);
  nand n70520(x70520, x68680, x68355);
  nand n70521(x70521, x68745, x67362);
  nand n70522(x70522, x70521, x70520);
  nand n70523(x70523, x68680, x86385);
  nand n70524(x70524, x68745, x62800);
  nand n70525(x70525, x70524, x70523);
  nand n70526(x70526, x68745, x60740);
  nand n70527(x70527, x68671, x70522);
  nand n70528(x70528, x68670, x70525);
  nand n70529(x70529, x68671, x86652);
  nand n70530(x70530, x70529, x70528);
  nand n70531(x70531, x68636, x86653);
  nand n70532(x70532, x68639, x70530);
  nand n70533(x70533, x70532, x70531);
  nand n70534(x70534, x68680, x68359);
  nand n70535(x70535, x68745, x67366);
  nand n70536(x70536, x70535, x70534);
  nand n70537(x70537, x68680, x86386);
  nand n70538(x70538, x68745, x62807);
  nand n70539(x70539, x70538, x70537);
  nand n70540(x70540, x68745, x60744);
  nand n70541(x70541, x68671, x70536);
  nand n70542(x70542, x68670, x70539);
  nand n70543(x70543, x68671, x86654);
  nand n70544(x70544, x70543, x70542);
  nand n70545(x70545, x68636, x86655);
  nand n70546(x70546, x68639, x70544);
  nand n70547(x70547, x70546, x70545);
  nand n70548(x70548, x68680, x68363);
  nand n70549(x70549, x68745, x67370);
  nand n70550(x70550, x70549, x70548);
  nand n70551(x70551, x68680, x86387);
  nand n70552(x70552, x68745, x62814);
  nand n70553(x70553, x70552, x70551);
  nand n70554(x70554, x68745, x60748);
  nand n70555(x70555, x68671, x70550);
  nand n70556(x70556, x68670, x70553);
  nand n70557(x70557, x68671, x86656);
  nand n70558(x70558, x70557, x70556);
  nand n70559(x70559, x68636, x86657);
  nand n70560(x70560, x68639, x70558);
  nand n70561(x70561, x70560, x70559);
  nand n70562(x70562, x68680, x68367);
  nand n70563(x70563, x68745, x67374);
  nand n70564(x70564, x70563, x70562);
  nand n70565(x70565, x68680, x86388);
  nand n70566(x70566, x68745, x62821);
  nand n70567(x70567, x70566, x70565);
  nand n70568(x70568, x68745, x60752);
  nand n70569(x70569, x68671, x70564);
  nand n70570(x70570, x68670, x70567);
  nand n70571(x70571, x68671, x86658);
  nand n70572(x70572, x70571, x70570);
  nand n70573(x70573, x68636, x86659);
  nand n70574(x70574, x68639, x70572);
  nand n70575(x70575, x70574, x70573);
  nand n70576(x70576, x68680, x68371);
  nand n70577(x70577, x68745, x67378);
  nand n70578(x70578, x70577, x70576);
  nand n70579(x70579, x68680, x86389);
  nand n70580(x70580, x68745, x62828);
  nand n70581(x70581, x70580, x70579);
  nand n70582(x70582, x68745, x60756);
  nand n70583(x70583, x68671, x70578);
  nand n70584(x70584, x68670, x70581);
  nand n70585(x70585, x68671, x86660);
  nand n70586(x70586, x70585, x70584);
  nand n70587(x70587, x68636, x86661);
  nand n70588(x70588, x68639, x70586);
  nand n70589(x70589, x70588, x70587);
  nand n70590(x70590, x68680, x68375);
  nand n70591(x70591, x68745, x67382);
  nand n70592(x70592, x70591, x70590);
  nand n70593(x70593, x68680, x86390);
  nand n70594(x70594, x68745, x62835);
  nand n70595(x70595, x70594, x70593);
  nand n70596(x70596, x68745, x60760);
  nand n70597(x70597, x68671, x70592);
  nand n70598(x70598, x68670, x70595);
  nand n70599(x70599, x68671, x86662);
  nand n70600(x70600, x70599, x70598);
  nand n70601(x70601, x68636, x86663);
  nand n70602(x70602, x68639, x70600);
  nand n70603(x70603, x70602, x70601);
  nand n70604(x70604, x68680, x68379);
  nand n70605(x70605, x68745, x67386);
  nand n70606(x70606, x70605, x70604);
  nand n70607(x70607, x68680, x86391);
  nand n70608(x70608, x68745, x62842);
  nand n70609(x70609, x70608, x70607);
  nand n70610(x70610, x68745, x60764);
  nand n70611(x70611, x68671, x70606);
  nand n70612(x70612, x68670, x70609);
  nand n70613(x70613, x68671, x86664);
  nand n70614(x70614, x70613, x70612);
  nand n70615(x70615, x68636, x86665);
  nand n70616(x70616, x68639, x70614);
  nand n70617(x70617, x70616, x70615);
  nand n70618(x70618, x68680, x68383);
  nand n70619(x70619, x68745, x67390);
  nand n70620(x70620, x70619, x70618);
  nand n70621(x70621, x68680, x86392);
  nand n70622(x70622, x68745, x62849);
  nand n70623(x70623, x70622, x70621);
  nand n70624(x70624, x68745, x60768);
  nand n70625(x70625, x68671, x70620);
  nand n70626(x70626, x68670, x70623);
  nand n70627(x70627, x68671, x86666);
  nand n70628(x70628, x70627, x70626);
  nand n70629(x70629, x68636, x86667);
  nand n70630(x70630, x68639, x70628);
  nand n70631(x70631, x70630, x70629);
  nand n70632(x70632, x68680, x68387);
  nand n70633(x70633, x68745, x67394);
  nand n70634(x70634, x70633, x70632);
  nand n70635(x70635, x68680, x86393);
  nand n70636(x70636, x68745, x62856);
  nand n70637(x70637, x70636, x70635);
  nand n70638(x70638, x68745, x60772);
  nand n70639(x70639, x68671, x70634);
  nand n70640(x70640, x68670, x70637);
  nand n70641(x70641, x68671, x86668);
  nand n70642(x70642, x70641, x70640);
  nand n70643(x70643, x68636, x86669);
  nand n70644(x70644, x68639, x70642);
  nand n70645(x70645, x70644, x70643);
  nand n70646(x70646, x68680, x68391);
  nand n70647(x70647, x68745, x67398);
  nand n70648(x70648, x70647, x70646);
  nand n70649(x70649, x68680, x86394);
  nand n70650(x70650, x68745, x62863);
  nand n70651(x70651, x70650, x70649);
  nand n70652(x70652, x68745, x60776);
  nand n70653(x70653, x68671, x70648);
  nand n70654(x70654, x68670, x70651);
  nand n70655(x70655, x68671, x86670);
  nand n70656(x70656, x70655, x70654);
  nand n70657(x70657, x68636, x86671);
  nand n70658(x70658, x68639, x70656);
  nand n70659(x70659, x70658, x70657);
  nand n70660(x70660, x68680, x68395);
  nand n70661(x70661, x68745, x67402);
  nand n70662(x70662, x70661, x70660);
  nand n70663(x70663, x68680, x86395);
  nand n70664(x70664, x68745, x62870);
  nand n70665(x70665, x70664, x70663);
  nand n70666(x70666, x68745, x60780);
  nand n70667(x70667, x68671, x70662);
  nand n70668(x70668, x68670, x70665);
  nand n70669(x70669, x68671, x86672);
  nand n70670(x70670, x70669, x70668);
  nand n70671(x70671, x68636, x86673);
  nand n70672(x70672, x68639, x70670);
  nand n70673(x70673, x70672, x70671);
  nand n70674(x70674, x68680, x68426);
  nand n70675(x70675, x68745, x67433);
  nand n70676(x70676, x70675, x70674);
  nand n70677(x70677, x68680, x66441);
  nand n70678(x70678, x68745, x62901);
  nand n70679(x70679, x70678, x70677);
  nand n70680(x70680, x68680, x61395);
  nand n70681(x70681, x68745, x60812);
  nand n70682(x70682, x70681, x70680);
  nand n70683(x70683, x68671, x70676);
  nand n70684(x70684, x68670, x70679);
  nand n70685(x70685, x68671, x70682);
  nand n70686(x70686, x70685, x70684);
  nand n70687(x70687, x68636, x86674);
  nand n70688(x70688, x68639, x70686);
  nand n70689(x70689, x70688, x70687);
  nand n70690(x70690, x68680, x68430);
  nand n70691(x70691, x68745, x67437);
  nand n70692(x70692, x70691, x70690);
  nand n70693(x70693, x68680, x66445);
  nand n70694(x70694, x68745, x62905);
  nand n70695(x70695, x70694, x70693);
  nand n70696(x70696, x68680, x61399);
  nand n70697(x70697, x68745, x60816);
  nand n70698(x70698, x70697, x70696);
  nand n70699(x70699, x68671, x70692);
  nand n70700(x70700, x68670, x70695);
  nand n70701(x70701, x68671, x70698);
  nand n70702(x70702, x70701, x70700);
  nand n70703(x70703, x68636, x86675);
  nand n70704(x70704, x68639, x70702);
  nand n70705(x70705, x70704, x70703);
  nand n70706(x70706, x68680, x68434);
  nand n70707(x70707, x68745, x67441);
  nand n70708(x70708, x70707, x70706);
  nand n70709(x70709, x68680, x66449);
  nand n70710(x70710, x68745, x62909);
  nand n70711(x70711, x70710, x70709);
  nand n70712(x70712, x68680, x61403);
  nand n70713(x70713, x68745, x60820);
  nand n70714(x70714, x70713, x70712);
  nand n70715(x70715, x68671, x70708);
  nand n70716(x70716, x68670, x70711);
  nand n70717(x70717, x68671, x70714);
  nand n70718(x70718, x70717, x70716);
  nand n70719(x70719, x68636, x86676);
  nand n70720(x70720, x68639, x70718);
  nand n70721(x70721, x70720, x70719);
  nand n70722(x70722, x68680, x68402);
  nand n70723(x70723, x68745, x67409);
  nand n70724(x70724, x70723, x70722);
  nand n70725(x70725, x68680, x66417);
  nand n70726(x70726, x68745, x62877);
  nand n70727(x70727, x70726, x70725);
  nand n70728(x70728, x68680, x61371);
  nand n70729(x70729, x68745, x60788);
  nand n70730(x70730, x70729, x70728);
  nand n70731(x70731, x68671, x70724);
  nand n70732(x70732, x68670, x70727);
  nand n70733(x70733, x68671, x70730);
  nand n70734(x70734, x70733, x70732);
  nand n70735(x70735, x68636, x86677);
  nand n70736(x70736, x68639, x70734);
  nand n70737(x70737, x70736, x70735);
  nand n70738(x70738, x68680, x68406);
  nand n70739(x70739, x68745, x67413);
  nand n70740(x70740, x70739, x70738);
  nand n70741(x70741, x68680, x66421);
  nand n70742(x70742, x68745, x62881);
  nand n70743(x70743, x70742, x70741);
  nand n70744(x70744, x68680, x61375);
  nand n70745(x70745, x68745, x60792);
  nand n70746(x70746, x70745, x70744);
  nand n70747(x70747, x68671, x70740);
  nand n70748(x70748, x68670, x70743);
  nand n70749(x70749, x68671, x70746);
  nand n70750(x70750, x70749, x70748);
  nand n70751(x70751, x68636, x86678);
  nand n70752(x70752, x68639, x70750);
  nand n70753(x70753, x70752, x70751);
  nand n70754(x70754, x68680, x68410);
  nand n70755(x70755, x68745, x67417);
  nand n70756(x70756, x70755, x70754);
  nand n70757(x70757, x68680, x66425);
  nand n70758(x70758, x68745, x62885);
  nand n70759(x70759, x70758, x70757);
  nand n70760(x70760, x68680, x61379);
  nand n70761(x70761, x68745, x60796);
  nand n70762(x70762, x70761, x70760);
  nand n70763(x70763, x68671, x70756);
  nand n70764(x70764, x68670, x70759);
  nand n70765(x70765, x68671, x70762);
  nand n70766(x70766, x70765, x70764);
  nand n70767(x70767, x68636, x86679);
  nand n70768(x70768, x68639, x70766);
  nand n70769(x70769, x70768, x70767);
  nand n70770(x70770, x68680, x68414);
  nand n70771(x70771, x68745, x67421);
  nand n70772(x70772, x70771, x70770);
  nand n70773(x70773, x68680, x66429);
  nand n70774(x70774, x68745, x62889);
  nand n70775(x70775, x70774, x70773);
  nand n70776(x70776, x68680, x61383);
  nand n70777(x70777, x68745, x60800);
  nand n70778(x70778, x70777, x70776);
  nand n70779(x70779, x68671, x70772);
  nand n70780(x70780, x68670, x70775);
  nand n70781(x70781, x68671, x70778);
  nand n70782(x70782, x70781, x70780);
  nand n70783(x70783, x68636, x86680);
  nand n70784(x70784, x68639, x70782);
  nand n70785(x70785, x70784, x70783);
  nand n70786(x70786, x68680, x68418);
  nand n70787(x70787, x68745, x67425);
  nand n70788(x70788, x70787, x70786);
  nand n70789(x70789, x68680, x66433);
  nand n70790(x70790, x68745, x62893);
  nand n70791(x70791, x70790, x70789);
  nand n70792(x70792, x68680, x61387);
  nand n70793(x70793, x68745, x60804);
  nand n70794(x70794, x70793, x70792);
  nand n70795(x70795, x68671, x70788);
  nand n70796(x70796, x68670, x70791);
  nand n70797(x70797, x68671, x70794);
  nand n70798(x70798, x70797, x70796);
  nand n70799(x70799, x68636, x86681);
  nand n70800(x70800, x68639, x70798);
  nand n70801(x70801, x70800, x70799);
  nand n70802(x70802, x68680, x68422);
  nand n70803(x70803, x68745, x67429);
  nand n70804(x70804, x70803, x70802);
  nand n70805(x70805, x68680, x66437);
  nand n70806(x70806, x68745, x62897);
  nand n70807(x70807, x70806, x70805);
  nand n70808(x70808, x68680, x61391);
  nand n70809(x70809, x68745, x60808);
  nand n70810(x70810, x70809, x70808);
  nand n70811(x70811, x68671, x70804);
  nand n70812(x70812, x68670, x70807);
  nand n70813(x70813, x68671, x70810);
  nand n70814(x70814, x70813, x70812);
  nand n70815(x70815, x68636, x86682);
  nand n70816(x70816, x68639, x70814);
  nand n70817(x70817, x70816, x70815);
  nand n70818(x70818, x68701, x67887);
  nand n70819(x70819, x68810, x66894);
  nand n70820(x70820, x70819, x70818);
  nand n70821(x70821, x68701, x64274);
  nand n70822(x70822, x68810, x61981);
  nand n70823(x70823, x70822, x70821);
  nand n70824(x70824, x68701, x60976);
  nand n70825(x70825, x68810, x27755);
  nand n70826(x70826, x70825, x70824);
  nand n70827(x70827, x68692, x70820);
  nand n70828(x70828, x68691, x70823);
  nand n70829(x70829, x68692, x70826);
  nand n70830(x70830, x70829, x70828);
  nand n70831(x70831, x68651, x86683);
  nand n70832(x70832, x68654, x70830);
  nand n70833(x70833, x70832, x70831);
  nand n70834(x70834, x68701, x68015);
  nand n70835(x70835, x68810, x67022);
  nand n70836(x70836, x70835, x70834);
  nand n70837(x70837, x68701, x65006);
  nand n70838(x70838, x68810, x62205);
  nand n70839(x70839, x70838, x70837);
  nand n70840(x70840, x68701, x61105);
  nand n70841(x70841, x68810, x38722);
  nand n70842(x70842, x70841, x70840);
  nand n70843(x70843, x68692, x70836);
  nand n70844(x70844, x68691, x70839);
  nand n70845(x70845, x68692, x70842);
  nand n70846(x70846, x70845, x70844);
  nand n70847(x70847, x68651, x86684);
  nand n70848(x70848, x68654, x70846);
  nand n70849(x70849, x70848, x70847);
  nand n70850(x70850, x68701, x68143);
  nand n70851(x70851, x68810, x67150);
  nand n70852(x70852, x70851, x70850);
  nand n70853(x70853, x68701, x65676);
  nand n70854(x70854, x68810, x62429);
  nand n70855(x70855, x70854, x70853);
  nand n70856(x70856, x68701, x61234);
  nand n70857(x70857, x68810, x49689);
  nand n70858(x70858, x70857, x70856);
  nand n70859(x70859, x68692, x70852);
  nand n70860(x70860, x68691, x70855);
  nand n70861(x70861, x68692, x70858);
  nand n70862(x70862, x70861, x70860);
  nand n70863(x70863, x68651, x86685);
  nand n70864(x70864, x68654, x70862);
  nand n70865(x70865, x70864, x70863);
  nand n70866(x70866, x68701, x68271);
  nand n70867(x70867, x68810, x67278);
  nand n70868(x70868, x70867, x70866);
  nand n70869(x70869, x68701, x66346);
  nand n70870(x70870, x68810, x62653);
  nand n70871(x70871, x70870, x70869);
  nand n70872(x70872, x68701, x61363);
  nand n70873(x70873, x68810, x60656);
  nand n70874(x70874, x70873, x70872);
  nand n70875(x70875, x68692, x70868);
  nand n70876(x70876, x68691, x70871);
  nand n70877(x70877, x68692, x70874);
  nand n70878(x70878, x70877, x70876);
  nand n70879(x70879, x68651, x86686);
  nand n70880(x70880, x68654, x70878);
  nand n70881(x70881, x70880, x70879);
  nand n70882(x70882, x68701, x68426);
  nand n70883(x70883, x68810, x67433);
  nand n70884(x70884, x70883, x70882);
  nand n70885(x70885, x68701, x66441);
  nand n70886(x70886, x68810, x62901);
  nand n70887(x70887, x70886, x70885);
  nand n70888(x70888, x68701, x61395);
  nand n70889(x70889, x68810, x60812);
  nand n70890(x70890, x70889, x70888);
  nand n70891(x70891, x68692, x70884);
  nand n70892(x70892, x68691, x70887);
  nand n70893(x70893, x68692, x70890);
  nand n70894(x70894, x70893, x70892);
  nand n70895(x70895, x68651, x86687);
  nand n70896(x70896, x68654, x70894);
  nand n70897(x70897, x70896, x70895);
  nand n70898(x70898, x68701, x68430);
  nand n70899(x70899, x68810, x67437);
  nand n70900(x70900, x70899, x70898);
  nand n70901(x70901, x68701, x66445);
  nand n70902(x70902, x68810, x62905);
  nand n70903(x70903, x70902, x70901);
  nand n70904(x70904, x68701, x61399);
  nand n70905(x70905, x68810, x60816);
  nand n70906(x70906, x70905, x70904);
  nand n70907(x70907, x68692, x70900);
  nand n70908(x70908, x68691, x70903);
  nand n70909(x70909, x68692, x70906);
  nand n70910(x70910, x70909, x70908);
  nand n70911(x70911, x68651, x86688);
  nand n70912(x70912, x68654, x70910);
  nand n70913(x70913, x70912, x70911);
  nand n70914(x70914, x68701, x68434);
  nand n70915(x70915, x68810, x67441);
  nand n70916(x70916, x70915, x70914);
  nand n70917(x70917, x68701, x66449);
  nand n70918(x70918, x68810, x62909);
  nand n70919(x70919, x70918, x70917);
  nand n70920(x70920, x68701, x61403);
  nand n70921(x70921, x68810, x60820);
  nand n70922(x70922, x70921, x70920);
  nand n70923(x70923, x68692, x70916);
  nand n70924(x70924, x68691, x70919);
  nand n70925(x70925, x68692, x70922);
  nand n70926(x70926, x70925, x70924);
  nand n70927(x70927, x68651, x86689);
  nand n70928(x70928, x68654, x70926);
  nand n70929(x70929, x70928, x70927);
  nand n70930(x70930, x68701, x68402);
  nand n70931(x70931, x68810, x67409);
  nand n70932(x70932, x70931, x70930);
  nand n70933(x70933, x68701, x66417);
  nand n70934(x70934, x68810, x62877);
  nand n70935(x70935, x70934, x70933);
  nand n70936(x70936, x68701, x61371);
  nand n70937(x70937, x68810, x60788);
  nand n70938(x70938, x70937, x70936);
  nand n70939(x70939, x68692, x70932);
  nand n70940(x70940, x68691, x70935);
  nand n70941(x70941, x68692, x70938);
  nand n70942(x70942, x70941, x70940);
  nand n70943(x70943, x68651, x86690);
  nand n70944(x70944, x68654, x70942);
  nand n70945(x70945, x70944, x70943);
  nand n70946(x70946, x68701, x68406);
  nand n70947(x70947, x68810, x67413);
  nand n70948(x70948, x70947, x70946);
  nand n70949(x70949, x68701, x66421);
  nand n70950(x70950, x68810, x62881);
  nand n70951(x70951, x70950, x70949);
  nand n70952(x70952, x68701, x61375);
  nand n70953(x70953, x68810, x60792);
  nand n70954(x70954, x70953, x70952);
  nand n70955(x70955, x68692, x70948);
  nand n70956(x70956, x68691, x70951);
  nand n70957(x70957, x68692, x70954);
  nand n70958(x70958, x70957, x70956);
  nand n70959(x70959, x68651, x86691);
  nand n70960(x70960, x68654, x70958);
  nand n70961(x70961, x70960, x70959);
  nand n70962(x70962, x68701, x68410);
  nand n70963(x70963, x68810, x67417);
  nand n70964(x70964, x70963, x70962);
  nand n70965(x70965, x68701, x66425);
  nand n70966(x70966, x68810, x62885);
  nand n70967(x70967, x70966, x70965);
  nand n70968(x70968, x68701, x61379);
  nand n70969(x70969, x68810, x60796);
  nand n70970(x70970, x70969, x70968);
  nand n70971(x70971, x68692, x70964);
  nand n70972(x70972, x68691, x70967);
  nand n70973(x70973, x68692, x70970);
  nand n70974(x70974, x70973, x70972);
  nand n70975(x70975, x68651, x86692);
  nand n70976(x70976, x68654, x70974);
  nand n70977(x70977, x70976, x70975);
  nand n70978(x70978, x68701, x68414);
  nand n70979(x70979, x68810, x67421);
  nand n70980(x70980, x70979, x70978);
  nand n70981(x70981, x68701, x66429);
  nand n70982(x70982, x68810, x62889);
  nand n70983(x70983, x70982, x70981);
  nand n70984(x70984, x68701, x61383);
  nand n70985(x70985, x68810, x60800);
  nand n70986(x70986, x70985, x70984);
  nand n70987(x70987, x68692, x70980);
  nand n70988(x70988, x68691, x70983);
  nand n70989(x70989, x68692, x70986);
  nand n70990(x70990, x70989, x70988);
  nand n70991(x70991, x68651, x86693);
  nand n70992(x70992, x68654, x70990);
  nand n70993(x70993, x70992, x70991);
  nand n70994(x70994, x68701, x68418);
  nand n70995(x70995, x68810, x67425);
  nand n70996(x70996, x70995, x70994);
  nand n70997(x70997, x68701, x66433);
  nand n70998(x70998, x68810, x62893);
  nand n70999(x70999, x70998, x70997);
  nand n71000(x71000, x68701, x61387);
  nand n71001(x71001, x68810, x60804);
  nand n71002(x71002, x71001, x71000);
  nand n71003(x71003, x68692, x70996);
  nand n71004(x71004, x68691, x70999);
  nand n71005(x71005, x68692, x71002);
  nand n71006(x71006, x71005, x71004);
  nand n71007(x71007, x68651, x86694);
  nand n71008(x71008, x68654, x71006);
  nand n71009(x71009, x71008, x71007);
  nand n71010(x71010, x68701, x68422);
  nand n71011(x71011, x68810, x67429);
  nand n71012(x71012, x71011, x71010);
  nand n71013(x71013, x68701, x66437);
  nand n71014(x71014, x68810, x62897);
  nand n71015(x71015, x71014, x71013);
  nand n71016(x71016, x68701, x61391);
  nand n71017(x71017, x68810, x60808);
  nand n71018(x71018, x71017, x71016);
  nand n71019(x71019, x68692, x71012);
  nand n71020(x71020, x68691, x71015);
  nand n71021(x71021, x68692, x71018);
  nand n71022(x71022, x71021, x71020);
  nand n71023(x71023, x68651, x86695);
  nand n71024(x71024, x68654, x71022);
  nand n71025(x71025, x71024, x71023);
  nand n71026(x71026, x70737, x14990);
  nand n71029(x71029, x71028, x71027);
  nand n71030(x71030, x71029, x71026);
  nand n71031(x71031, x70753, x15011);
  nand n71034(x71034, x71033, x71032);
  nand n71035(x71035, x71034, x71031);
  nand n71036(x71036, x70769, x15032);
  nand n71039(x71039, x71038, x71037);
  nand n71040(x71040, x71039, x71036);
  nand n71041(x71041, x70785, x15053);
  nand n71044(x71044, x71043, x71042);
  nand n71045(x71045, x71044, x71041);
  nand n71046(x71046, x70801, x15074);
  nand n71049(x71049, x71048, x71047);
  nand n71050(x71050, x71049, x71046);
  nand n71051(x71051, x70817, x15095);
  nand n71054(x71054, x71053, x71052);
  nand n71055(x71055, x71054, x71051);
  nand n71056(x71056, x71050, x71055);
  nand n71058(x71058, x71040, x71045);
  nand n71060(x71060, x71030, x71035);
  nand n71062(x71062, x71059, x71057);
  nand n71064(x71064, x71063, x71061);
  nand n71066(x71066, x68644, x71065);
  nand n71068(x71068, x71067, x68760);
  nand n71070(x71070, x71067, x68776);
  nand n71072(x71072, x71067, x68792);
  nand n71074(x71074, x71067, x68808);
  nand n71076(x71076, x70945, x2137);
  nand n71079(x71079, x71078, x71077);
  nand n71080(x71080, x71079, x71076);
  nand n71081(x71081, x70961, x2158);
  nand n71084(x71084, x71083, x71082);
  nand n71085(x71085, x71084, x71081);
  nand n71086(x71086, x70977, x2179);
  nand n71089(x71089, x71088, x71087);
  nand n71090(x71090, x71089, x71086);
  nand n71091(x71091, x70993, x2200);
  nand n71094(x71094, x71093, x71092);
  nand n71095(x71095, x71094, x71091);
  nand n71096(x71096, x71009, x2221);
  nand n71099(x71099, x71098, x71097);
  nand n71100(x71100, x71099, x71096);
  nand n71101(x71101, x71025, x2242);
  nand n71104(x71104, x71103, x71102);
  nand n71105(x71105, x71104, x71101);
  nand n71106(x71106, x71100, x71105);
  nand n71108(x71108, x71090, x71095);
  nand n71110(x71110, x71080, x71085);
  nand n71112(x71112, x71109, x71107);
  nand n71114(x71114, x71113, x71111);
  nand n71116(x71116, x68659, x71115);
  nand n71118(x71118, x71117, x68825);
  nand n71120(x71120, x71117, x68841);
  nand n71122(x71122, x71117, x68857);
  nand n71124(x71124, x71117, x68873);
  nand n71128(x71128, x71127, x71126);
  nand n71129(x71129, x1895, x1898);
  nand n71130(x71130, x1900, x14745);
  nand n71131(x71131, x14750, x14753);
  nand n71134(x71134, x71133, x71132);
  nand n71137(x71137, x71136, x71135);
  nand n71140(x71140, x71139, x71138);
  nand n71141(x71141, x678, x1);
  nand n71142(x71142, x15228, x71141);
  nand n71143(x71143, x0, x83429);
  nand n71144(x71144, x1, x86696);
  nand n71145(x71145, x71140, x71147);
  nand n71146(x71146, x71145, x71144);
  nand n71148(x71148, x0, x83435);
  nand n71149(x71149, x1, x86697);
  nand n71150(x71150, x71140, x71152);
  nand n71151(x71151, x71150, x71149);
  nand n71153(x71153, x0, x83441);
  nand n71154(x71154, x1, x86698);
  nand n71155(x71155, x71140, x71157);
  nand n71156(x71156, x71155, x71154);
  nand n71158(x71158, x0, x83447);
  nand n71159(x71159, x1, x86699);
  nand n71160(x71160, x71140, x71162);
  nand n71161(x71161, x71160, x71159);
  nand n71163(x71163, x0, x83452);
  nand n71164(x71164, x1, x86700);
  nand n71165(x71165, x71140, x71167);
  nand n71166(x71166, x71165, x71164);
  nand n71168(x71168, x0, x83456);
  nand n71169(x71169, x1, x86701);
  nand n71170(x71170, x71140, x71172);
  nand n71171(x71171, x71170, x71169);
  nand n71173(x71173, x0, x83459);
  nand n71174(x71174, x1, x86702);
  nand n71175(x71175, x71140, x71177);
  nand n71176(x71176, x71175, x71174);
  nand n71178(x71178, x0, x83464);
  nand n71179(x71179, x1, x86703);
  nand n71180(x71180, x71140, x71182);
  nand n71181(x71181, x71180, x71179);
  nand n71183(x71183, x71140, x71185);
  nand n71184(x71184, x71183, x71179);
  nand n71186(x71186, x71140, x71188);
  nand n71187(x71187, x71186, x71179);
  nand n71189(x71189, x71140, x71191);
  nand n71190(x71190, x71189, x71179);
  nand n71192(x71192, x71140, x71194);
  nand n71193(x71193, x71192, x71179);
  nand n71195(x71195, x71140, x71197);
  nand n71196(x71196, x71195, x71179);
  nand n71198(x71198, x0, x83468);
  nand n71199(x71199, x1, x86704);
  nand n71200(x71200, x71140, x71202);
  nand n71201(x71201, x71200, x71199);
  nand n71203(x71203, x71140, x71205);
  nand n71204(x71204, x71203, x71199);
  nand n71206(x71206, x0, x83471);
  nand n71207(x71207, x1, x86705);
  nand n71208(x71208, x71140, x71210);
  nand n71209(x71209, x71208, x71207);
  nand n71211(x71211, x0, x83475);
  nand n71212(x71212, x1, x86706);
  nand n71213(x71213, x71140, x71215);
  nand n71214(x71214, x71213, x71212);
  nand n71216(x71216, x0, x83479);
  nand n71217(x71217, x1, x86707);
  nand n71218(x71218, x71140, x71220);
  nand n71219(x71219, x71218, x71217);
  nand n71221(x71221, x0, x83482);
  nand n71222(x71222, x1, x86708);
  nand n71223(x71223, x71140, x71225);
  nand n71224(x71224, x71223, x71222);
  nand n71226(x71226, x0, x83487);
  nand n71227(x71227, x1, x86709);
  nand n71228(x71228, x71140, x71230);
  nand n71229(x71229, x71228, x71227);
  nand n71231(x71231, x0, x83489);
  nand n71232(x71232, x1, x86710);
  nand n71233(x71233, x71140, x71235);
  nand n71234(x71234, x71233, x71232);
  nand n71236(x71236, x0, x83492);
  nand n71237(x71237, x1, x86711);
  nand n71238(x71238, x71140, x71240);
  nand n71239(x71239, x71238, x71237);
  nand n71241(x71241, x0, x83495);
  nand n71242(x71242, x1, x86712);
  nand n71243(x71243, x71140, x71245);
  nand n71244(x71244, x71243, x71242);
  nand n71246(x71246, x0, x83497);
  nand n71247(x71247, x1, x86713);
  nand n71248(x71248, x71140, x71250);
  nand n71249(x71249, x71248, x71247);
  nand n71251(x71251, x0, x83499);
  nand n71252(x71252, x1, x86714);
  nand n71253(x71253, x71140, x71255);
  nand n71254(x71254, x71253, x71252);
  nand n71256(x71256, x0, x83501);
  nand n71257(x71257, x1, x86715);
  nand n71258(x71258, x71140, x71260);
  nand n71259(x71259, x71258, x71257);
  nand n71261(x71261, x0, x83503);
  nand n71262(x71262, x1, x86716);
  nand n71263(x71263, x71140, x71265);
  nand n71264(x71264, x71263, x71262);
  nand n71266(x71266, x0, x83506);
  nand n71267(x71267, x1, x86717);
  nand n71268(x71268, x71140, x71270);
  nand n71269(x71269, x71268, x71267);
  nand n71271(x71271, x0, x83512);
  nand n71272(x71272, x1, x86718);
  nand n71273(x71273, x71140, x71275);
  nand n71274(x71274, x71273, x71272);
  nand n71276(x71276, x71140, x71277);
  nand n71278(x71278, x71140, x71279);
  nand n71280(x71280, x0, x83515);
  nand n71281(x71281, x1, x86721);
  nand n71282(x71282, x71140, x71284);
  nand n71283(x71283, x71282, x71281);
  nand n71285(x71285, x15228, x602);
  nand n71286(x71286, x1, x86722);
  nand n71287(x71287, x71140, x71289);
  nand n71288(x71288, x71287, x71286);
  nand n71290(x71290, x15228, x603);
  nand n71291(x71291, x1, x86723);
  nand n71292(x71292, x71140, x71294);
  nand n71293(x71293, x71292, x71291);
  nand n71295(x71295, x15228, x604);
  nand n71296(x71296, x1, x86724);
  nand n71297(x71297, x71140, x71299);
  nand n71298(x71298, x71297, x71296);
  nand n71300(x71300, x15228, x605);
  nand n71301(x71301, x1, x86725);
  nand n71302(x71302, x71140, x71304);
  nand n71303(x71303, x71302, x71301);
  nand n71305(x71305, x15228, x606);
  nand n71306(x71306, x1, x86726);
  nand n71307(x71307, x71140, x71309);
  nand n71308(x71308, x71307, x71306);
  nand n71310(x71310, x15228, x607);
  nand n71311(x71311, x1, x86727);
  nand n71312(x71312, x71140, x71314);
  nand n71313(x71313, x71312, x71311);
  nand n71315(x71315, x15228, x608);
  nand n71316(x71316, x1, x86728);
  nand n71317(x71317, x71140, x71319);
  nand n71318(x71318, x71317, x71316);
  nand n71320(x71320, x15228, x609);
  nand n71321(x71321, x1, x86729);
  nand n71322(x71322, x71140, x71324);
  nand n71323(x71323, x71322, x71321);
  nand n71325(x71325, x15228, x610);
  nand n71326(x71326, x1, x86730);
  nand n71327(x71327, x71140, x71329);
  nand n71328(x71328, x71327, x71326);
  nand n71330(x71330, x15228, x611);
  nand n71331(x71331, x1, x86731);
  nand n71332(x71332, x71140, x71334);
  nand n71333(x71333, x71332, x71331);
  nand n71335(x71335, x15228, x612);
  nand n71336(x71336, x1, x86732);
  nand n71337(x71337, x71140, x71339);
  nand n71338(x71338, x71337, x71336);
  nand n71340(x71340, x15228, x613);
  nand n71341(x71341, x1, x86733);
  nand n71342(x71342, x71140, x71344);
  nand n71343(x71343, x71342, x71341);
  nand n71345(x71345, x15228, x614);
  nand n71346(x71346, x1, x86734);
  nand n71347(x71347, x71140, x71349);
  nand n71348(x71348, x71347, x71346);
  nand n71350(x71350, x15228, x615);
  nand n71351(x71351, x1, x86735);
  nand n71352(x71352, x71140, x71354);
  nand n71353(x71353, x71352, x71351);
  nand n71355(x71355, x15228, x616);
  nand n71356(x71356, x1, x86736);
  nand n71357(x71357, x71140, x71359);
  nand n71358(x71358, x71357, x71356);
  nand n71360(x71360, x15228, x617);
  nand n71361(x71361, x1, x86737);
  nand n71362(x71362, x71140, x71364);
  nand n71363(x71363, x71362, x71361);
  nand n71365(x71365, x15228, x618);
  nand n71366(x71366, x1, x86738);
  nand n71367(x71367, x71140, x71369);
  nand n71368(x71368, x71367, x71366);
  nand n71370(x71370, x15228, x619);
  nand n71371(x71371, x1, x86739);
  nand n71372(x71372, x71140, x71374);
  nand n71373(x71373, x71372, x71371);
  nand n71375(x71375, x15228, x620);
  nand n71376(x71376, x1, x86740);
  nand n71377(x71377, x71140, x71379);
  nand n71378(x71378, x71377, x71376);
  nand n71380(x71380, x15228, x621);
  nand n71381(x71381, x1, x86741);
  nand n71382(x71382, x71140, x71384);
  nand n71383(x71383, x71382, x71381);
  nand n71385(x71385, x15228, x622);
  nand n71386(x71386, x1, x86742);
  nand n71387(x71387, x71140, x71389);
  nand n71388(x71388, x71387, x71386);
  nand n71390(x71390, x15228, x623);
  nand n71391(x71391, x1, x86743);
  nand n71392(x71392, x71140, x71394);
  nand n71393(x71393, x71392, x71391);
  nand n71395(x71395, x15228, x624);
  nand n71396(x71396, x1, x86744);
  nand n71397(x71397, x71140, x71399);
  nand n71398(x71398, x71397, x71396);
  nand n71400(x71400, x15228, x625);
  nand n71401(x71401, x1, x86745);
  nand n71402(x71402, x71140, x71404);
  nand n71403(x71403, x71402, x71401);
  nand n71405(x71405, x15228, x626);
  nand n71406(x71406, x1, x86746);
  nand n71407(x71407, x71140, x71409);
  nand n71408(x71408, x71407, x71406);
  nand n71410(x71410, x15228, x627);
  nand n71411(x71411, x1, x86747);
  nand n71412(x71412, x71140, x71414);
  nand n71413(x71413, x71412, x71411);
  nand n71415(x71415, x15228, x628);
  nand n71416(x71416, x1, x86748);
  nand n71417(x71417, x71140, x71419);
  nand n71418(x71418, x71417, x71416);
  nand n71420(x71420, x15228, x629);
  nand n71421(x71421, x1, x86749);
  nand n71422(x71422, x71140, x71424);
  nand n71423(x71423, x71422, x71421);
  nand n71425(x71425, x15228, x630);
  nand n71426(x71426, x1, x86750);
  nand n71427(x71427, x71140, x71429);
  nand n71428(x71428, x71427, x71426);
  nand n71430(x71430, x15228, x631);
  nand n71431(x71431, x1, x86751);
  nand n71432(x71432, x71140, x71434);
  nand n71433(x71433, x71432, x71431);
  nand n71435(x71435, x15228, x632);
  nand n71436(x71436, x1, x86752);
  nand n71437(x71437, x71140, x71439);
  nand n71438(x71438, x71437, x71436);
  nand n71440(x71440, x15228, x633);
  nand n71441(x71441, x1, x86753);
  nand n71442(x71442, x71140, x71444);
  nand n71443(x71443, x71442, x71441);
  nand n71445(x71445, x15228, x0);
  nand n71446(x71446, x1, x86754);
  nand n71447(x71447, x71140, x71449);
  nand n71448(x71448, x71447, x71446);
  nand n71450(x71450, x15228, x58);
  nand n71451(x71451, x1, x86755);
  nand n71452(x71452, x71140, x71454);
  nand n71453(x71453, x71452, x71451);
  nand n71455(x71455, x15228, x59);
  nand n71456(x71456, x1, x86756);
  nand n71457(x71457, x71140, x71459);
  nand n71458(x71458, x71457, x71456);
  nand n71460(x71460, x15228, x60);
  nand n71461(x71461, x1, x86757);
  nand n71462(x71462, x71140, x71464);
  nand n71463(x71463, x71462, x71461);
  nand n71465(x71465, x15228, x61);
  nand n71466(x71466, x1, x86758);
  nand n71467(x71467, x71140, x71469);
  nand n71468(x71468, x71467, x71466);
  nand n71470(x71470, x15228, x62);
  nand n71471(x71471, x1, x86759);
  nand n71472(x71472, x71140, x71474);
  nand n71473(x71473, x71472, x71471);
  nand n71475(x71475, x15228, x63);
  nand n71476(x71476, x1, x86760);
  nand n71477(x71477, x71140, x71479);
  nand n71478(x71478, x71477, x71476);
  nand n71480(x71480, x71140, x71482);
  nand n71481(x71481, x71480, x71286);
  nand n71483(x71483, x71140, x71485);
  nand n71484(x71484, x71483, x71291);
  nand n71486(x71486, x15228, x93);
  nand n71487(x71487, x1, x86761);
  nand n71488(x71488, x71140, x71490);
  nand n71489(x71489, x71488, x71487);
  nand n71491(x71491, x15228, x296);
  nand n71492(x71492, x1, x86762);
  nand n71493(x71493, x71140, x71495);
  nand n71494(x71494, x71493, x71492);
  nand n71496(x71496, x15228, x300);
  nand n71497(x71497, x1, x86763);
  nand n71498(x71498, x71140, x71500);
  nand n71499(x71499, x71498, x71497);
  nand n71501(x71501, x15228, x304);
  nand n71502(x71502, x1, x86764);
  nand n71503(x71503, x71140, x71505);
  nand n71504(x71504, x71503, x71502);
  nand n71506(x71506, x15228, x308);
  nand n71507(x71507, x1, x86765);
  nand n71508(x71508, x71140, x71510);
  nand n71509(x71509, x71508, x71507);
  nand n71511(x71511, x15228, x312);
  nand n71512(x71512, x1, x86766);
  nand n71513(x71513, x71140, x71515);
  nand n71514(x71514, x71513, x71512);
  nand n71516(x71516, x15228, x316);
  nand n71517(x71517, x1, x86767);
  nand n71518(x71518, x71140, x71520);
  nand n71519(x71519, x71518, x71517);
  nand n71521(x71521, x15228, x320);
  nand n71522(x71522, x1, x86768);
  nand n71523(x71523, x71140, x71525);
  nand n71524(x71524, x71523, x71522);
  nand n71526(x71526, x15228, x324);
  nand n71527(x71527, x1, x86769);
  nand n71528(x71528, x71140, x71530);
  nand n71529(x71529, x71528, x71527);
  nand n71531(x71531, x15228, x328);
  nand n71532(x71532, x1, x86770);
  nand n71533(x71533, x71140, x71535);
  nand n71534(x71534, x71533, x71532);
  nand n71536(x71536, x15228, x332);
  nand n71537(x71537, x1, x86771);
  nand n71538(x71538, x71140, x71540);
  nand n71539(x71539, x71538, x71537);
  nand n71541(x71541, x15228, x336);
  nand n71542(x71542, x1, x86772);
  nand n71543(x71543, x71140, x71545);
  nand n71544(x71544, x71543, x71542);
  nand n71546(x71546, x15228, x340);
  nand n71547(x71547, x1, x86773);
  nand n71548(x71548, x71140, x71550);
  nand n71549(x71549, x71548, x71547);
  nand n71551(x71551, x15228, x344);
  nand n71552(x71552, x1, x86774);
  nand n71553(x71553, x71140, x71555);
  nand n71554(x71554, x71553, x71552);
  nand n71556(x71556, x15228, x348);
  nand n71557(x71557, x1, x86775);
  nand n71558(x71558, x71140, x71560);
  nand n71559(x71559, x71558, x71557);
  nand n71561(x71561, x15228, x352);
  nand n71562(x71562, x1, x86776);
  nand n71563(x71563, x71140, x71565);
  nand n71564(x71564, x71563, x71562);
  nand n71566(x71566, x15228, x356);
  nand n71567(x71567, x1, x86777);
  nand n71568(x71568, x71140, x71570);
  nand n71569(x71569, x71568, x71567);
  nand n71571(x71571, x15228, x360);
  nand n71572(x71572, x1, x86778);
  nand n71573(x71573, x71140, x71575);
  nand n71574(x71574, x71573, x71572);
  nand n71576(x71576, x15228, x364);
  nand n71577(x71577, x1, x86779);
  nand n71578(x71578, x71140, x71580);
  nand n71579(x71579, x71578, x71577);
  nand n71581(x71581, x15228, x368);
  nand n71582(x71582, x1, x86780);
  nand n71583(x71583, x71140, x71585);
  nand n71584(x71584, x71583, x71582);
  nand n71586(x71586, x15228, x372);
  nand n71587(x71587, x1, x86781);
  nand n71588(x71588, x71140, x71590);
  nand n71589(x71589, x71588, x71587);
  nand n71591(x71591, x15228, x376);
  nand n71592(x71592, x1, x86782);
  nand n71593(x71593, x71140, x71595);
  nand n71594(x71594, x71593, x71592);
  nand n71596(x71596, x15228, x380);
  nand n71597(x71597, x1, x86783);
  nand n71598(x71598, x71140, x71600);
  nand n71599(x71599, x71598, x71597);
  nand n71601(x71601, x15228, x384);
  nand n71602(x71602, x1, x86784);
  nand n71603(x71603, x71140, x71605);
  nand n71604(x71604, x71603, x71602);
  nand n71606(x71606, x15228, x388);
  nand n71607(x71607, x1, x86785);
  nand n71608(x71608, x71140, x71610);
  nand n71609(x71609, x71608, x71607);
  nand n71611(x71611, x15228, x392);
  nand n71612(x71612, x1, x86786);
  nand n71613(x71613, x71140, x71615);
  nand n71614(x71614, x71613, x71612);
  nand n71616(x71616, x15228, x396);
  nand n71617(x71617, x1, x86787);
  nand n71618(x71618, x71140, x71620);
  nand n71619(x71619, x71618, x71617);
  nand n71621(x71621, x15228, x400);
  nand n71622(x71622, x1, x86788);
  nand n71623(x71623, x71140, x71625);
  nand n71624(x71624, x71623, x71622);
  nand n71626(x71626, x15228, x404);
  nand n71627(x71627, x1, x86789);
  nand n71628(x71628, x71140, x71630);
  nand n71629(x71629, x71628, x71627);
  nand n71631(x71631, x15228, x408);
  nand n71632(x71632, x1, x86790);
  nand n71633(x71633, x71140, x71635);
  nand n71634(x71634, x71633, x71632);
  nand n71636(x71636, x71139, x71136);
  nand n71637(x71637, x71636, x71135);
  nand n71638(x71638, x71637, x71482);
  nand n71639(x71639, x71135, x86791);
  nand n71640(x71640, x68462, x71642);
  nand n71641(x71641, x71640, x71639);
  nand n71643(x71643, x71637, x71485);
  nand n71644(x71644, x71135, x86792);
  nand n71645(x71645, x68462, x71647);
  nand n71646(x71646, x71645, x71644);
  nand n71648(x71648, x71637, x71490);
  nand n71649(x71649, x71135, x86793);
  nand n71650(x71650, x68462, x71652);
  nand n71651(x71651, x71650, x71649);
  nand n71653(x71653, x71637, x71495);
  nand n71654(x71654, x71135, x86794);
  nand n71655(x71655, x68462, x71657);
  nand n71656(x71656, x71655, x71654);
  nand n71658(x71658, x71637, x71500);
  nand n71659(x71659, x71135, x86795);
  nand n71660(x71660, x68462, x71662);
  nand n71661(x71661, x71660, x71659);
  nand n71663(x71663, x71637, x71505);
  nand n71664(x71664, x71135, x86796);
  nand n71665(x71665, x68462, x71667);
  nand n71666(x71666, x71665, x71664);
  nand n71668(x71668, x71637, x71510);
  nand n71669(x71669, x71135, x86797);
  nand n71670(x71670, x68462, x71672);
  nand n71671(x71671, x71670, x71669);
  nand n71673(x71673, x71637, x71515);
  nand n71674(x71674, x71135, x86798);
  nand n71675(x71675, x68462, x71677);
  nand n71676(x71676, x71675, x71674);
  nand n71678(x71678, x71637, x71520);
  nand n71679(x71679, x71135, x86799);
  nand n71680(x71680, x68462, x71682);
  nand n71681(x71681, x71680, x71679);
  nand n71683(x71683, x71637, x71525);
  nand n71684(x71684, x71135, x86800);
  nand n71685(x71685, x68462, x71687);
  nand n71686(x71686, x71685, x71684);
  nand n71688(x71688, x71637, x71530);
  nand n71689(x71689, x71135, x86801);
  nand n71690(x71690, x68462, x71692);
  nand n71691(x71691, x71690, x71689);
  nand n71693(x71693, x71637, x71535);
  nand n71694(x71694, x71135, x86802);
  nand n71695(x71695, x68462, x71697);
  nand n71696(x71696, x71695, x71694);
  nand n71698(x71698, x71637, x71540);
  nand n71699(x71699, x71135, x86803);
  nand n71700(x71700, x68462, x71702);
  nand n71701(x71701, x71700, x71699);
  nand n71703(x71703, x71637, x71545);
  nand n71704(x71704, x71135, x86804);
  nand n71705(x71705, x68462, x71707);
  nand n71706(x71706, x71705, x71704);
  nand n71708(x71708, x71637, x71550);
  nand n71709(x71709, x71135, x86805);
  nand n71710(x71710, x68462, x71712);
  nand n71711(x71711, x71710, x71709);
  nand n71713(x71713, x71637, x71555);
  nand n71714(x71714, x71135, x86806);
  nand n71715(x71715, x68462, x71717);
  nand n71716(x71716, x71715, x71714);
  nand n71718(x71718, x71637, x71560);
  nand n71719(x71719, x71135, x86807);
  nand n71720(x71720, x68462, x71722);
  nand n71721(x71721, x71720, x71719);
  nand n71723(x71723, x71637, x71565);
  nand n71724(x71724, x71135, x86808);
  nand n71725(x71725, x68462, x71727);
  nand n71726(x71726, x71725, x71724);
  nand n71728(x71728, x71637, x71570);
  nand n71729(x71729, x71135, x86809);
  nand n71730(x71730, x68462, x71732);
  nand n71731(x71731, x71730, x71729);
  nand n71733(x71733, x71637, x71575);
  nand n71734(x71734, x71135, x86810);
  nand n71735(x71735, x68462, x71737);
  nand n71736(x71736, x71735, x71734);
  nand n71738(x71738, x71637, x71580);
  nand n71739(x71739, x71135, x86811);
  nand n71740(x71740, x68462, x71742);
  nand n71741(x71741, x71740, x71739);
  nand n71743(x71743, x71637, x71585);
  nand n71744(x71744, x71135, x86812);
  nand n71745(x71745, x68462, x71747);
  nand n71746(x71746, x71745, x71744);
  nand n71748(x71748, x71637, x71590);
  nand n71749(x71749, x71135, x86813);
  nand n71750(x71750, x68462, x71752);
  nand n71751(x71751, x71750, x71749);
  nand n71753(x71753, x71637, x71595);
  nand n71754(x71754, x71135, x86814);
  nand n71755(x71755, x68462, x71757);
  nand n71756(x71756, x71755, x71754);
  nand n71758(x71758, x71637, x71600);
  nand n71759(x71759, x71135, x86815);
  nand n71760(x71760, x68462, x71762);
  nand n71761(x71761, x71760, x71759);
  nand n71763(x71763, x71637, x71605);
  nand n71764(x71764, x71135, x86816);
  nand n71765(x71765, x68462, x71767);
  nand n71766(x71766, x71765, x71764);
  nand n71768(x71768, x71637, x71610);
  nand n71769(x71769, x71135, x86817);
  nand n71770(x71770, x68462, x71772);
  nand n71771(x71771, x71770, x71769);
  nand n71773(x71773, x71637, x71615);
  nand n71774(x71774, x71135, x86818);
  nand n71775(x71775, x68462, x71777);
  nand n71776(x71776, x71775, x71774);
  nand n71778(x71778, x71637, x71620);
  nand n71779(x71779, x71135, x86819);
  nand n71780(x71780, x68462, x71782);
  nand n71781(x71781, x71780, x71779);
  nand n71783(x71783, x71637, x71625);
  nand n71784(x71784, x71135, x86820);
  nand n71785(x71785, x68462, x71787);
  nand n71786(x71786, x71785, x71784);
  nand n71788(x71788, x71637, x71630);
  nand n71789(x71789, x71135, x86821);
  nand n71790(x71790, x68462, x71792);
  nand n71791(x71791, x71790, x71789);
  nand n71793(x71793, x71637, x71635);
  nand n71794(x71794, x71135, x86822);
  nand n71795(x71795, x68462, x71797);
  nand n71796(x71796, x71795, x71794);
  nand n71798(x71798, x71637, x15155);
  nand n71799(x71799, x71135, x86823);
  nand n71800(x71800, x68462, x71802);
  nand n71801(x71801, x71800, x71799);
  nand n71803(x71803, x71637, x15158);
  nand n71804(x71804, x71135, x86824);
  nand n71805(x71805, x68462, x71807);
  nand n71806(x71806, x71805, x71804);
  nand n71808(x71808, x71637, x15161);
  nand n71809(x71809, x71135, x86825);
  nand n71810(x71810, x68462, x71812);
  nand n71811(x71811, x71810, x71809);
  nand n71813(x71813, x71637, x15164);
  nand n71814(x71814, x71135, x86826);
  nand n71815(x71815, x68462, x71817);
  nand n71816(x71816, x71815, x71814);
  nand n71818(x71818, x71637, x15167);
  nand n71819(x71819, x71135, x86827);
  nand n71820(x71820, x68462, x71822);
  nand n71821(x71821, x71820, x71819);
  nand n71823(x71823, x71637, x15170);
  nand n71824(x71824, x71135, x86828);
  nand n71825(x71825, x68462, x71827);
  nand n71826(x71826, x71825, x71824);
  nand n71828(x71828, x71637, x15173);
  nand n71829(x71829, x71135, x86829);
  nand n71830(x71830, x68462, x71832);
  nand n71831(x71831, x71830, x71829);
  nand n71833(x71833, x71637, x15176);
  nand n71834(x71834, x71135, x86830);
  nand n71835(x71835, x68462, x71837);
  nand n71836(x71836, x71835, x71834);
  nand n71838(x71838, x71637, x15179);
  nand n71839(x71839, x71135, x86831);
  nand n71840(x71840, x68462, x71842);
  nand n71841(x71841, x71840, x71839);
  nand n71843(x71843, x71637, x15182);
  nand n71844(x71844, x71135, x86832);
  nand n71845(x71845, x68462, x71847);
  nand n71846(x71846, x71845, x71844);
  nand n71848(x71848, x71637, x15185);
  nand n71849(x71849, x71135, x86833);
  nand n71850(x71850, x68462, x71852);
  nand n71851(x71851, x71850, x71849);
  nand n71853(x71853, x71637, x15188);
  nand n71854(x71854, x71135, x86834);
  nand n71855(x71855, x68462, x71857);
  nand n71856(x71856, x71855, x71854);
  nand n71858(x71858, x71637, x15191);
  nand n71859(x71859, x71135, x86835);
  nand n71860(x71860, x68462, x71862);
  nand n71861(x71861, x71860, x71859);
  nand n71863(x71863, x71637, x15194);
  nand n71864(x71864, x71135, x86836);
  nand n71865(x71865, x68462, x71867);
  nand n71866(x71866, x71865, x71864);
  nand n71868(x71868, x71637, x15197);
  nand n71869(x71869, x71135, x86837);
  nand n71870(x71870, x68462, x71872);
  nand n71871(x71871, x71870, x71869);
  nand n71873(x71873, x71637, x15200);
  nand n71874(x71874, x71135, x86838);
  nand n71875(x71875, x68462, x71877);
  nand n71876(x71876, x71875, x71874);
  nand n71878(x71878, x71637, x15203);
  nand n71879(x71879, x71135, x86839);
  nand n71880(x71880, x68462, x71882);
  nand n71881(x71881, x71880, x71879);
  nand n71883(x71883, x71637, x15206);
  nand n71884(x71884, x71135, x86840);
  nand n71885(x71885, x68462, x71887);
  nand n71886(x71886, x71885, x71884);
  nand n71888(x71888, x71637, x15209);
  nand n71889(x71889, x71135, x86841);
  nand n71890(x71890, x68462, x71892);
  nand n71891(x71891, x71890, x71889);
  nand n71893(x71893, x71637, x15211);
  nand n71894(x71894, x71135, x86842);
  nand n71895(x71895, x68462, x71897);
  nand n71896(x71896, x71895, x71894);
  nand n71898(x71898, x71637, x15213);
  nand n71899(x71899, x71135, x86843);
  nand n71900(x71900, x68462, x71902);
  nand n71901(x71901, x71900, x71899);
  nand n71903(x71903, x71637, x15215);
  nand n71904(x71904, x71135, x86844);
  nand n71905(x71905, x68462, x71907);
  nand n71906(x71906, x71905, x71904);
  nand n71908(x71908, x68462, x71910);
  nand n71909(x71909, x71908, x71904);
  nand n71911(x71911, x68462, x71913);
  nand n71912(x71912, x71911, x71904);
  nand n71914(x71914, x68462, x71916);
  nand n71915(x71915, x71914, x71904);
  nand n71917(x71917, x68462, x71919);
  nand n71918(x71918, x71917, x71904);
  nand n71920(x71920, x68462, x71922);
  nand n71921(x71921, x71920, x71904);
  nand n71923(x71923, x68462, x71925);
  nand n71924(x71924, x71923, x71904);
  nand n71926(x71926, x68462, x71928);
  nand n71927(x71927, x71926, x71904);
  nand n71929(x71929, x68462, x71931);
  nand n71930(x71930, x71929, x71904);
  nand n71932(x71932, x68462, x71934);
  nand n71933(x71933, x71932, x71904);
  nand n71935(x71935, x68462, x71937);
  nand n71936(x71936, x71935, x71904);
  nand n71938(x71938, x71637, x15220);
  nand n71939(x71939, x71135, x86845);
  nand n71940(x71940, x68462, x71942);
  nand n71941(x71941, x71940, x71939);
  nand n71943(x71943, x71637, x71454);
  nand n71944(x71944, x71135, x86846);
  nand n71945(x71945, x68462, x71947);
  nand n71946(x71946, x71945, x71944);
  nand n71948(x71948, x71637, x71459);
  nand n71949(x71949, x71135, x86847);
  nand n71950(x71950, x68462, x71952);
  nand n71951(x71951, x71950, x71949);
  nand n71953(x71953, x71637, x71464);
  nand n71954(x71954, x71135, x86848);
  nand n71955(x71955, x68462, x71957);
  nand n71956(x71956, x71955, x71954);
  nand n71958(x71958, x71637, x71469);
  nand n71959(x71959, x71135, x86849);
  nand n71960(x71960, x68462, x71962);
  nand n71961(x71961, x71960, x71959);
  nand n71963(x71963, x71637, x71474);
  nand n71964(x71964, x71135, x86850);
  nand n71965(x71965, x68462, x71967);
  nand n71966(x71966, x71965, x71964);
  nand n71968(x71968, x71637, x71479);
  nand n71969(x71969, x71135, x86851);
  nand n71970(x71970, x68462, x71972);
  nand n71971(x71971, x71970, x71969);
  nand n71973(x71973, x71637, x71245);
  nand n71974(x71974, x71135, x86852);
  nand n71975(x71975, x68462, x71977);
  nand n71976(x71976, x71975, x71974);
  nand n71978(x71978, x71637, x71250);
  nand n71979(x71979, x71135, x86853);
  nand n71980(x71980, x68462, x71982);
  nand n71981(x71981, x71980, x71979);
  nand n71983(x71983, x71637, x71255);
  nand n71984(x71984, x71135, x86854);
  nand n71985(x71985, x68462, x71987);
  nand n71986(x71986, x71985, x71984);
  nand n71988(x71988, x71637, x71260);
  nand n71989(x71989, x71135, x86855);
  nand n71990(x71990, x68462, x71992);
  nand n71991(x71991, x71990, x71989);
  nand n71993(x71993, x71637, x71265);
  nand n71994(x71994, x71135, x86856);
  nand n71995(x71995, x68462, x71997);
  nand n71996(x71996, x71995, x71994);
  nand n71998(x71998, x71637, x71270);
  nand n71999(x71999, x71135, x86857);
  nand n72000(x72000, x68462, x72002);
  nand n72001(x72001, x72000, x71999);
  nand n72003(x72003, x71637, x71230);
  nand n72004(x72004, x71135, x86858);
  nand n72005(x72005, x68462, x72007);
  nand n72006(x72006, x72005, x72004);
  nand n72008(x72008, x71637, x71235);
  nand n72009(x72009, x71135, x86859);
  nand n72010(x72010, x68462, x72012);
  nand n72011(x72011, x72010, x72009);
  nand n72013(x72013, x71637, x71240);
  nand n72014(x72014, x71135, x86860);
  nand n72015(x72015, x68462, x72017);
  nand n72016(x72016, x72015, x72014);
  nand n72018(x72018, x71637, x1715);
  nand n72019(x72019, x71135, x86861);
  nand n72020(x72020, x68462, x72022);
  nand n72021(x72021, x72020, x72019);
  nand n72023(x72023, x71637, x1693);
  nand n72024(x72024, x71135, x86862);
  nand n72025(x72025, x68462, x72027);
  nand n72026(x72026, x72025, x72024);
  nand n72028(x72028, x71637, x1695);
  nand n72029(x72029, x71135, x86863);
  nand n72030(x72030, x68462, x72032);
  nand n72031(x72031, x72030, x72029);
  nand n72033(x72033, x71637, x1697);
  nand n72034(x72034, x71135, x86864);
  nand n72035(x72035, x68462, x72037);
  nand n72036(x72036, x72035, x72034);
  nand n72038(x72038, x71637, x1699);
  nand n72039(x72039, x71135, x86865);
  nand n72040(x72040, x68462, x72042);
  nand n72041(x72041, x72040, x72039);
  nand n72043(x72043, x71637, x6503);
  nand n72044(x72044, x71135, x86866);
  nand n72045(x72045, x68462, x72047);
  nand n72046(x72046, x72045, x72044);
  nand n72048(x72048, x71637, x6524);
  nand n72049(x72049, x71135, x86867);
  nand n72050(x72050, x68462, x72052);
  nand n72051(x72051, x72050, x72049);
  nand n72053(x72053, x71637, x6545);
  nand n72054(x72054, x71135, x86868);
  nand n72055(x72055, x68462, x72057);
  nand n72056(x72056, x72055, x72054);
  nand n72058(x72058, x71637, x6566);
  nand n72059(x72059, x71135, x86869);
  nand n72060(x72060, x68462, x72062);
  nand n72061(x72061, x72060, x72059);
  nand n72063(x72063, x71637, x6587);
  nand n72064(x72064, x71135, x86870);
  nand n72065(x72065, x68462, x72067);
  nand n72066(x72066, x72065, x72064);
  nand n72068(x72068, x71637, x6608);
  nand n72069(x72069, x71135, x86871);
  nand n72070(x72070, x68462, x72072);
  nand n72071(x72071, x72070, x72069);
  nand n72073(x72073, x71637, x6629);
  nand n72074(x72074, x71135, x86872);
  nand n72075(x72075, x68462, x72077);
  nand n72076(x72076, x72075, x72074);
  nand n72078(x72078, x71637, x6650);
  nand n72079(x72079, x71135, x86873);
  nand n72080(x72080, x68462, x72082);
  nand n72081(x72081, x72080, x72079);
  nand n72083(x72083, x71637, x6671);
  nand n72084(x72084, x71135, x86874);
  nand n72085(x72085, x68462, x72087);
  nand n72086(x72086, x72085, x72084);
  nand n72088(x72088, x71637, x6692);
  nand n72089(x72089, x71135, x86875);
  nand n72090(x72090, x68462, x72092);
  nand n72091(x72091, x72090, x72089);
  nand n72093(x72093, x71637, x6713);
  nand n72094(x72094, x71135, x86876);
  nand n72095(x72095, x68462, x72097);
  nand n72096(x72096, x72095, x72094);
  nand n72098(x72098, x71637, x6734);
  nand n72099(x72099, x71135, x86877);
  nand n72100(x72100, x68462, x72102);
  nand n72101(x72101, x72100, x72099);
  nand n72103(x72103, x71637, x6755);
  nand n72104(x72104, x71135, x86878);
  nand n72105(x72105, x68462, x72107);
  nand n72106(x72106, x72105, x72104);
  nand n72108(x72108, x71637, x6776);
  nand n72109(x72109, x71135, x86879);
  nand n72110(x72110, x68462, x72112);
  nand n72111(x72111, x72110, x72109);
  nand n72113(x72113, x71637, x6797);
  nand n72114(x72114, x71135, x86880);
  nand n72115(x72115, x68462, x72117);
  nand n72116(x72116, x72115, x72114);
  nand n72118(x72118, x71637, x6818);
  nand n72119(x72119, x71135, x86881);
  nand n72120(x72120, x68462, x72122);
  nand n72121(x72121, x72120, x72119);
  nand n72123(x72123, x71637, x6839);
  nand n72124(x72124, x71135, x86882);
  nand n72125(x72125, x68462, x72127);
  nand n72126(x72126, x72125, x72124);
  nand n72128(x72128, x71637, x6860);
  nand n72129(x72129, x71135, x86883);
  nand n72130(x72130, x68462, x72132);
  nand n72131(x72131, x72130, x72129);
  nand n72133(x72133, x71637, x6881);
  nand n72134(x72134, x71135, x86884);
  nand n72135(x72135, x68462, x72137);
  nand n72136(x72136, x72135, x72134);
  nand n72138(x72138, x71637, x6902);
  nand n72139(x72139, x71135, x86885);
  nand n72140(x72140, x68462, x72142);
  nand n72141(x72141, x72140, x72139);
  nand n72143(x72143, x71637, x6923);
  nand n72144(x72144, x71135, x86886);
  nand n72145(x72145, x68462, x72147);
  nand n72146(x72146, x72145, x72144);
  nand n72148(x72148, x71637, x6944);
  nand n72149(x72149, x71135, x86887);
  nand n72150(x72150, x68462, x72152);
  nand n72151(x72151, x72150, x72149);
  nand n72153(x72153, x71637, x6965);
  nand n72154(x72154, x71135, x86888);
  nand n72155(x72155, x68462, x72157);
  nand n72156(x72156, x72155, x72154);
  nand n72158(x72158, x71637, x6986);
  nand n72159(x72159, x71135, x86889);
  nand n72160(x72160, x68462, x72162);
  nand n72161(x72161, x72160, x72159);
  nand n72163(x72163, x71637, x7007);
  nand n72164(x72164, x71135, x86890);
  nand n72165(x72165, x68462, x72167);
  nand n72166(x72166, x72165, x72164);
  nand n72168(x72168, x71637, x7028);
  nand n72169(x72169, x71135, x86891);
  nand n72170(x72170, x68462, x72172);
  nand n72171(x72171, x72170, x72169);
  nand n72173(x72173, x71637, x7049);
  nand n72174(x72174, x71135, x86892);
  nand n72175(x72175, x68462, x72177);
  nand n72176(x72176, x72175, x72174);
  nand n72178(x72178, x71637, x7070);
  nand n72179(x72179, x71135, x86893);
  nand n72180(x72180, x68462, x72182);
  nand n72181(x72181, x72180, x72179);
  nand n72183(x72183, x71637, x7091);
  nand n72184(x72184, x71135, x86894);
  nand n72185(x72185, x68462, x72187);
  nand n72186(x72186, x72185, x72184);
  nand n72188(x72188, x71637, x7112);
  nand n72189(x72189, x71135, x86895);
  nand n72190(x72190, x68462, x72192);
  nand n72191(x72191, x72190, x72189);
  nand n72193(x72193, x71637, x7133);
  nand n72194(x72194, x71135, x86896);
  nand n72195(x72195, x68462, x72197);
  nand n72196(x72196, x72195, x72194);
  nand n72198(x72198, x71637, x7154);
  nand n72199(x72199, x71135, x86897);
  nand n72200(x72200, x68462, x72202);
  nand n72201(x72201, x72200, x72199);
  nand n72203(x72203, x71637, x7178);
  nand n72204(x72204, x71135, x86898);
  nand n72205(x72205, x68462, x72207);
  nand n72206(x72206, x72205, x72204);
  nand n72208(x72208, x71637, x7199);
  nand n72209(x72209, x71135, x86899);
  nand n72210(x72210, x68462, x72212);
  nand n72211(x72211, x72210, x72209);
  nand n72213(x72213, x71637, x7220);
  nand n72214(x72214, x71135, x86900);
  nand n72215(x72215, x68462, x72217);
  nand n72216(x72216, x72215, x72214);
  nand n72218(x72218, x71637, x7241);
  nand n72219(x72219, x71135, x86901);
  nand n72220(x72220, x68462, x72222);
  nand n72221(x72221, x72220, x72219);
  nand n72223(x72223, x71637, x7262);
  nand n72224(x72224, x71135, x86902);
  nand n72225(x72225, x68462, x72227);
  nand n72226(x72226, x72225, x72224);
  nand n72228(x72228, x71637, x7283);
  nand n72229(x72229, x71135, x86903);
  nand n72230(x72230, x68462, x72232);
  nand n72231(x72231, x72230, x72229);
  nand n72233(x72233, x71637, x7304);
  nand n72234(x72234, x71135, x86904);
  nand n72235(x72235, x68462, x72237);
  nand n72236(x72236, x72235, x72234);
  nand n72238(x72238, x71637, x7325);
  nand n72239(x72239, x71135, x86905);
  nand n72240(x72240, x68462, x72242);
  nand n72241(x72241, x72240, x72239);
  nand n72243(x72243, x71637, x7346);
  nand n72244(x72244, x71135, x86906);
  nand n72245(x72245, x68462, x72247);
  nand n72246(x72246, x72245, x72244);
  nand n72248(x72248, x71637, x7367);
  nand n72249(x72249, x71135, x86907);
  nand n72250(x72250, x68462, x72252);
  nand n72251(x72251, x72250, x72249);
  nand n72253(x72253, x71637, x7388);
  nand n72254(x72254, x71135, x86908);
  nand n72255(x72255, x68462, x72257);
  nand n72256(x72256, x72255, x72254);
  nand n72258(x72258, x71637, x7409);
  nand n72259(x72259, x71135, x86909);
  nand n72260(x72260, x68462, x72262);
  nand n72261(x72261, x72260, x72259);
  nand n72263(x72263, x71637, x7430);
  nand n72264(x72264, x71135, x86910);
  nand n72265(x72265, x68462, x72267);
  nand n72266(x72266, x72265, x72264);
  nand n72268(x72268, x71637, x7451);
  nand n72269(x72269, x71135, x86911);
  nand n72270(x72270, x68462, x72272);
  nand n72271(x72271, x72270, x72269);
  nand n72273(x72273, x71637, x7472);
  nand n72274(x72274, x71135, x86912);
  nand n72275(x72275, x68462, x72277);
  nand n72276(x72276, x72275, x72274);
  nand n72278(x72278, x71637, x7493);
  nand n72279(x72279, x71135, x86913);
  nand n72280(x72280, x68462, x72282);
  nand n72281(x72281, x72280, x72279);
  nand n72283(x72283, x71637, x7514);
  nand n72284(x72284, x71135, x86914);
  nand n72285(x72285, x68462, x72287);
  nand n72286(x72286, x72285, x72284);
  nand n72288(x72288, x71637, x7535);
  nand n72289(x72289, x71135, x86915);
  nand n72290(x72290, x68462, x72292);
  nand n72291(x72291, x72290, x72289);
  nand n72293(x72293, x71637, x7556);
  nand n72294(x72294, x71135, x86916);
  nand n72295(x72295, x68462, x72297);
  nand n72296(x72296, x72295, x72294);
  nand n72298(x72298, x71637, x7577);
  nand n72299(x72299, x71135, x86917);
  nand n72300(x72300, x68462, x72302);
  nand n72301(x72301, x72300, x72299);
  nand n72303(x72303, x71637, x7598);
  nand n72304(x72304, x71135, x86918);
  nand n72305(x72305, x68462, x72307);
  nand n72306(x72306, x72305, x72304);
  nand n72308(x72308, x71637, x7619);
  nand n72309(x72309, x71135, x86919);
  nand n72310(x72310, x68462, x72312);
  nand n72311(x72311, x72310, x72309);
  nand n72313(x72313, x71637, x7640);
  nand n72314(x72314, x71135, x86920);
  nand n72315(x72315, x68462, x72317);
  nand n72316(x72316, x72315, x72314);
  nand n72318(x72318, x71637, x7661);
  nand n72319(x72319, x71135, x86921);
  nand n72320(x72320, x68462, x72322);
  nand n72321(x72321, x72320, x72319);
  nand n72323(x72323, x71637, x7682);
  nand n72324(x72324, x71135, x86922);
  nand n72325(x72325, x68462, x72327);
  nand n72326(x72326, x72325, x72324);
  nand n72328(x72328, x71637, x7703);
  nand n72329(x72329, x71135, x86923);
  nand n72330(x72330, x68462, x72332);
  nand n72331(x72331, x72330, x72329);
  nand n72333(x72333, x71637, x7724);
  nand n72334(x72334, x71135, x86924);
  nand n72335(x72335, x68462, x72337);
  nand n72336(x72336, x72335, x72334);
  nand n72338(x72338, x71637, x7745);
  nand n72339(x72339, x71135, x86925);
  nand n72340(x72340, x68462, x72342);
  nand n72341(x72341, x72340, x72339);
  nand n72343(x72343, x71637, x7766);
  nand n72344(x72344, x71135, x86926);
  nand n72345(x72345, x68462, x72347);
  nand n72346(x72346, x72345, x72344);
  nand n72348(x72348, x71637, x7787);
  nand n72349(x72349, x71135, x86927);
  nand n72350(x72350, x68462, x72352);
  nand n72351(x72351, x72350, x72349);
  nand n72353(x72353, x71637, x7808);
  nand n72354(x72354, x71135, x86928);
  nand n72355(x72355, x68462, x72357);
  nand n72356(x72356, x72355, x72354);
  nand n72358(x72358, x71637, x7829);
  nand n72359(x72359, x71135, x86929);
  nand n72360(x72360, x68462, x72362);
  nand n72361(x72361, x72360, x72359);
  nand n72363(x72363, x71637, x7850);
  nand n72364(x72364, x71135, x86930);
  nand n72365(x72365, x68462, x72367);
  nand n72366(x72366, x72365, x72364);
  nand n72368(x72368, x71637, x7871);
  nand n72369(x72369, x71135, x86931);
  nand n72370(x72370, x68462, x72372);
  nand n72371(x72371, x72370, x72369);
  nand n72373(x72373, x71637, x7892);
  nand n72374(x72374, x71135, x86932);
  nand n72375(x72375, x68462, x72377);
  nand n72376(x72376, x72375, x72374);
  nand n72378(x72378, x71637, x7913);
  nand n72379(x72379, x71135, x86933);
  nand n72380(x72380, x68462, x72382);
  nand n72381(x72381, x72380, x72379);
  nand n72383(x72383, x71637, x7934);
  nand n72384(x72384, x71135, x86934);
  nand n72385(x72385, x68462, x72387);
  nand n72386(x72386, x72385, x72384);
  nand n72388(x72388, x71637, x7955);
  nand n72389(x72389, x71135, x86935);
  nand n72390(x72390, x68462, x72392);
  nand n72391(x72391, x72390, x72389);
  nand n72393(x72393, x71637, x7976);
  nand n72394(x72394, x71135, x86936);
  nand n72395(x72395, x68462, x72397);
  nand n72396(x72396, x72395, x72394);
  nand n72398(x72398, x71637, x7997);
  nand n72399(x72399, x71135, x86937);
  nand n72400(x72400, x68462, x72402);
  nand n72401(x72401, x72400, x72399);
  nand n72403(x72403, x71637, x8018);
  nand n72404(x72404, x71135, x86938);
  nand n72405(x72405, x68462, x72407);
  nand n72406(x72406, x72405, x72404);
  nand n72408(x72408, x71637, x8039);
  nand n72409(x72409, x71135, x86939);
  nand n72410(x72410, x68462, x72412);
  nand n72411(x72411, x72410, x72409);
  nand n72413(x72413, x71637, x8060);
  nand n72414(x72414, x71135, x86940);
  nand n72415(x72415, x68462, x72417);
  nand n72416(x72416, x72415, x72414);
  nand n72418(x72418, x71637, x8081);
  nand n72419(x72419, x71135, x86941);
  nand n72420(x72420, x68462, x72422);
  nand n72421(x72421, x72420, x72419);
  nand n72423(x72423, x71637, x8102);
  nand n72424(x72424, x71135, x86942);
  nand n72425(x72425, x68462, x72427);
  nand n72426(x72426, x72425, x72424);
  nand n72428(x72428, x71637, x8123);
  nand n72429(x72429, x71135, x86943);
  nand n72430(x72430, x68462, x72432);
  nand n72431(x72431, x72430, x72429);
  nand n72433(x72433, x71637, x8144);
  nand n72434(x72434, x71135, x86944);
  nand n72435(x72435, x68462, x72437);
  nand n72436(x72436, x72435, x72434);
  nand n72438(x72438, x71637, x8165);
  nand n72439(x72439, x71135, x86945);
  nand n72440(x72440, x68462, x72442);
  nand n72441(x72441, x72440, x72439);
  nand n72443(x72443, x71637, x8186);
  nand n72444(x72444, x71135, x86946);
  nand n72445(x72445, x68462, x72447);
  nand n72446(x72446, x72445, x72444);
  nand n72448(x72448, x71637, x8207);
  nand n72449(x72449, x71135, x86947);
  nand n72450(x72450, x68462, x72452);
  nand n72451(x72451, x72450, x72449);
  nand n72453(x72453, x71637, x8228);
  nand n72454(x72454, x71135, x86948);
  nand n72455(x72455, x68462, x72457);
  nand n72456(x72456, x72455, x72454);
  nand n72458(x72458, x71637, x8249);
  nand n72459(x72459, x71135, x86949);
  nand n72460(x72460, x68462, x72462);
  nand n72461(x72461, x72460, x72459);
  nand n72463(x72463, x71637, x8270);
  nand n72464(x72464, x71135, x86950);
  nand n72465(x72465, x68462, x72467);
  nand n72466(x72466, x72465, x72464);
  nand n72468(x72468, x71637, x8291);
  nand n72469(x72469, x71135, x86951);
  nand n72470(x72470, x68462, x72472);
  nand n72471(x72471, x72470, x72469);
  nand n72473(x72473, x71637, x8312);
  nand n72474(x72474, x71135, x86952);
  nand n72475(x72475, x68462, x72477);
  nand n72476(x72476, x72475, x72474);
  nand n72478(x72478, x71637, x8333);
  nand n72479(x72479, x71135, x86953);
  nand n72480(x72480, x68462, x72482);
  nand n72481(x72481, x72480, x72479);
  nand n72483(x72483, x71637, x8354);
  nand n72484(x72484, x71135, x86954);
  nand n72485(x72485, x68462, x72487);
  nand n72486(x72486, x72485, x72484);
  nand n72488(x72488, x71637, x8375);
  nand n72489(x72489, x71135, x86955);
  nand n72490(x72490, x68462, x72492);
  nand n72491(x72491, x72490, x72489);
  nand n72493(x72493, x71637, x8396);
  nand n72494(x72494, x71135, x86956);
  nand n72495(x72495, x68462, x72497);
  nand n72496(x72496, x72495, x72494);
  nand n72498(x72498, x71637, x8417);
  nand n72499(x72499, x71135, x86957);
  nand n72500(x72500, x68462, x72502);
  nand n72501(x72501, x72500, x72499);
  nand n72503(x72503, x71637, x8438);
  nand n72504(x72504, x71135, x86958);
  nand n72505(x72505, x68462, x72507);
  nand n72506(x72506, x72505, x72504);
  nand n72508(x72508, x71637, x8459);
  nand n72509(x72509, x71135, x86959);
  nand n72510(x72510, x68462, x72512);
  nand n72511(x72511, x72510, x72509);
  nand n72513(x72513, x71637, x8480);
  nand n72514(x72514, x71135, x86960);
  nand n72515(x72515, x68462, x72517);
  nand n72516(x72516, x72515, x72514);
  nand n72518(x72518, x71637, x8501);
  nand n72519(x72519, x71135, x86961);
  nand n72520(x72520, x68462, x72522);
  nand n72521(x72521, x72520, x72519);
  nand n72523(x72523, x71637, x1446);
  nand n72524(x72524, x71135, x86962);
  nand n72525(x72525, x68462, x72527);
  nand n72526(x72526, x72525, x72524);
  nand n72528(x72528, x71637, x1470);
  nand n72529(x72529, x71135, x86963);
  nand n72530(x72530, x68462, x72532);
  nand n72531(x72531, x72530, x72529);
  nand n72533(x72533, x71637, x8522);
  nand n72534(x72534, x71135, x86964);
  nand n72535(x72535, x68462, x72537);
  nand n72536(x72536, x72535, x72534);
  nand n72538(x72538, x71637, x8543);
  nand n72539(x72539, x71135, x86965);
  nand n72540(x72540, x68462, x72542);
  nand n72541(x72541, x72540, x72539);
  nand n72543(x72543, x71637, x8564);
  nand n72544(x72544, x71135, x86966);
  nand n72545(x72545, x68462, x72547);
  nand n72546(x72546, x72545, x72544);
  nand n72548(x72548, x71637, x8585);
  nand n72549(x72549, x71135, x86967);
  nand n72550(x72550, x68462, x72552);
  nand n72551(x72551, x72550, x72549);
  nand n72553(x72553, x71637, x8606);
  nand n72554(x72554, x71135, x86968);
  nand n72555(x72555, x68462, x72557);
  nand n72556(x72556, x72555, x72554);
  nand n72558(x72558, x71637, x8627);
  nand n72559(x72559, x71135, x86969);
  nand n72560(x72560, x68462, x72562);
  nand n72561(x72561, x72560, x72559);
  nand n72563(x72563, x71637, x8648);
  nand n72564(x72564, x71135, x86970);
  nand n72565(x72565, x68462, x72567);
  nand n72566(x72566, x72565, x72564);
  nand n72568(x72568, x71637, x8669);
  nand n72569(x72569, x71135, x86971);
  nand n72570(x72570, x68462, x72572);
  nand n72571(x72571, x72570, x72569);
  nand n72573(x72573, x71637, x8690);
  nand n72574(x72574, x71135, x86972);
  nand n72575(x72575, x68462, x72577);
  nand n72576(x72576, x72575, x72574);
  nand n72578(x72578, x71637, x8711);
  nand n72579(x72579, x71135, x86973);
  nand n72580(x72580, x68462, x72582);
  nand n72581(x72581, x72580, x72579);
  nand n72583(x72583, x71637, x8732);
  nand n72584(x72584, x71135, x86974);
  nand n72585(x72585, x68462, x72587);
  nand n72586(x72586, x72585, x72584);
  nand n72588(x72588, x71637, x8753);
  nand n72589(x72589, x71135, x86975);
  nand n72590(x72590, x68462, x72592);
  nand n72591(x72591, x72590, x72589);
  nand n72593(x72593, x71637, x8774);
  nand n72594(x72594, x71135, x86976);
  nand n72595(x72595, x68462, x72597);
  nand n72596(x72596, x72595, x72594);
  nand n72598(x72598, x71637, x8795);
  nand n72599(x72599, x71135, x86977);
  nand n72600(x72600, x68462, x72602);
  nand n72601(x72601, x72600, x72599);
  nand n72603(x72603, x71637, x8816);
  nand n72604(x72604, x71135, x86978);
  nand n72605(x72605, x68462, x72607);
  nand n72606(x72606, x72605, x72604);
  nand n72608(x72608, x71637, x8837);
  nand n72609(x72609, x71135, x86979);
  nand n72610(x72610, x68462, x72612);
  nand n72611(x72611, x72610, x72609);
  nand n72613(x72613, x71637, x8858);
  nand n72614(x72614, x71135, x86980);
  nand n72615(x72615, x68462, x72617);
  nand n72616(x72616, x72615, x72614);
  nand n72618(x72618, x71637, x8879);
  nand n72619(x72619, x71135, x86981);
  nand n72620(x72620, x68462, x72622);
  nand n72621(x72621, x72620, x72619);
  nand n72623(x72623, x71637, x8900);
  nand n72624(x72624, x71135, x86982);
  nand n72625(x72625, x68462, x72627);
  nand n72626(x72626, x72625, x72624);
  nand n72628(x72628, x71637, x8921);
  nand n72629(x72629, x71135, x86983);
  nand n72630(x72630, x68462, x72632);
  nand n72631(x72631, x72630, x72629);
  nand n72633(x72633, x71637, x8942);
  nand n72634(x72634, x71135, x86984);
  nand n72635(x72635, x68462, x72637);
  nand n72636(x72636, x72635, x72634);
  nand n72638(x72638, x71637, x8963);
  nand n72639(x72639, x71135, x86985);
  nand n72640(x72640, x68462, x72642);
  nand n72641(x72641, x72640, x72639);
  nand n72643(x72643, x71637, x8984);
  nand n72644(x72644, x71135, x86986);
  nand n72645(x72645, x68462, x72647);
  nand n72646(x72646, x72645, x72644);
  nand n72648(x72648, x71637, x9005);
  nand n72649(x72649, x71135, x86987);
  nand n72650(x72650, x68462, x72652);
  nand n72651(x72651, x72650, x72649);
  nand n72653(x72653, x71637, x9026);
  nand n72654(x72654, x71135, x86988);
  nand n72655(x72655, x68462, x72657);
  nand n72656(x72656, x72655, x72654);
  nand n72658(x72658, x71637, x9047);
  nand n72659(x72659, x71135, x86989);
  nand n72660(x72660, x68462, x72662);
  nand n72661(x72661, x72660, x72659);
  nand n72663(x72663, x71637, x9068);
  nand n72664(x72664, x71135, x86990);
  nand n72665(x72665, x68462, x72667);
  nand n72666(x72666, x72665, x72664);
  nand n72668(x72668, x71637, x9089);
  nand n72669(x72669, x71135, x86991);
  nand n72670(x72670, x68462, x72672);
  nand n72671(x72671, x72670, x72669);
  nand n72673(x72673, x71637, x9110);
  nand n72674(x72674, x71135, x86992);
  nand n72675(x72675, x68462, x72677);
  nand n72676(x72676, x72675, x72674);
  nand n72678(x72678, x71637, x9131);
  nand n72679(x72679, x71135, x86993);
  nand n72680(x72680, x68462, x72682);
  nand n72681(x72681, x72680, x72679);
  nand n72683(x72683, x71637, x9152);
  nand n72684(x72684, x71135, x86994);
  nand n72685(x72685, x68462, x72687);
  nand n72686(x72686, x72685, x72684);
  nand n72688(x72688, x71637, x9173);
  nand n72689(x72689, x71135, x86995);
  nand n72690(x72690, x68462, x72692);
  nand n72691(x72691, x72690, x72689);
  nand n72693(x72693, x71637, x9194);
  nand n72694(x72694, x71135, x86996);
  nand n72695(x72695, x68462, x72697);
  nand n72696(x72696, x72695, x72694);
  nand n72698(x72698, x71637, x9215);
  nand n72699(x72699, x71135, x86997);
  nand n72700(x72700, x68462, x72702);
  nand n72701(x72701, x72700, x72699);
  nand n72703(x72703, x71637, x9236);
  nand n72704(x72704, x71135, x86998);
  nand n72705(x72705, x68462, x72707);
  nand n72706(x72706, x72705, x72704);
  nand n72708(x72708, x71637, x9257);
  nand n72709(x72709, x71135, x86999);
  nand n72710(x72710, x68462, x72712);
  nand n72711(x72711, x72710, x72709);
  nand n72713(x72713, x71637, x9278);
  nand n72714(x72714, x71135, x87000);
  nand n72715(x72715, x68462, x72717);
  nand n72716(x72716, x72715, x72714);
  nand n72718(x72718, x71637, x9299);
  nand n72719(x72719, x71135, x87001);
  nand n72720(x72720, x68462, x72722);
  nand n72721(x72721, x72720, x72719);
  nand n72723(x72723, x71637, x9320);
  nand n72724(x72724, x71135, x87002);
  nand n72725(x72725, x68462, x72727);
  nand n72726(x72726, x72725, x72724);
  nand n72728(x72728, x71637, x9341);
  nand n72729(x72729, x71135, x87003);
  nand n72730(x72730, x68462, x72732);
  nand n72731(x72731, x72730, x72729);
  nand n72733(x72733, x71637, x9362);
  nand n72734(x72734, x71135, x87004);
  nand n72735(x72735, x68462, x72737);
  nand n72736(x72736, x72735, x72734);
  nand n72738(x72738, x71637, x9383);
  nand n72739(x72739, x71135, x87005);
  nand n72740(x72740, x68462, x72742);
  nand n72741(x72741, x72740, x72739);
  nand n72743(x72743, x71637, x9404);
  nand n72744(x72744, x71135, x87006);
  nand n72745(x72745, x68462, x72747);
  nand n72746(x72746, x72745, x72744);
  nand n72748(x72748, x71637, x9425);
  nand n72749(x72749, x71135, x87007);
  nand n72750(x72750, x68462, x72752);
  nand n72751(x72751, x72750, x72749);
  nand n72753(x72753, x71637, x9446);
  nand n72754(x72754, x71135, x87008);
  nand n72755(x72755, x68462, x72757);
  nand n72756(x72756, x72755, x72754);
  nand n72758(x72758, x71637, x9467);
  nand n72759(x72759, x71135, x87009);
  nand n72760(x72760, x68462, x72762);
  nand n72761(x72761, x72760, x72759);
  nand n72763(x72763, x71637, x9488);
  nand n72764(x72764, x71135, x87010);
  nand n72765(x72765, x68462, x72767);
  nand n72766(x72766, x72765, x72764);
  nand n72768(x72768, x71637, x9509);
  nand n72769(x72769, x71135, x87011);
  nand n72770(x72770, x68462, x72772);
  nand n72771(x72771, x72770, x72769);
  nand n72773(x72773, x71637, x9530);
  nand n72774(x72774, x71135, x87012);
  nand n72775(x72775, x68462, x72777);
  nand n72776(x72776, x72775, x72774);
  nand n72778(x72778, x71637, x9551);
  nand n72779(x72779, x71135, x87013);
  nand n72780(x72780, x68462, x72782);
  nand n72781(x72781, x72780, x72779);
  nand n72783(x72783, x71637, x9572);
  nand n72784(x72784, x71135, x87014);
  nand n72785(x72785, x68462, x72787);
  nand n72786(x72786, x72785, x72784);
  nand n72788(x72788, x71637, x9593);
  nand n72789(x72789, x71135, x87015);
  nand n72790(x72790, x68462, x72792);
  nand n72791(x72791, x72790, x72789);
  nand n72793(x72793, x71637, x9614);
  nand n72794(x72794, x71135, x87016);
  nand n72795(x72795, x68462, x72797);
  nand n72796(x72796, x72795, x72794);
  nand n72798(x72798, x71637, x9635);
  nand n72799(x72799, x71135, x87017);
  nand n72800(x72800, x68462, x72802);
  nand n72801(x72801, x72800, x72799);
  nand n72803(x72803, x71637, x9656);
  nand n72804(x72804, x71135, x87018);
  nand n72805(x72805, x68462, x72807);
  nand n72806(x72806, x72805, x72804);
  nand n72808(x72808, x71637, x9677);
  nand n72809(x72809, x71135, x87019);
  nand n72810(x72810, x68462, x72812);
  nand n72811(x72811, x72810, x72809);
  nand n72813(x72813, x71637, x9698);
  nand n72814(x72814, x71135, x87020);
  nand n72815(x72815, x68462, x72817);
  nand n72816(x72816, x72815, x72814);
  nand n72818(x72818, x71637, x9719);
  nand n72819(x72819, x71135, x87021);
  nand n72820(x72820, x68462, x72822);
  nand n72821(x72821, x72820, x72819);
  nand n72823(x72823, x71637, x9740);
  nand n72824(x72824, x71135, x87022);
  nand n72825(x72825, x68462, x72827);
  nand n72826(x72826, x72825, x72824);
  nand n72828(x72828, x71637, x9761);
  nand n72829(x72829, x71135, x87023);
  nand n72830(x72830, x68462, x72832);
  nand n72831(x72831, x72830, x72829);
  nand n72833(x72833, x71637, x9782);
  nand n72834(x72834, x71135, x87024);
  nand n72835(x72835, x68462, x72837);
  nand n72836(x72836, x72835, x72834);
  nand n72838(x72838, x71637, x9803);
  nand n72839(x72839, x71135, x87025);
  nand n72840(x72840, x68462, x72842);
  nand n72841(x72841, x72840, x72839);
  nand n72843(x72843, x71637, x9824);
  nand n72844(x72844, x71135, x87026);
  nand n72845(x72845, x68462, x72847);
  nand n72846(x72846, x72845, x72844);
  nand n72848(x72848, x71637, x9845);
  nand n72849(x72849, x71135, x87027);
  nand n72850(x72850, x68462, x72852);
  nand n72851(x72851, x72850, x72849);
  nand n72853(x72853, x71637, x9866);
  nand n72854(x72854, x71135, x87028);
  nand n72855(x72855, x68462, x72857);
  nand n72856(x72856, x72855, x72854);
  nand n72858(x72858, x71637, x9887);
  nand n72859(x72859, x71135, x87029);
  nand n72860(x72860, x68462, x72862);
  nand n72861(x72861, x72860, x72859);
  nand n72863(x72863, x71637, x9908);
  nand n72864(x72864, x71135, x87030);
  nand n72865(x72865, x68462, x72867);
  nand n72866(x72866, x72865, x72864);
  nand n72868(x72868, x71637, x9929);
  nand n72869(x72869, x71135, x87031);
  nand n72870(x72870, x68462, x72872);
  nand n72871(x72871, x72870, x72869);
  nand n72873(x72873, x71637, x9950);
  nand n72874(x72874, x71135, x87032);
  nand n72875(x72875, x68462, x72877);
  nand n72876(x72876, x72875, x72874);
  nand n72878(x72878, x71637, x9971);
  nand n72879(x72879, x71135, x87033);
  nand n72880(x72880, x68462, x72882);
  nand n72881(x72881, x72880, x72879);
  nand n72883(x72883, x71637, x9992);
  nand n72884(x72884, x71135, x87034);
  nand n72885(x72885, x68462, x72887);
  nand n72886(x72886, x72885, x72884);
  nand n72888(x72888, x71637, x10013);
  nand n72889(x72889, x71135, x87035);
  nand n72890(x72890, x68462, x72892);
  nand n72891(x72891, x72890, x72889);
  nand n72893(x72893, x71637, x10034);
  nand n72894(x72894, x71135, x87036);
  nand n72895(x72895, x68462, x72897);
  nand n72896(x72896, x72895, x72894);
  nand n72898(x72898, x71637, x10055);
  nand n72899(x72899, x71135, x87037);
  nand n72900(x72900, x68462, x72902);
  nand n72901(x72901, x72900, x72899);
  nand n72903(x72903, x71637, x10076);
  nand n72904(x72904, x71135, x87038);
  nand n72905(x72905, x68462, x72907);
  nand n72906(x72906, x72905, x72904);
  nand n72908(x72908, x71637, x10097);
  nand n72909(x72909, x71135, x87039);
  nand n72910(x72910, x68462, x72912);
  nand n72911(x72911, x72910, x72909);
  nand n72913(x72913, x71637, x10118);
  nand n72914(x72914, x71135, x87040);
  nand n72915(x72915, x68462, x72917);
  nand n72916(x72916, x72915, x72914);
  nand n72918(x72918, x71637, x10139);
  nand n72919(x72919, x71135, x87041);
  nand n72920(x72920, x68462, x72922);
  nand n72921(x72921, x72920, x72919);
  nand n72923(x72923, x71637, x10160);
  nand n72924(x72924, x71135, x87042);
  nand n72925(x72925, x68462, x72927);
  nand n72926(x72926, x72925, x72924);
  nand n72928(x72928, x71637, x10181);
  nand n72929(x72929, x71135, x87043);
  nand n72930(x72930, x68462, x72932);
  nand n72931(x72931, x72930, x72929);
  nand n72933(x72933, x71637, x10202);
  nand n72934(x72934, x71135, x87044);
  nand n72935(x72935, x68462, x72937);
  nand n72936(x72936, x72935, x72934);
  nand n72938(x72938, x71637, x10223);
  nand n72939(x72939, x71135, x87045);
  nand n72940(x72940, x68462, x72942);
  nand n72941(x72941, x72940, x72939);
  nand n72943(x72943, x71637, x10244);
  nand n72944(x72944, x71135, x87046);
  nand n72945(x72945, x68462, x72947);
  nand n72946(x72946, x72945, x72944);
  nand n72948(x72948, x71637, x10265);
  nand n72949(x72949, x71135, x87047);
  nand n72950(x72950, x68462, x72952);
  nand n72951(x72951, x72950, x72949);
  nand n72953(x72953, x71637, x10286);
  nand n72954(x72954, x71135, x87048);
  nand n72955(x72955, x68462, x72957);
  nand n72956(x72956, x72955, x72954);
  nand n72958(x72958, x71637, x10307);
  nand n72959(x72959, x71135, x87049);
  nand n72960(x72960, x68462, x72962);
  nand n72961(x72961, x72960, x72959);
  nand n72963(x72963, x71637, x10328);
  nand n72964(x72964, x71135, x87050);
  nand n72965(x72965, x68462, x72967);
  nand n72966(x72966, x72965, x72964);
  nand n72968(x72968, x71637, x10349);
  nand n72969(x72969, x71135, x87051);
  nand n72970(x72970, x68462, x72972);
  nand n72971(x72971, x72970, x72969);
  nand n72973(x72973, x71637, x10370);
  nand n72974(x72974, x71135, x87052);
  nand n72975(x72975, x68462, x72977);
  nand n72976(x72976, x72975, x72974);
  nand n72978(x72978, x71637, x10391);
  nand n72979(x72979, x71135, x87053);
  nand n72980(x72980, x68462, x72982);
  nand n72981(x72981, x72980, x72979);
  nand n72983(x72983, x71637, x10412);
  nand n72984(x72984, x71135, x87054);
  nand n72985(x72985, x68462, x72987);
  nand n72986(x72986, x72985, x72984);
  nand n72988(x72988, x71637, x10433);
  nand n72989(x72989, x71135, x87055);
  nand n72990(x72990, x68462, x72992);
  nand n72991(x72991, x72990, x72989);
  nand n72993(x72993, x71637, x10454);
  nand n72994(x72994, x71135, x87056);
  nand n72995(x72995, x68462, x72997);
  nand n72996(x72996, x72995, x72994);
  nand n72998(x72998, x71637, x10475);
  nand n72999(x72999, x71135, x87057);
  nand n73000(x73000, x68462, x73002);
  nand n73001(x73001, x73000, x72999);
  nand n73003(x73003, x71637, x10496);
  nand n73004(x73004, x71135, x87058);
  nand n73005(x73005, x68462, x73007);
  nand n73006(x73006, x73005, x73004);
  nand n73008(x73008, x71637, x10517);
  nand n73009(x73009, x71135, x87059);
  nand n73010(x73010, x68462, x73012);
  nand n73011(x73011, x73010, x73009);
  nand n73013(x73013, x71637, x1515);
  nand n73014(x73014, x71135, x87060);
  nand n73015(x73015, x68462, x73017);
  nand n73016(x73016, x73015, x73014);
  nand n73018(x73018, x71637, x1536);
  nand n73019(x73019, x71135, x87061);
  nand n73020(x73020, x68462, x73022);
  nand n73021(x73021, x73020, x73019);
  nand n73023(x73023, x71637, x10538);
  nand n73024(x73024, x71135, x87062);
  nand n73025(x73025, x68462, x73027);
  nand n73026(x73026, x73025, x73024);
  nand n73028(x73028, x71637, x10559);
  nand n73029(x73029, x71135, x87063);
  nand n73030(x73030, x68462, x73032);
  nand n73031(x73031, x73030, x73029);
  nand n73033(x73033, x71637, x10580);
  nand n73034(x73034, x71135, x87064);
  nand n73035(x73035, x68462, x73037);
  nand n73036(x73036, x73035, x73034);
  nand n73038(x73038, x71637, x10601);
  nand n73039(x73039, x71135, x87065);
  nand n73040(x73040, x68462, x73042);
  nand n73041(x73041, x73040, x73039);
  nand n73043(x73043, x71637, x10622);
  nand n73044(x73044, x71135, x87066);
  nand n73045(x73045, x68462, x73047);
  nand n73046(x73046, x73045, x73044);
  nand n73048(x73048, x71637, x10643);
  nand n73049(x73049, x71135, x87067);
  nand n73050(x73050, x68462, x73052);
  nand n73051(x73051, x73050, x73049);
  nand n73053(x73053, x71637, x10664);
  nand n73054(x73054, x71135, x87068);
  nand n73055(x73055, x68462, x73057);
  nand n73056(x73056, x73055, x73054);
  nand n73058(x73058, x71637, x10685);
  nand n73059(x73059, x71135, x87069);
  nand n73060(x73060, x68462, x73062);
  nand n73061(x73061, x73060, x73059);
  nand n73063(x73063, x71637, x10706);
  nand n73064(x73064, x71135, x87070);
  nand n73065(x73065, x68462, x73067);
  nand n73066(x73066, x73065, x73064);
  nand n73068(x73068, x71637, x10727);
  nand n73069(x73069, x71135, x87071);
  nand n73070(x73070, x68462, x73072);
  nand n73071(x73071, x73070, x73069);
  nand n73073(x73073, x71637, x10748);
  nand n73074(x73074, x71135, x87072);
  nand n73075(x73075, x68462, x73077);
  nand n73076(x73076, x73075, x73074);
  nand n73078(x73078, x71637, x10769);
  nand n73079(x73079, x71135, x87073);
  nand n73080(x73080, x68462, x73082);
  nand n73081(x73081, x73080, x73079);
  nand n73083(x73083, x71637, x10790);
  nand n73084(x73084, x71135, x87074);
  nand n73085(x73085, x68462, x73087);
  nand n73086(x73086, x73085, x73084);
  nand n73088(x73088, x71637, x10811);
  nand n73089(x73089, x71135, x87075);
  nand n73090(x73090, x68462, x73092);
  nand n73091(x73091, x73090, x73089);
  nand n73093(x73093, x71637, x10832);
  nand n73094(x73094, x71135, x87076);
  nand n73095(x73095, x68462, x73097);
  nand n73096(x73096, x73095, x73094);
  nand n73098(x73098, x71637, x10853);
  nand n73099(x73099, x71135, x87077);
  nand n73100(x73100, x68462, x73102);
  nand n73101(x73101, x73100, x73099);
  nand n73103(x73103, x71637, x10874);
  nand n73104(x73104, x71135, x87078);
  nand n73105(x73105, x68462, x73107);
  nand n73106(x73106, x73105, x73104);
  nand n73108(x73108, x71637, x10895);
  nand n73109(x73109, x71135, x87079);
  nand n73110(x73110, x68462, x73112);
  nand n73111(x73111, x73110, x73109);
  nand n73113(x73113, x71637, x10916);
  nand n73114(x73114, x71135, x87080);
  nand n73115(x73115, x68462, x73117);
  nand n73116(x73116, x73115, x73114);
  nand n73118(x73118, x71637, x10937);
  nand n73119(x73119, x71135, x87081);
  nand n73120(x73120, x68462, x73122);
  nand n73121(x73121, x73120, x73119);
  nand n73123(x73123, x71637, x10958);
  nand n73124(x73124, x71135, x87082);
  nand n73125(x73125, x68462, x73127);
  nand n73126(x73126, x73125, x73124);
  nand n73128(x73128, x71637, x10979);
  nand n73129(x73129, x71135, x87083);
  nand n73130(x73130, x68462, x73132);
  nand n73131(x73131, x73130, x73129);
  nand n73133(x73133, x71637, x11000);
  nand n73134(x73134, x71135, x87084);
  nand n73135(x73135, x68462, x73137);
  nand n73136(x73136, x73135, x73134);
  nand n73138(x73138, x71637, x11021);
  nand n73139(x73139, x71135, x87085);
  nand n73140(x73140, x68462, x73142);
  nand n73141(x73141, x73140, x73139);
  nand n73143(x73143, x71637, x11042);
  nand n73144(x73144, x71135, x87086);
  nand n73145(x73145, x68462, x73147);
  nand n73146(x73146, x73145, x73144);
  nand n73148(x73148, x71637, x11063);
  nand n73149(x73149, x71135, x87087);
  nand n73150(x73150, x68462, x73152);
  nand n73151(x73151, x73150, x73149);
  nand n73153(x73153, x71637, x11084);
  nand n73154(x73154, x71135, x87088);
  nand n73155(x73155, x68462, x73157);
  nand n73156(x73156, x73155, x73154);
  nand n73158(x73158, x71637, x11105);
  nand n73159(x73159, x71135, x87089);
  nand n73160(x73160, x68462, x73162);
  nand n73161(x73161, x73160, x73159);
  nand n73163(x73163, x71637, x11126);
  nand n73164(x73164, x71135, x87090);
  nand n73165(x73165, x68462, x73167);
  nand n73166(x73166, x73165, x73164);
  nand n73168(x73168, x71637, x11147);
  nand n73169(x73169, x71135, x87091);
  nand n73170(x73170, x68462, x73172);
  nand n73171(x73171, x73170, x73169);
  nand n73173(x73173, x71637, x11168);
  nand n73174(x73174, x71135, x87092);
  nand n73175(x73175, x68462, x73177);
  nand n73176(x73176, x73175, x73174);
  nand n73178(x73178, x71637, x11189);
  nand n73179(x73179, x71135, x87093);
  nand n73180(x73180, x68462, x73182);
  nand n73181(x73181, x73180, x73179);
  nand n73183(x73183, x71637, x11210);
  nand n73184(x73184, x71135, x87094);
  nand n73185(x73185, x68462, x73187);
  nand n73186(x73186, x73185, x73184);
  nand n73188(x73188, x71637, x11231);
  nand n73189(x73189, x71135, x87095);
  nand n73190(x73190, x68462, x73192);
  nand n73191(x73191, x73190, x73189);
  nand n73193(x73193, x71637, x11252);
  nand n73194(x73194, x71135, x87096);
  nand n73195(x73195, x68462, x73197);
  nand n73196(x73196, x73195, x73194);
  nand n73198(x73198, x71637, x11273);
  nand n73199(x73199, x71135, x87097);
  nand n73200(x73200, x68462, x73202);
  nand n73201(x73201, x73200, x73199);
  nand n73203(x73203, x71637, x11294);
  nand n73204(x73204, x71135, x87098);
  nand n73205(x73205, x68462, x73207);
  nand n73206(x73206, x73205, x73204);
  nand n73208(x73208, x71637, x11315);
  nand n73209(x73209, x71135, x87099);
  nand n73210(x73210, x68462, x73212);
  nand n73211(x73211, x73210, x73209);
  nand n73213(x73213, x71637, x11336);
  nand n73214(x73214, x71135, x87100);
  nand n73215(x73215, x68462, x73217);
  nand n73216(x73216, x73215, x73214);
  nand n73218(x73218, x71637, x11357);
  nand n73219(x73219, x71135, x87101);
  nand n73220(x73220, x68462, x73222);
  nand n73221(x73221, x73220, x73219);
  nand n73223(x73223, x71637, x11378);
  nand n73224(x73224, x71135, x87102);
  nand n73225(x73225, x68462, x73227);
  nand n73226(x73226, x73225, x73224);
  nand n73228(x73228, x71637, x11399);
  nand n73229(x73229, x71135, x87103);
  nand n73230(x73230, x68462, x73232);
  nand n73231(x73231, x73230, x73229);
  nand n73233(x73233, x71637, x11420);
  nand n73234(x73234, x71135, x87104);
  nand n73235(x73235, x68462, x73237);
  nand n73236(x73236, x73235, x73234);
  nand n73238(x73238, x71637, x11441);
  nand n73239(x73239, x71135, x87105);
  nand n73240(x73240, x68462, x73242);
  nand n73241(x73241, x73240, x73239);
  nand n73243(x73243, x71637, x11462);
  nand n73244(x73244, x71135, x87106);
  nand n73245(x73245, x68462, x73247);
  nand n73246(x73246, x73245, x73244);
  nand n73248(x73248, x71637, x11483);
  nand n73249(x73249, x71135, x87107);
  nand n73250(x73250, x68462, x73252);
  nand n73251(x73251, x73250, x73249);
  nand n73253(x73253, x71637, x11504);
  nand n73254(x73254, x71135, x87108);
  nand n73255(x73255, x68462, x73257);
  nand n73256(x73256, x73255, x73254);
  nand n73258(x73258, x71637, x11525);
  nand n73259(x73259, x71135, x87109);
  nand n73260(x73260, x68462, x73262);
  nand n73261(x73261, x73260, x73259);
  nand n73263(x73263, x71637, x11546);
  nand n73264(x73264, x71135, x87110);
  nand n73265(x73265, x68462, x73267);
  nand n73266(x73266, x73265, x73264);
  nand n73268(x73268, x71637, x11567);
  nand n73269(x73269, x71135, x87111);
  nand n73270(x73270, x68462, x73272);
  nand n73271(x73271, x73270, x73269);
  nand n73273(x73273, x71637, x11588);
  nand n73274(x73274, x71135, x87112);
  nand n73275(x73275, x68462, x73277);
  nand n73276(x73276, x73275, x73274);
  nand n73278(x73278, x71637, x11609);
  nand n73279(x73279, x71135, x87113);
  nand n73280(x73280, x68462, x73282);
  nand n73281(x73281, x73280, x73279);
  nand n73283(x73283, x71637, x11630);
  nand n73284(x73284, x71135, x87114);
  nand n73285(x73285, x68462, x73287);
  nand n73286(x73286, x73285, x73284);
  nand n73288(x73288, x71637, x11651);
  nand n73289(x73289, x71135, x87115);
  nand n73290(x73290, x68462, x73292);
  nand n73291(x73291, x73290, x73289);
  nand n73293(x73293, x71637, x11672);
  nand n73294(x73294, x71135, x87116);
  nand n73295(x73295, x68462, x73297);
  nand n73296(x73296, x73295, x73294);
  nand n73298(x73298, x71637, x11693);
  nand n73299(x73299, x71135, x87117);
  nand n73300(x73300, x68462, x73302);
  nand n73301(x73301, x73300, x73299);
  nand n73303(x73303, x71637, x11714);
  nand n73304(x73304, x71135, x87118);
  nand n73305(x73305, x68462, x73307);
  nand n73306(x73306, x73305, x73304);
  nand n73308(x73308, x71637, x11735);
  nand n73309(x73309, x71135, x87119);
  nand n73310(x73310, x68462, x73312);
  nand n73311(x73311, x73310, x73309);
  nand n73313(x73313, x71637, x11756);
  nand n73314(x73314, x71135, x87120);
  nand n73315(x73315, x68462, x73317);
  nand n73316(x73316, x73315, x73314);
  nand n73318(x73318, x71637, x11777);
  nand n73319(x73319, x71135, x87121);
  nand n73320(x73320, x68462, x73322);
  nand n73321(x73321, x73320, x73319);
  nand n73323(x73323, x71637, x11798);
  nand n73324(x73324, x71135, x87122);
  nand n73325(x73325, x68462, x73327);
  nand n73326(x73326, x73325, x73324);
  nand n73328(x73328, x71637, x11819);
  nand n73329(x73329, x71135, x87123);
  nand n73330(x73330, x68462, x73332);
  nand n73331(x73331, x73330, x73329);
  nand n73333(x73333, x71637, x11840);
  nand n73334(x73334, x71135, x87124);
  nand n73335(x73335, x68462, x73337);
  nand n73336(x73336, x73335, x73334);
  nand n73338(x73338, x71637, x11861);
  nand n73339(x73339, x71135, x87125);
  nand n73340(x73340, x68462, x73342);
  nand n73341(x73341, x73340, x73339);
  nand n73343(x73343, x71637, x11882);
  nand n73344(x73344, x71135, x87126);
  nand n73345(x73345, x68462, x73347);
  nand n73346(x73346, x73345, x73344);
  nand n73348(x73348, x71637, x11903);
  nand n73349(x73349, x71135, x87127);
  nand n73350(x73350, x68462, x73352);
  nand n73351(x73351, x73350, x73349);
  nand n73353(x73353, x71637, x11924);
  nand n73354(x73354, x71135, x87128);
  nand n73355(x73355, x68462, x73357);
  nand n73356(x73356, x73355, x73354);
  nand n73358(x73358, x71637, x11945);
  nand n73359(x73359, x71135, x87129);
  nand n73360(x73360, x68462, x73362);
  nand n73361(x73361, x73360, x73359);
  nand n73363(x73363, x71637, x11966);
  nand n73364(x73364, x71135, x87130);
  nand n73365(x73365, x68462, x73367);
  nand n73366(x73366, x73365, x73364);
  nand n73368(x73368, x71637, x11987);
  nand n73369(x73369, x71135, x87131);
  nand n73370(x73370, x68462, x73372);
  nand n73371(x73371, x73370, x73369);
  nand n73373(x73373, x71637, x12008);
  nand n73374(x73374, x71135, x87132);
  nand n73375(x73375, x68462, x73377);
  nand n73376(x73376, x73375, x73374);
  nand n73378(x73378, x71637, x12029);
  nand n73379(x73379, x71135, x87133);
  nand n73380(x73380, x68462, x73382);
  nand n73381(x73381, x73380, x73379);
  nand n73383(x73383, x71637, x12050);
  nand n73384(x73384, x71135, x87134);
  nand n73385(x73385, x68462, x73387);
  nand n73386(x73386, x73385, x73384);
  nand n73388(x73388, x71637, x12071);
  nand n73389(x73389, x71135, x87135);
  nand n73390(x73390, x68462, x73392);
  nand n73391(x73391, x73390, x73389);
  nand n73393(x73393, x71637, x12092);
  nand n73394(x73394, x71135, x87136);
  nand n73395(x73395, x68462, x73397);
  nand n73396(x73396, x73395, x73394);
  nand n73398(x73398, x71637, x12113);
  nand n73399(x73399, x71135, x87137);
  nand n73400(x73400, x68462, x73402);
  nand n73401(x73401, x73400, x73399);
  nand n73403(x73403, x71637, x12134);
  nand n73404(x73404, x71135, x87138);
  nand n73405(x73405, x68462, x73407);
  nand n73406(x73406, x73405, x73404);
  nand n73408(x73408, x71637, x12155);
  nand n73409(x73409, x71135, x87139);
  nand n73410(x73410, x68462, x73412);
  nand n73411(x73411, x73410, x73409);
  nand n73413(x73413, x71637, x12176);
  nand n73414(x73414, x71135, x87140);
  nand n73415(x73415, x68462, x73417);
  nand n73416(x73416, x73415, x73414);
  nand n73418(x73418, x71637, x12197);
  nand n73419(x73419, x71135, x87141);
  nand n73420(x73420, x68462, x73422);
  nand n73421(x73421, x73420, x73419);
  nand n73423(x73423, x71637, x12218);
  nand n73424(x73424, x71135, x87142);
  nand n73425(x73425, x68462, x73427);
  nand n73426(x73426, x73425, x73424);
  nand n73428(x73428, x71637, x12239);
  nand n73429(x73429, x71135, x87143);
  nand n73430(x73430, x68462, x73432);
  nand n73431(x73431, x73430, x73429);
  nand n73433(x73433, x71637, x12260);
  nand n73434(x73434, x71135, x87144);
  nand n73435(x73435, x68462, x73437);
  nand n73436(x73436, x73435, x73434);
  nand n73438(x73438, x71637, x12281);
  nand n73439(x73439, x71135, x87145);
  nand n73440(x73440, x68462, x73442);
  nand n73441(x73441, x73440, x73439);
  nand n73443(x73443, x71637, x12302);
  nand n73444(x73444, x71135, x87146);
  nand n73445(x73445, x68462, x73447);
  nand n73446(x73446, x73445, x73444);
  nand n73448(x73448, x71637, x12323);
  nand n73449(x73449, x71135, x87147);
  nand n73450(x73450, x68462, x73452);
  nand n73451(x73451, x73450, x73449);
  nand n73453(x73453, x71637, x12344);
  nand n73454(x73454, x71135, x87148);
  nand n73455(x73455, x68462, x73457);
  nand n73456(x73456, x73455, x73454);
  nand n73458(x73458, x71637, x12365);
  nand n73459(x73459, x71135, x87149);
  nand n73460(x73460, x68462, x73462);
  nand n73461(x73461, x73460, x73459);
  nand n73463(x73463, x71637, x12386);
  nand n73464(x73464, x71135, x87150);
  nand n73465(x73465, x68462, x73467);
  nand n73466(x73466, x73465, x73464);
  nand n73468(x73468, x71637, x12407);
  nand n73469(x73469, x71135, x87151);
  nand n73470(x73470, x68462, x73472);
  nand n73471(x73471, x73470, x73469);
  nand n73473(x73473, x71637, x12428);
  nand n73474(x73474, x71135, x87152);
  nand n73475(x73475, x68462, x73477);
  nand n73476(x73476, x73475, x73474);
  nand n73478(x73478, x71637, x12449);
  nand n73479(x73479, x71135, x87153);
  nand n73480(x73480, x68462, x73482);
  nand n73481(x73481, x73480, x73479);
  nand n73483(x73483, x71637, x12470);
  nand n73484(x73484, x71135, x87154);
  nand n73485(x73485, x68462, x73487);
  nand n73486(x73486, x73485, x73484);
  nand n73488(x73488, x71637, x12491);
  nand n73489(x73489, x71135, x87155);
  nand n73490(x73490, x68462, x73492);
  nand n73491(x73491, x73490, x73489);
  nand n73493(x73493, x71637, x12512);
  nand n73494(x73494, x71135, x87156);
  nand n73495(x73495, x68462, x73497);
  nand n73496(x73496, x73495, x73494);
  nand n73498(x73498, x71637, x12533);
  nand n73499(x73499, x71135, x87157);
  nand n73500(x73500, x68462, x73502);
  nand n73501(x73501, x73500, x73499);
  nand n73503(x73503, x71637, x1578);
  nand n73504(x73504, x71135, x87158);
  nand n73505(x73505, x68462, x73507);
  nand n73506(x73506, x73505, x73504);
  nand n73508(x73508, x71637, x1599);
  nand n73509(x73509, x71135, x87159);
  nand n73510(x73510, x68462, x73512);
  nand n73511(x73511, x73510, x73509);
  nand n73513(x73513, x71637, x12554);
  nand n73514(x73514, x71135, x87160);
  nand n73515(x73515, x68462, x73517);
  nand n73516(x73516, x73515, x73514);
  nand n73518(x73518, x71637, x12575);
  nand n73519(x73519, x71135, x87161);
  nand n73520(x73520, x68462, x73522);
  nand n73521(x73521, x73520, x73519);
  nand n73523(x73523, x71637, x12596);
  nand n73524(x73524, x71135, x87162);
  nand n73525(x73525, x68462, x73527);
  nand n73526(x73526, x73525, x73524);
  nand n73528(x73528, x71637, x12617);
  nand n73529(x73529, x71135, x87163);
  nand n73530(x73530, x68462, x73532);
  nand n73531(x73531, x73530, x73529);
  nand n73533(x73533, x71637, x12638);
  nand n73534(x73534, x71135, x87164);
  nand n73535(x73535, x68462, x73537);
  nand n73536(x73536, x73535, x73534);
  nand n73538(x73538, x71637, x12659);
  nand n73539(x73539, x71135, x87165);
  nand n73540(x73540, x68462, x73542);
  nand n73541(x73541, x73540, x73539);
  nand n73543(x73543, x71637, x12680);
  nand n73544(x73544, x71135, x87166);
  nand n73545(x73545, x68462, x73547);
  nand n73546(x73546, x73545, x73544);
  nand n73548(x73548, x71637, x12701);
  nand n73549(x73549, x71135, x87167);
  nand n73550(x73550, x68462, x73552);
  nand n73551(x73551, x73550, x73549);
  nand n73553(x73553, x71637, x12722);
  nand n73554(x73554, x71135, x87168);
  nand n73555(x73555, x68462, x73557);
  nand n73556(x73556, x73555, x73554);
  nand n73558(x73558, x71637, x12743);
  nand n73559(x73559, x71135, x87169);
  nand n73560(x73560, x68462, x73562);
  nand n73561(x73561, x73560, x73559);
  nand n73563(x73563, x71637, x12764);
  nand n73564(x73564, x71135, x87170);
  nand n73565(x73565, x68462, x73567);
  nand n73566(x73566, x73565, x73564);
  nand n73568(x73568, x71637, x12785);
  nand n73569(x73569, x71135, x87171);
  nand n73570(x73570, x68462, x73572);
  nand n73571(x73571, x73570, x73569);
  nand n73573(x73573, x71637, x12806);
  nand n73574(x73574, x71135, x87172);
  nand n73575(x73575, x68462, x73577);
  nand n73576(x73576, x73575, x73574);
  nand n73578(x73578, x71637, x12827);
  nand n73579(x73579, x71135, x87173);
  nand n73580(x73580, x68462, x73582);
  nand n73581(x73581, x73580, x73579);
  nand n73583(x73583, x71637, x12848);
  nand n73584(x73584, x71135, x87174);
  nand n73585(x73585, x68462, x73587);
  nand n73586(x73586, x73585, x73584);
  nand n73588(x73588, x71637, x12869);
  nand n73589(x73589, x71135, x87175);
  nand n73590(x73590, x68462, x73592);
  nand n73591(x73591, x73590, x73589);
  nand n73593(x73593, x71637, x12890);
  nand n73594(x73594, x71135, x87176);
  nand n73595(x73595, x68462, x73597);
  nand n73596(x73596, x73595, x73594);
  nand n73598(x73598, x71637, x12911);
  nand n73599(x73599, x71135, x87177);
  nand n73600(x73600, x68462, x73602);
  nand n73601(x73601, x73600, x73599);
  nand n73603(x73603, x71637, x12932);
  nand n73604(x73604, x71135, x87178);
  nand n73605(x73605, x68462, x73607);
  nand n73606(x73606, x73605, x73604);
  nand n73608(x73608, x71637, x12953);
  nand n73609(x73609, x71135, x87179);
  nand n73610(x73610, x68462, x73612);
  nand n73611(x73611, x73610, x73609);
  nand n73613(x73613, x71637, x12974);
  nand n73614(x73614, x71135, x87180);
  nand n73615(x73615, x68462, x73617);
  nand n73616(x73616, x73615, x73614);
  nand n73618(x73618, x71637, x12995);
  nand n73619(x73619, x71135, x87181);
  nand n73620(x73620, x68462, x73622);
  nand n73621(x73621, x73620, x73619);
  nand n73623(x73623, x71637, x13016);
  nand n73624(x73624, x71135, x87182);
  nand n73625(x73625, x68462, x73627);
  nand n73626(x73626, x73625, x73624);
  nand n73628(x73628, x71637, x13037);
  nand n73629(x73629, x71135, x87183);
  nand n73630(x73630, x68462, x73632);
  nand n73631(x73631, x73630, x73629);
  nand n73633(x73633, x71637, x13058);
  nand n73634(x73634, x71135, x87184);
  nand n73635(x73635, x68462, x73637);
  nand n73636(x73636, x73635, x73634);
  nand n73638(x73638, x71637, x13079);
  nand n73639(x73639, x71135, x87185);
  nand n73640(x73640, x68462, x73642);
  nand n73641(x73641, x73640, x73639);
  nand n73643(x73643, x71637, x13100);
  nand n73644(x73644, x71135, x87186);
  nand n73645(x73645, x68462, x73647);
  nand n73646(x73646, x73645, x73644);
  nand n73648(x73648, x71637, x13121);
  nand n73649(x73649, x71135, x87187);
  nand n73650(x73650, x68462, x73652);
  nand n73651(x73651, x73650, x73649);
  nand n73653(x73653, x71637, x13142);
  nand n73654(x73654, x71135, x87188);
  nand n73655(x73655, x68462, x73657);
  nand n73656(x73656, x73655, x73654);
  nand n73658(x73658, x71637, x13163);
  nand n73659(x73659, x71135, x87189);
  nand n73660(x73660, x68462, x73662);
  nand n73661(x73661, x73660, x73659);
  nand n73663(x73663, x71637, x13184);
  nand n73664(x73664, x71135, x87190);
  nand n73665(x73665, x68462, x73667);
  nand n73666(x73666, x73665, x73664);
  nand n73668(x73668, x71637, x13205);
  nand n73669(x73669, x71135, x87191);
  nand n73670(x73670, x68462, x73672);
  nand n73671(x73671, x73670, x73669);
  nand n73673(x73673, x71637, x13226);
  nand n73674(x73674, x71135, x87192);
  nand n73675(x73675, x68462, x73677);
  nand n73676(x73676, x73675, x73674);
  nand n73678(x73678, x71637, x13247);
  nand n73679(x73679, x71135, x87193);
  nand n73680(x73680, x68462, x73682);
  nand n73681(x73681, x73680, x73679);
  nand n73683(x73683, x71637, x13268);
  nand n73684(x73684, x71135, x87194);
  nand n73685(x73685, x68462, x73687);
  nand n73686(x73686, x73685, x73684);
  nand n73688(x73688, x71637, x13289);
  nand n73689(x73689, x71135, x87195);
  nand n73690(x73690, x68462, x73692);
  nand n73691(x73691, x73690, x73689);
  nand n73693(x73693, x71637, x13310);
  nand n73694(x73694, x71135, x87196);
  nand n73695(x73695, x68462, x73697);
  nand n73696(x73696, x73695, x73694);
  nand n73698(x73698, x71637, x13331);
  nand n73699(x73699, x71135, x87197);
  nand n73700(x73700, x68462, x73702);
  nand n73701(x73701, x73700, x73699);
  nand n73703(x73703, x71637, x13352);
  nand n73704(x73704, x71135, x87198);
  nand n73705(x73705, x68462, x73707);
  nand n73706(x73706, x73705, x73704);
  nand n73708(x73708, x71637, x13373);
  nand n73709(x73709, x71135, x87199);
  nand n73710(x73710, x68462, x73712);
  nand n73711(x73711, x73710, x73709);
  nand n73713(x73713, x71637, x13394);
  nand n73714(x73714, x71135, x87200);
  nand n73715(x73715, x68462, x73717);
  nand n73716(x73716, x73715, x73714);
  nand n73718(x73718, x71637, x13415);
  nand n73719(x73719, x71135, x87201);
  nand n73720(x73720, x68462, x73722);
  nand n73721(x73721, x73720, x73719);
  nand n73723(x73723, x71637, x13436);
  nand n73724(x73724, x71135, x87202);
  nand n73725(x73725, x68462, x73727);
  nand n73726(x73726, x73725, x73724);
  nand n73728(x73728, x71637, x13457);
  nand n73729(x73729, x71135, x87203);
  nand n73730(x73730, x68462, x73732);
  nand n73731(x73731, x73730, x73729);
  nand n73733(x73733, x71637, x13478);
  nand n73734(x73734, x71135, x87204);
  nand n73735(x73735, x68462, x73737);
  nand n73736(x73736, x73735, x73734);
  nand n73738(x73738, x71637, x13499);
  nand n73739(x73739, x71135, x87205);
  nand n73740(x73740, x68462, x73742);
  nand n73741(x73741, x73740, x73739);
  nand n73743(x73743, x71637, x13520);
  nand n73744(x73744, x71135, x87206);
  nand n73745(x73745, x68462, x73747);
  nand n73746(x73746, x73745, x73744);
  nand n73748(x73748, x71637, x13541);
  nand n73749(x73749, x71135, x87207);
  nand n73750(x73750, x68462, x73752);
  nand n73751(x73751, x73750, x73749);
  nand n73753(x73753, x71637, x13562);
  nand n73754(x73754, x71135, x87208);
  nand n73755(x73755, x68462, x73757);
  nand n73756(x73756, x73755, x73754);
  nand n73758(x73758, x71637, x13583);
  nand n73759(x73759, x71135, x87209);
  nand n73760(x73760, x68462, x73762);
  nand n73761(x73761, x73760, x73759);
  nand n73763(x73763, x71637, x13604);
  nand n73764(x73764, x71135, x87210);
  nand n73765(x73765, x68462, x73767);
  nand n73766(x73766, x73765, x73764);
  nand n73768(x73768, x71637, x13625);
  nand n73769(x73769, x71135, x87211);
  nand n73770(x73770, x68462, x73772);
  nand n73771(x73771, x73770, x73769);
  nand n73773(x73773, x71637, x13646);
  nand n73774(x73774, x71135, x87212);
  nand n73775(x73775, x68462, x73777);
  nand n73776(x73776, x73775, x73774);
  nand n73778(x73778, x71637, x13667);
  nand n73779(x73779, x71135, x87213);
  nand n73780(x73780, x68462, x73782);
  nand n73781(x73781, x73780, x73779);
  nand n73783(x73783, x71637, x13688);
  nand n73784(x73784, x71135, x87214);
  nand n73785(x73785, x68462, x73787);
  nand n73786(x73786, x73785, x73784);
  nand n73788(x73788, x71637, x13709);
  nand n73789(x73789, x71135, x87215);
  nand n73790(x73790, x68462, x73792);
  nand n73791(x73791, x73790, x73789);
  nand n73793(x73793, x71637, x13730);
  nand n73794(x73794, x71135, x87216);
  nand n73795(x73795, x68462, x73797);
  nand n73796(x73796, x73795, x73794);
  nand n73798(x73798, x71637, x13751);
  nand n73799(x73799, x71135, x87217);
  nand n73800(x73800, x68462, x73802);
  nand n73801(x73801, x73800, x73799);
  nand n73803(x73803, x71637, x13772);
  nand n73804(x73804, x71135, x87218);
  nand n73805(x73805, x68462, x73807);
  nand n73806(x73806, x73805, x73804);
  nand n73808(x73808, x71637, x13793);
  nand n73809(x73809, x71135, x87219);
  nand n73810(x73810, x68462, x73812);
  nand n73811(x73811, x73810, x73809);
  nand n73813(x73813, x71637, x13814);
  nand n73814(x73814, x71135, x87220);
  nand n73815(x73815, x68462, x73817);
  nand n73816(x73816, x73815, x73814);
  nand n73818(x73818, x71637, x13835);
  nand n73819(x73819, x71135, x87221);
  nand n73820(x73820, x68462, x73822);
  nand n73821(x73821, x73820, x73819);
  nand n73823(x73823, x71637, x13856);
  nand n73824(x73824, x71135, x87222);
  nand n73825(x73825, x68462, x73827);
  nand n73826(x73826, x73825, x73824);
  nand n73828(x73828, x71637, x13877);
  nand n73829(x73829, x71135, x87223);
  nand n73830(x73830, x68462, x73832);
  nand n73831(x73831, x73830, x73829);
  nand n73833(x73833, x71637, x13898);
  nand n73834(x73834, x71135, x87224);
  nand n73835(x73835, x68462, x73837);
  nand n73836(x73836, x73835, x73834);
  nand n73838(x73838, x71637, x13919);
  nand n73839(x73839, x71135, x87225);
  nand n73840(x73840, x68462, x73842);
  nand n73841(x73841, x73840, x73839);
  nand n73843(x73843, x71637, x13940);
  nand n73844(x73844, x71135, x87226);
  nand n73845(x73845, x68462, x73847);
  nand n73846(x73846, x73845, x73844);
  nand n73848(x73848, x71637, x13961);
  nand n73849(x73849, x71135, x87227);
  nand n73850(x73850, x68462, x73852);
  nand n73851(x73851, x73850, x73849);
  nand n73853(x73853, x71637, x13982);
  nand n73854(x73854, x71135, x87228);
  nand n73855(x73855, x68462, x73857);
  nand n73856(x73856, x73855, x73854);
  nand n73858(x73858, x71637, x14003);
  nand n73859(x73859, x71135, x87229);
  nand n73860(x73860, x68462, x73862);
  nand n73861(x73861, x73860, x73859);
  nand n73863(x73863, x71637, x14024);
  nand n73864(x73864, x71135, x87230);
  nand n73865(x73865, x68462, x73867);
  nand n73866(x73866, x73865, x73864);
  nand n73868(x73868, x71637, x14045);
  nand n73869(x73869, x71135, x87231);
  nand n73870(x73870, x68462, x73872);
  nand n73871(x73871, x73870, x73869);
  nand n73873(x73873, x71637, x14066);
  nand n73874(x73874, x71135, x87232);
  nand n73875(x73875, x68462, x73877);
  nand n73876(x73876, x73875, x73874);
  nand n73878(x73878, x71637, x14087);
  nand n73879(x73879, x71135, x87233);
  nand n73880(x73880, x68462, x73882);
  nand n73881(x73881, x73880, x73879);
  nand n73883(x73883, x71637, x14108);
  nand n73884(x73884, x71135, x87234);
  nand n73885(x73885, x68462, x73887);
  nand n73886(x73886, x73885, x73884);
  nand n73888(x73888, x71637, x14129);
  nand n73889(x73889, x71135, x87235);
  nand n73890(x73890, x68462, x73892);
  nand n73891(x73891, x73890, x73889);
  nand n73893(x73893, x71637, x14150);
  nand n73894(x73894, x71135, x87236);
  nand n73895(x73895, x68462, x73897);
  nand n73896(x73896, x73895, x73894);
  nand n73898(x73898, x71637, x14171);
  nand n73899(x73899, x71135, x87237);
  nand n73900(x73900, x68462, x73902);
  nand n73901(x73901, x73900, x73899);
  nand n73903(x73903, x71637, x14192);
  nand n73904(x73904, x71135, x87238);
  nand n73905(x73905, x68462, x73907);
  nand n73906(x73906, x73905, x73904);
  nand n73908(x73908, x71637, x14213);
  nand n73909(x73909, x71135, x87239);
  nand n73910(x73910, x68462, x73912);
  nand n73911(x73911, x73910, x73909);
  nand n73913(x73913, x71637, x14234);
  nand n73914(x73914, x71135, x87240);
  nand n73915(x73915, x68462, x73917);
  nand n73916(x73916, x73915, x73914);
  nand n73918(x73918, x71637, x14255);
  nand n73919(x73919, x71135, x87241);
  nand n73920(x73920, x68462, x73922);
  nand n73921(x73921, x73920, x73919);
  nand n73923(x73923, x71637, x14276);
  nand n73924(x73924, x71135, x87242);
  nand n73925(x73925, x68462, x73927);
  nand n73926(x73926, x73925, x73924);
  nand n73928(x73928, x71637, x14297);
  nand n73929(x73929, x71135, x87243);
  nand n73930(x73930, x68462, x73932);
  nand n73931(x73931, x73930, x73929);
  nand n73933(x73933, x71637, x14318);
  nand n73934(x73934, x71135, x87244);
  nand n73935(x73935, x68462, x73937);
  nand n73936(x73936, x73935, x73934);
  nand n73938(x73938, x71637, x14339);
  nand n73939(x73939, x71135, x87245);
  nand n73940(x73940, x68462, x73942);
  nand n73941(x73941, x73940, x73939);
  nand n73943(x73943, x71637, x14360);
  nand n73944(x73944, x71135, x87246);
  nand n73945(x73945, x68462, x73947);
  nand n73946(x73946, x73945, x73944);
  nand n73948(x73948, x71637, x14381);
  nand n73949(x73949, x71135, x87247);
  nand n73950(x73950, x68462, x73952);
  nand n73951(x73951, x73950, x73949);
  nand n73953(x73953, x71637, x14402);
  nand n73954(x73954, x71135, x87248);
  nand n73955(x73955, x68462, x73957);
  nand n73956(x73956, x73955, x73954);
  nand n73958(x73958, x71637, x14423);
  nand n73959(x73959, x71135, x87249);
  nand n73960(x73960, x68462, x73962);
  nand n73961(x73961, x73960, x73959);
  nand n73963(x73963, x71637, x14444);
  nand n73964(x73964, x71135, x87250);
  nand n73965(x73965, x68462, x73967);
  nand n73966(x73966, x73965, x73964);
  nand n73968(x73968, x71637, x14465);
  nand n73969(x73969, x71135, x87251);
  nand n73970(x73970, x68462, x73972);
  nand n73971(x73971, x73970, x73969);
  nand n73973(x73973, x71637, x14486);
  nand n73974(x73974, x71135, x87252);
  nand n73975(x73975, x68462, x73977);
  nand n73976(x73976, x73975, x73974);
  nand n73978(x73978, x71637, x14507);
  nand n73979(x73979, x71135, x87253);
  nand n73980(x73980, x68462, x73982);
  nand n73981(x73981, x73980, x73979);
  nand n73983(x73983, x71637, x14528);
  nand n73984(x73984, x71135, x87254);
  nand n73985(x73985, x68462, x73987);
  nand n73986(x73986, x73985, x73984);
  nand n73988(x73988, x71637, x14549);
  nand n73989(x73989, x71135, x87255);
  nand n73990(x73990, x68462, x73992);
  nand n73991(x73991, x73990, x73989);
  nand n73993(x73993, x71637, x1641);
  nand n73994(x73994, x71135, x87256);
  nand n73995(x73995, x68462, x73997);
  nand n73996(x73996, x73995, x73994);
  nand n73998(x73998, x71637, x1662);
  nand n73999(x73999, x71135, x87257);
  nand n74000(x74000, x68462, x74002);
  nand n74001(x74001, x74000, x73999);
  nand n74003(x74003, x68462, x74005);
  nand n74004(x74004, x74003, x71799);
  nand n74006(x74006, x68462, x74008);
  nand n74007(x74007, x74006, x71804);
  nand n74009(x74009, x68462, x74011);
  nand n74010(x74010, x74009, x71809);
  nand n74012(x74012, x68462, x74014);
  nand n74013(x74013, x74012, x71814);
  nand n74015(x74015, x68462, x74017);
  nand n74016(x74016, x74015, x71819);
  nand n74018(x74018, x68462, x74020);
  nand n74019(x74019, x74018, x71824);
  nand n74021(x74021, x68462, x74023);
  nand n74022(x74022, x74021, x71829);
  nand n74024(x74024, x68462, x74026);
  nand n74025(x74025, x74024, x71834);
  nand n74027(x74027, x68462, x74029);
  nand n74028(x74028, x74027, x71839);
  nand n74030(x74030, x68462, x74032);
  nand n74031(x74031, x74030, x71844);
  nand n74033(x74033, x68462, x74035);
  nand n74034(x74034, x74033, x71849);
  nand n74036(x74036, x68462, x74038);
  nand n74037(x74037, x74036, x71854);
  nand n74039(x74039, x68462, x74041);
  nand n74040(x74040, x74039, x71859);
  nand n74042(x74042, x68462, x74044);
  nand n74043(x74043, x74042, x71864);
  nand n74045(x74045, x68462, x74047);
  nand n74046(x74046, x74045, x71869);
  nand n74048(x74048, x68462, x74050);
  nand n74049(x74049, x74048, x71874);
  nand n74051(x74051, x68462, x74053);
  nand n74052(x74052, x74051, x71879);
  nand n74054(x74054, x68462, x74056);
  nand n74055(x74055, x74054, x71884);
  nand n74057(x74057, x68462, x74059);
  nand n74058(x74058, x74057, x71889);
  nand n74060(x74060, x68462, x74062);
  nand n74061(x74061, x74060, x71894);
  nand n74063(x74063, x68462, x74065);
  nand n74064(x74064, x74063, x71899);
  nand n74066(x74066, x68462, x74068);
  nand n74067(x74067, x74066, x71904);
  nand n74069(x74069, x68462, x74071);
  nand n74070(x74070, x74069, x71904);
  nand n74072(x74072, x68462, x74074);
  nand n74073(x74073, x74072, x71904);
  nand n74075(x74075, x68462, x74077);
  nand n74076(x74076, x74075, x71904);
  nand n74078(x74078, x68462, x74080);
  nand n74079(x74079, x74078, x71904);
  nand n74081(x74081, x68462, x74083);
  nand n74082(x74082, x74081, x71904);
  nand n74084(x74084, x68462, x74086);
  nand n74085(x74085, x74084, x71904);
  nand n74087(x74087, x68462, x74089);
  nand n74088(x74088, x74087, x71904);
  nand n74090(x74090, x68462, x74092);
  nand n74091(x74091, x74090, x71904);
  nand n74093(x74093, x68462, x74095);
  nand n74094(x74094, x74093, x71904);
  nand n74096(x74096, x68462, x74098);
  nand n74097(x74097, x74096, x71904);
  nand n74099(x74099, x68462, x74101);
  nand n74100(x74100, x74099, x71939);
  nand n74102(x74102, x68462, x74104);
  nand n74103(x74103, x74102, x71944);
  nand n74105(x74105, x68462, x74107);
  nand n74106(x74106, x74105, x71949);
  nand n74108(x74108, x68462, x74110);
  nand n74109(x74109, x74108, x71954);
  nand n74111(x74111, x68462, x74113);
  nand n74112(x74112, x74111, x71959);
  nand n74114(x74114, x68462, x74116);
  nand n74115(x74115, x74114, x71964);
  nand n74117(x74117, x68462, x74119);
  nand n74118(x74118, x74117, x71969);
  nand n74120(x74120, x68462, x74122);
  nand n74121(x74121, x74120, x71974);
  nand n74123(x74123, x68462, x74125);
  nand n74124(x74124, x74123, x71979);
  nand n74126(x74126, x68462, x74128);
  nand n74127(x74127, x74126, x71984);
  nand n74129(x74129, x68462, x74131);
  nand n74130(x74130, x74129, x71989);
  nand n74132(x74132, x68462, x74134);
  nand n74133(x74133, x74132, x71994);
  nand n74135(x74135, x68462, x74137);
  nand n74136(x74136, x74135, x71999);
  nand n74138(x74138, x68462, x74140);
  nand n74139(x74139, x74138, x72004);
  nand n74141(x74141, x68462, x74143);
  nand n74142(x74142, x74141, x72009);
  nand n74144(x74144, x68462, x74146);
  nand n74145(x74145, x74144, x72014);
  nand n74147(x74147, x68462, x74149);
  nand n74148(x74148, x74147, x72019);
  nand n74150(x74150, x68462, x74152);
  nand n74151(x74151, x74150, x72024);
  nand n74153(x74153, x68462, x74155);
  nand n74154(x74154, x74153, x72029);
  nand n74156(x74156, x68462, x74158);
  nand n74157(x74157, x74156, x72034);
  nand n74159(x74159, x68462, x74161);
  nand n74160(x74160, x74159, x72039);
  nand n74162(x74162, x68462, x74164);
  nand n74163(x74163, x74162, x72044);
  nand n74165(x74165, x68462, x74167);
  nand n74166(x74166, x74165, x72049);
  nand n74168(x74168, x68462, x74170);
  nand n74169(x74169, x74168, x72054);
  nand n74171(x74171, x68462, x74173);
  nand n74172(x74172, x74171, x72059);
  nand n74174(x74174, x68462, x74176);
  nand n74175(x74175, x74174, x72064);
  nand n74177(x74177, x68462, x74179);
  nand n74178(x74178, x74177, x72069);
  nand n74180(x74180, x68462, x74182);
  nand n74181(x74181, x74180, x72074);
  nand n74183(x74183, x68462, x74185);
  nand n74184(x74184, x74183, x72079);
  nand n74186(x74186, x68462, x74188);
  nand n74187(x74187, x74186, x72084);
  nand n74189(x74189, x68462, x74191);
  nand n74190(x74190, x74189, x72089);
  nand n74192(x74192, x68462, x74194);
  nand n74193(x74193, x74192, x72094);
  nand n74195(x74195, x68462, x74197);
  nand n74196(x74196, x74195, x72099);
  nand n74198(x74198, x68462, x74200);
  nand n74199(x74199, x74198, x72104);
  nand n74201(x74201, x68462, x74203);
  nand n74202(x74202, x74201, x72109);
  nand n74204(x74204, x68462, x74206);
  nand n74205(x74205, x74204, x72114);
  nand n74207(x74207, x68462, x74209);
  nand n74208(x74208, x74207, x72119);
  nand n74210(x74210, x68462, x74212);
  nand n74211(x74211, x74210, x72124);
  nand n74213(x74213, x68462, x74215);
  nand n74214(x74214, x74213, x72129);
  nand n74216(x74216, x68462, x74218);
  nand n74217(x74217, x74216, x72134);
  nand n74219(x74219, x68462, x74221);
  nand n74220(x74220, x74219, x72139);
  nand n74222(x74222, x68462, x74224);
  nand n74223(x74223, x74222, x72144);
  nand n74225(x74225, x68462, x74227);
  nand n74226(x74226, x74225, x72149);
  nand n74228(x74228, x68462, x74230);
  nand n74229(x74229, x74228, x72154);
  nand n74231(x74231, x68462, x74233);
  nand n74232(x74232, x74231, x72159);
  nand n74234(x74234, x68462, x74236);
  nand n74235(x74235, x74234, x72164);
  nand n74237(x74237, x68462, x74239);
  nand n74238(x74238, x74237, x72169);
  nand n74240(x74240, x68462, x74242);
  nand n74241(x74241, x74240, x72174);
  nand n74243(x74243, x68462, x74245);
  nand n74244(x74244, x74243, x72179);
  nand n74246(x74246, x68462, x74248);
  nand n74247(x74247, x74246, x72184);
  nand n74249(x74249, x68462, x74251);
  nand n74250(x74250, x74249, x72189);
  nand n74252(x74252, x68462, x74254);
  nand n74253(x74253, x74252, x72194);
  nand n74255(x74255, x68462, x74257);
  nand n74256(x74256, x74255, x72199);
  nand n74258(x74258, x68462, x74260);
  nand n74259(x74259, x74258, x72204);
  nand n74261(x74261, x68462, x74263);
  nand n74262(x74262, x74261, x72209);
  nand n74264(x74264, x68462, x74266);
  nand n74265(x74265, x74264, x72214);
  nand n74267(x74267, x68462, x74269);
  nand n74268(x74268, x74267, x72219);
  nand n74270(x74270, x68462, x74272);
  nand n74271(x74271, x74270, x72224);
  nand n74273(x74273, x68462, x74275);
  nand n74274(x74274, x74273, x72229);
  nand n74276(x74276, x68462, x74278);
  nand n74277(x74277, x74276, x72234);
  nand n74279(x74279, x68462, x74281);
  nand n74280(x74280, x74279, x72239);
  nand n74282(x74282, x68462, x74284);
  nand n74283(x74283, x74282, x72244);
  nand n74285(x74285, x68462, x74287);
  nand n74286(x74286, x74285, x72249);
  nand n74288(x74288, x68462, x74290);
  nand n74289(x74289, x74288, x72254);
  nand n74291(x74291, x68462, x74293);
  nand n74292(x74292, x74291, x72259);
  nand n74294(x74294, x68462, x74296);
  nand n74295(x74295, x74294, x72264);
  nand n74297(x74297, x68462, x74299);
  nand n74298(x74298, x74297, x72269);
  nand n74300(x74300, x68462, x74302);
  nand n74301(x74301, x74300, x72274);
  nand n74303(x74303, x68462, x74305);
  nand n74304(x74304, x74303, x72279);
  nand n74306(x74306, x68462, x74308);
  nand n74307(x74307, x74306, x72284);
  nand n74309(x74309, x68462, x74311);
  nand n74310(x74310, x74309, x72289);
  nand n74312(x74312, x68462, x74314);
  nand n74313(x74313, x74312, x72294);
  nand n74315(x74315, x68462, x74317);
  nand n74316(x74316, x74315, x72299);
  nand n74318(x74318, x68462, x74320);
  nand n74319(x74319, x74318, x72304);
  nand n74321(x74321, x68462, x74323);
  nand n74322(x74322, x74321, x72309);
  nand n74324(x74324, x68462, x74326);
  nand n74325(x74325, x74324, x72314);
  nand n74327(x74327, x68462, x74329);
  nand n74328(x74328, x74327, x72319);
  nand n74330(x74330, x68462, x74332);
  nand n74331(x74331, x74330, x72324);
  nand n74333(x74333, x68462, x74335);
  nand n74334(x74334, x74333, x72329);
  nand n74336(x74336, x68462, x74338);
  nand n74337(x74337, x74336, x72334);
  nand n74339(x74339, x68462, x74341);
  nand n74340(x74340, x74339, x72339);
  nand n74342(x74342, x68462, x74344);
  nand n74343(x74343, x74342, x72344);
  nand n74345(x74345, x68462, x74347);
  nand n74346(x74346, x74345, x72349);
  nand n74348(x74348, x68462, x74350);
  nand n74349(x74349, x74348, x72354);
  nand n74351(x74351, x68462, x74353);
  nand n74352(x74352, x74351, x72359);
  nand n74354(x74354, x68462, x74356);
  nand n74355(x74355, x74354, x72364);
  nand n74357(x74357, x68462, x74359);
  nand n74358(x74358, x74357, x72369);
  nand n74360(x74360, x68462, x74362);
  nand n74361(x74361, x74360, x72374);
  nand n74363(x74363, x68462, x74365);
  nand n74364(x74364, x74363, x72379);
  nand n74366(x74366, x68462, x74368);
  nand n74367(x74367, x74366, x72384);
  nand n74369(x74369, x68462, x74371);
  nand n74370(x74370, x74369, x72389);
  nand n74372(x74372, x68462, x74374);
  nand n74373(x74373, x74372, x72394);
  nand n74375(x74375, x68462, x74377);
  nand n74376(x74376, x74375, x72399);
  nand n74378(x74378, x68462, x74380);
  nand n74379(x74379, x74378, x72404);
  nand n74381(x74381, x68462, x74383);
  nand n74382(x74382, x74381, x72409);
  nand n74384(x74384, x68462, x74386);
  nand n74385(x74385, x74384, x72414);
  nand n74387(x74387, x68462, x74389);
  nand n74388(x74388, x74387, x72419);
  nand n74390(x74390, x68462, x74392);
  nand n74391(x74391, x74390, x72424);
  nand n74393(x74393, x68462, x74395);
  nand n74394(x74394, x74393, x72429);
  nand n74396(x74396, x68462, x74398);
  nand n74397(x74397, x74396, x72434);
  nand n74399(x74399, x68462, x74401);
  nand n74400(x74400, x74399, x72439);
  nand n74402(x74402, x68462, x74404);
  nand n74403(x74403, x74402, x72444);
  nand n74405(x74405, x68462, x74407);
  nand n74406(x74406, x74405, x72449);
  nand n74408(x74408, x68462, x74410);
  nand n74409(x74409, x74408, x72454);
  nand n74411(x74411, x68462, x74413);
  nand n74412(x74412, x74411, x72459);
  nand n74414(x74414, x68462, x74416);
  nand n74415(x74415, x74414, x72464);
  nand n74417(x74417, x68462, x74419);
  nand n74418(x74418, x74417, x72469);
  nand n74420(x74420, x68462, x74422);
  nand n74421(x74421, x74420, x72474);
  nand n74423(x74423, x68462, x74425);
  nand n74424(x74424, x74423, x72479);
  nand n74426(x74426, x68462, x74428);
  nand n74427(x74427, x74426, x72484);
  nand n74429(x74429, x68462, x74431);
  nand n74430(x74430, x74429, x72489);
  nand n74432(x74432, x68462, x74434);
  nand n74433(x74433, x74432, x72494);
  nand n74435(x74435, x68462, x74437);
  nand n74436(x74436, x74435, x72499);
  nand n74438(x74438, x68462, x74440);
  nand n74439(x74439, x74438, x72504);
  nand n74441(x74441, x68462, x74443);
  nand n74442(x74442, x74441, x72509);
  nand n74444(x74444, x68462, x74446);
  nand n74445(x74445, x74444, x72514);
  nand n74447(x74447, x68462, x74449);
  nand n74448(x74448, x74447, x72519);
  nand n74450(x74450, x68462, x74452);
  nand n74451(x74451, x74450, x72524);
  nand n74453(x74453, x68462, x74455);
  nand n74454(x74454, x74453, x72529);
  nand n74456(x74456, x68462, x74458);
  nand n74457(x74457, x74456, x72534);
  nand n74459(x74459, x68462, x74461);
  nand n74460(x74460, x74459, x72539);
  nand n74462(x74462, x68462, x74464);
  nand n74463(x74463, x74462, x72544);
  nand n74465(x74465, x68462, x74467);
  nand n74466(x74466, x74465, x72549);
  nand n74468(x74468, x68462, x74470);
  nand n74469(x74469, x74468, x72554);
  nand n74471(x74471, x68462, x74473);
  nand n74472(x74472, x74471, x72559);
  nand n74474(x74474, x68462, x74476);
  nand n74475(x74475, x74474, x72564);
  nand n74477(x74477, x68462, x74479);
  nand n74478(x74478, x74477, x72569);
  nand n74480(x74480, x68462, x74482);
  nand n74481(x74481, x74480, x72574);
  nand n74483(x74483, x68462, x74485);
  nand n74484(x74484, x74483, x72579);
  nand n74486(x74486, x68462, x74488);
  nand n74487(x74487, x74486, x72584);
  nand n74489(x74489, x68462, x74491);
  nand n74490(x74490, x74489, x72589);
  nand n74492(x74492, x68462, x74494);
  nand n74493(x74493, x74492, x72594);
  nand n74495(x74495, x68462, x74497);
  nand n74496(x74496, x74495, x72599);
  nand n74498(x74498, x68462, x74500);
  nand n74499(x74499, x74498, x72604);
  nand n74501(x74501, x68462, x74503);
  nand n74502(x74502, x74501, x72609);
  nand n74504(x74504, x68462, x74506);
  nand n74505(x74505, x74504, x72614);
  nand n74507(x74507, x68462, x74509);
  nand n74508(x74508, x74507, x72619);
  nand n74510(x74510, x68462, x74512);
  nand n74511(x74511, x74510, x72624);
  nand n74513(x74513, x68462, x74515);
  nand n74514(x74514, x74513, x72629);
  nand n74516(x74516, x68462, x74518);
  nand n74517(x74517, x74516, x72634);
  nand n74519(x74519, x68462, x74521);
  nand n74520(x74520, x74519, x72639);
  nand n74522(x74522, x68462, x74524);
  nand n74523(x74523, x74522, x72644);
  nand n74525(x74525, x68462, x74527);
  nand n74526(x74526, x74525, x72649);
  nand n74528(x74528, x68462, x74530);
  nand n74529(x74529, x74528, x72654);
  nand n74531(x74531, x68462, x74533);
  nand n74532(x74532, x74531, x72659);
  nand n74534(x74534, x68462, x74536);
  nand n74535(x74535, x74534, x72664);
  nand n74537(x74537, x68462, x74539);
  nand n74538(x74538, x74537, x72669);
  nand n74540(x74540, x68462, x74542);
  nand n74541(x74541, x74540, x72674);
  nand n74543(x74543, x68462, x74545);
  nand n74544(x74544, x74543, x72679);
  nand n74546(x74546, x68462, x74548);
  nand n74547(x74547, x74546, x72684);
  nand n74549(x74549, x68462, x74551);
  nand n74550(x74550, x74549, x72689);
  nand n74552(x74552, x68462, x74554);
  nand n74553(x74553, x74552, x72694);
  nand n74555(x74555, x68462, x74557);
  nand n74556(x74556, x74555, x72699);
  nand n74558(x74558, x68462, x74560);
  nand n74559(x74559, x74558, x72704);
  nand n74561(x74561, x68462, x74563);
  nand n74562(x74562, x74561, x72709);
  nand n74564(x74564, x68462, x74566);
  nand n74565(x74565, x74564, x72714);
  nand n74567(x74567, x68462, x74569);
  nand n74568(x74568, x74567, x72719);
  nand n74570(x74570, x68462, x74572);
  nand n74571(x74571, x74570, x72724);
  nand n74573(x74573, x68462, x74575);
  nand n74574(x74574, x74573, x72729);
  nand n74576(x74576, x68462, x74578);
  nand n74577(x74577, x74576, x72734);
  nand n74579(x74579, x68462, x74581);
  nand n74580(x74580, x74579, x72739);
  nand n74582(x74582, x68462, x74584);
  nand n74583(x74583, x74582, x72744);
  nand n74585(x74585, x68462, x74587);
  nand n74586(x74586, x74585, x72749);
  nand n74588(x74588, x68462, x74590);
  nand n74589(x74589, x74588, x72754);
  nand n74591(x74591, x68462, x74593);
  nand n74592(x74592, x74591, x72759);
  nand n74594(x74594, x68462, x74596);
  nand n74595(x74595, x74594, x72764);
  nand n74597(x74597, x68462, x74599);
  nand n74598(x74598, x74597, x72769);
  nand n74600(x74600, x68462, x74602);
  nand n74601(x74601, x74600, x72774);
  nand n74603(x74603, x68462, x74605);
  nand n74604(x74604, x74603, x72779);
  nand n74606(x74606, x68462, x74608);
  nand n74607(x74607, x74606, x72784);
  nand n74609(x74609, x68462, x74611);
  nand n74610(x74610, x74609, x72789);
  nand n74612(x74612, x68462, x74614);
  nand n74613(x74613, x74612, x72794);
  nand n74615(x74615, x68462, x74617);
  nand n74616(x74616, x74615, x72799);
  nand n74618(x74618, x68462, x74620);
  nand n74619(x74619, x74618, x72804);
  nand n74621(x74621, x68462, x74623);
  nand n74622(x74622, x74621, x72809);
  nand n74624(x74624, x68462, x74626);
  nand n74625(x74625, x74624, x72814);
  nand n74627(x74627, x68462, x74629);
  nand n74628(x74628, x74627, x72819);
  nand n74630(x74630, x68462, x74632);
  nand n74631(x74631, x74630, x72824);
  nand n74633(x74633, x68462, x74635);
  nand n74634(x74634, x74633, x72829);
  nand n74636(x74636, x68462, x74638);
  nand n74637(x74637, x74636, x72834);
  nand n74639(x74639, x68462, x74641);
  nand n74640(x74640, x74639, x72839);
  nand n74642(x74642, x68462, x74644);
  nand n74643(x74643, x74642, x72844);
  nand n74645(x74645, x68462, x74647);
  nand n74646(x74646, x74645, x72849);
  nand n74648(x74648, x68462, x74650);
  nand n74649(x74649, x74648, x72854);
  nand n74651(x74651, x68462, x74653);
  nand n74652(x74652, x74651, x72859);
  nand n74654(x74654, x68462, x74656);
  nand n74655(x74655, x74654, x72864);
  nand n74657(x74657, x68462, x74659);
  nand n74658(x74658, x74657, x72869);
  nand n74660(x74660, x68462, x74662);
  nand n74661(x74661, x74660, x72874);
  nand n74663(x74663, x68462, x74665);
  nand n74664(x74664, x74663, x72879);
  nand n74666(x74666, x68462, x74668);
  nand n74667(x74667, x74666, x72884);
  nand n74669(x74669, x68462, x74671);
  nand n74670(x74670, x74669, x72889);
  nand n74672(x74672, x68462, x74674);
  nand n74673(x74673, x74672, x72894);
  nand n74675(x74675, x68462, x74677);
  nand n74676(x74676, x74675, x72899);
  nand n74678(x74678, x68462, x74680);
  nand n74679(x74679, x74678, x72904);
  nand n74681(x74681, x68462, x74683);
  nand n74682(x74682, x74681, x72909);
  nand n74684(x74684, x68462, x74686);
  nand n74685(x74685, x74684, x72914);
  nand n74687(x74687, x68462, x74689);
  nand n74688(x74688, x74687, x72919);
  nand n74690(x74690, x68462, x74692);
  nand n74691(x74691, x74690, x72924);
  nand n74693(x74693, x68462, x74695);
  nand n74694(x74694, x74693, x72929);
  nand n74696(x74696, x68462, x74698);
  nand n74697(x74697, x74696, x72934);
  nand n74699(x74699, x68462, x74701);
  nand n74700(x74700, x74699, x72939);
  nand n74702(x74702, x68462, x74704);
  nand n74703(x74703, x74702, x72944);
  nand n74705(x74705, x68462, x74707);
  nand n74706(x74706, x74705, x72949);
  nand n74708(x74708, x68462, x74710);
  nand n74709(x74709, x74708, x72954);
  nand n74711(x74711, x68462, x74713);
  nand n74712(x74712, x74711, x72959);
  nand n74714(x74714, x68462, x74716);
  nand n74715(x74715, x74714, x72964);
  nand n74717(x74717, x68462, x74719);
  nand n74718(x74718, x74717, x72969);
  nand n74720(x74720, x68462, x74722);
  nand n74721(x74721, x74720, x72974);
  nand n74723(x74723, x68462, x74725);
  nand n74724(x74724, x74723, x72979);
  nand n74726(x74726, x68462, x74728);
  nand n74727(x74727, x74726, x72984);
  nand n74729(x74729, x68462, x74731);
  nand n74730(x74730, x74729, x72989);
  nand n74732(x74732, x68462, x74734);
  nand n74733(x74733, x74732, x72994);
  nand n74735(x74735, x68462, x74737);
  nand n74736(x74736, x74735, x72999);
  nand n74738(x74738, x68462, x74740);
  nand n74739(x74739, x74738, x73004);
  nand n74741(x74741, x68462, x74743);
  nand n74742(x74742, x74741, x73009);
  nand n74744(x74744, x68462, x74746);
  nand n74745(x74745, x74744, x73014);
  nand n74747(x74747, x68462, x74749);
  nand n74748(x74748, x74747, x73019);
  nand n74750(x74750, x68462, x74752);
  nand n74751(x74751, x74750, x73024);
  nand n74753(x74753, x68462, x74755);
  nand n74754(x74754, x74753, x73029);
  nand n74756(x74756, x68462, x74758);
  nand n74757(x74757, x74756, x73034);
  nand n74759(x74759, x68462, x74761);
  nand n74760(x74760, x74759, x73039);
  nand n74762(x74762, x68462, x74764);
  nand n74763(x74763, x74762, x73044);
  nand n74765(x74765, x68462, x74767);
  nand n74766(x74766, x74765, x73049);
  nand n74768(x74768, x68462, x74770);
  nand n74769(x74769, x74768, x73054);
  nand n74771(x74771, x68462, x74773);
  nand n74772(x74772, x74771, x73059);
  nand n74774(x74774, x68462, x74776);
  nand n74775(x74775, x74774, x73064);
  nand n74777(x74777, x68462, x74779);
  nand n74778(x74778, x74777, x73069);
  nand n74780(x74780, x68462, x74782);
  nand n74781(x74781, x74780, x73074);
  nand n74783(x74783, x68462, x74785);
  nand n74784(x74784, x74783, x73079);
  nand n74786(x74786, x68462, x74788);
  nand n74787(x74787, x74786, x73084);
  nand n74789(x74789, x68462, x74791);
  nand n74790(x74790, x74789, x73089);
  nand n74792(x74792, x68462, x74794);
  nand n74793(x74793, x74792, x73094);
  nand n74795(x74795, x68462, x74797);
  nand n74796(x74796, x74795, x73099);
  nand n74798(x74798, x68462, x74800);
  nand n74799(x74799, x74798, x73104);
  nand n74801(x74801, x68462, x74803);
  nand n74802(x74802, x74801, x73109);
  nand n74804(x74804, x68462, x74806);
  nand n74805(x74805, x74804, x73114);
  nand n74807(x74807, x68462, x74809);
  nand n74808(x74808, x74807, x73119);
  nand n74810(x74810, x68462, x74812);
  nand n74811(x74811, x74810, x73124);
  nand n74813(x74813, x68462, x74815);
  nand n74814(x74814, x74813, x73129);
  nand n74816(x74816, x68462, x74818);
  nand n74817(x74817, x74816, x73134);
  nand n74819(x74819, x68462, x74821);
  nand n74820(x74820, x74819, x73139);
  nand n74822(x74822, x68462, x74824);
  nand n74823(x74823, x74822, x73144);
  nand n74825(x74825, x68462, x74827);
  nand n74826(x74826, x74825, x73149);
  nand n74828(x74828, x68462, x74830);
  nand n74829(x74829, x74828, x73154);
  nand n74831(x74831, x68462, x74833);
  nand n74832(x74832, x74831, x73159);
  nand n74834(x74834, x68462, x74836);
  nand n74835(x74835, x74834, x73164);
  nand n74837(x74837, x68462, x74839);
  nand n74838(x74838, x74837, x73169);
  nand n74840(x74840, x68462, x74842);
  nand n74841(x74841, x74840, x73174);
  nand n74843(x74843, x68462, x74845);
  nand n74844(x74844, x74843, x73179);
  nand n74846(x74846, x68462, x74848);
  nand n74847(x74847, x74846, x73184);
  nand n74849(x74849, x68462, x74851);
  nand n74850(x74850, x74849, x73189);
  nand n74852(x74852, x68462, x74854);
  nand n74853(x74853, x74852, x73194);
  nand n74855(x74855, x68462, x74857);
  nand n74856(x74856, x74855, x73199);
  nand n74858(x74858, x68462, x74860);
  nand n74859(x74859, x74858, x73204);
  nand n74861(x74861, x68462, x74863);
  nand n74862(x74862, x74861, x73209);
  nand n74864(x74864, x68462, x74866);
  nand n74865(x74865, x74864, x73214);
  nand n74867(x74867, x68462, x74869);
  nand n74868(x74868, x74867, x73219);
  nand n74870(x74870, x68462, x74872);
  nand n74871(x74871, x74870, x73224);
  nand n74873(x74873, x68462, x74875);
  nand n74874(x74874, x74873, x73229);
  nand n74876(x74876, x68462, x74878);
  nand n74877(x74877, x74876, x73234);
  nand n74879(x74879, x68462, x74881);
  nand n74880(x74880, x74879, x73239);
  nand n74882(x74882, x68462, x74884);
  nand n74883(x74883, x74882, x73244);
  nand n74885(x74885, x68462, x74887);
  nand n74886(x74886, x74885, x73249);
  nand n74888(x74888, x68462, x74890);
  nand n74889(x74889, x74888, x73254);
  nand n74891(x74891, x68462, x74893);
  nand n74892(x74892, x74891, x73259);
  nand n74894(x74894, x68462, x74896);
  nand n74895(x74895, x74894, x73264);
  nand n74897(x74897, x68462, x74899);
  nand n74898(x74898, x74897, x73269);
  nand n74900(x74900, x68462, x74902);
  nand n74901(x74901, x74900, x73274);
  nand n74903(x74903, x68462, x74905);
  nand n74904(x74904, x74903, x73279);
  nand n74906(x74906, x68462, x74908);
  nand n74907(x74907, x74906, x73284);
  nand n74909(x74909, x68462, x74911);
  nand n74910(x74910, x74909, x73289);
  nand n74912(x74912, x68462, x74914);
  nand n74913(x74913, x74912, x73294);
  nand n74915(x74915, x68462, x74917);
  nand n74916(x74916, x74915, x73299);
  nand n74918(x74918, x68462, x74920);
  nand n74919(x74919, x74918, x73304);
  nand n74921(x74921, x68462, x74923);
  nand n74922(x74922, x74921, x73309);
  nand n74924(x74924, x68462, x74926);
  nand n74925(x74925, x74924, x73314);
  nand n74927(x74927, x68462, x74929);
  nand n74928(x74928, x74927, x73319);
  nand n74930(x74930, x68462, x74932);
  nand n74931(x74931, x74930, x73324);
  nand n74933(x74933, x68462, x74935);
  nand n74934(x74934, x74933, x73329);
  nand n74936(x74936, x68462, x74938);
  nand n74937(x74937, x74936, x73334);
  nand n74939(x74939, x68462, x74941);
  nand n74940(x74940, x74939, x73339);
  nand n74942(x74942, x68462, x74944);
  nand n74943(x74943, x74942, x73344);
  nand n74945(x74945, x68462, x74947);
  nand n74946(x74946, x74945, x73349);
  nand n74948(x74948, x68462, x74950);
  nand n74949(x74949, x74948, x73354);
  nand n74951(x74951, x68462, x74953);
  nand n74952(x74952, x74951, x73359);
  nand n74954(x74954, x68462, x74956);
  nand n74955(x74955, x74954, x73364);
  nand n74957(x74957, x68462, x74959);
  nand n74958(x74958, x74957, x73369);
  nand n74960(x74960, x68462, x74962);
  nand n74961(x74961, x74960, x73374);
  nand n74963(x74963, x68462, x74965);
  nand n74964(x74964, x74963, x73379);
  nand n74966(x74966, x68462, x74968);
  nand n74967(x74967, x74966, x73384);
  nand n74969(x74969, x68462, x74971);
  nand n74970(x74970, x74969, x73389);
  nand n74972(x74972, x68462, x74974);
  nand n74973(x74973, x74972, x73394);
  nand n74975(x74975, x68462, x74977);
  nand n74976(x74976, x74975, x73399);
  nand n74978(x74978, x68462, x74980);
  nand n74979(x74979, x74978, x73404);
  nand n74981(x74981, x68462, x74983);
  nand n74982(x74982, x74981, x73409);
  nand n74984(x74984, x68462, x74986);
  nand n74985(x74985, x74984, x73414);
  nand n74987(x74987, x68462, x74989);
  nand n74988(x74988, x74987, x73419);
  nand n74990(x74990, x68462, x74992);
  nand n74991(x74991, x74990, x73424);
  nand n74993(x74993, x68462, x74995);
  nand n74994(x74994, x74993, x73429);
  nand n74996(x74996, x68462, x74998);
  nand n74997(x74997, x74996, x73434);
  nand n74999(x74999, x68462, x75001);
  nand n75000(x75000, x74999, x73439);
  nand n75002(x75002, x68462, x75004);
  nand n75003(x75003, x75002, x73444);
  nand n75005(x75005, x68462, x75007);
  nand n75006(x75006, x75005, x73449);
  nand n75008(x75008, x68462, x75010);
  nand n75009(x75009, x75008, x73454);
  nand n75011(x75011, x68462, x75013);
  nand n75012(x75012, x75011, x73459);
  nand n75014(x75014, x68462, x75016);
  nand n75015(x75015, x75014, x73464);
  nand n75017(x75017, x68462, x75019);
  nand n75018(x75018, x75017, x73469);
  nand n75020(x75020, x68462, x75022);
  nand n75021(x75021, x75020, x73474);
  nand n75023(x75023, x68462, x75025);
  nand n75024(x75024, x75023, x73479);
  nand n75026(x75026, x68462, x75028);
  nand n75027(x75027, x75026, x73484);
  nand n75029(x75029, x68462, x75031);
  nand n75030(x75030, x75029, x73489);
  nand n75032(x75032, x68462, x75034);
  nand n75033(x75033, x75032, x73494);
  nand n75035(x75035, x68462, x75037);
  nand n75036(x75036, x75035, x73499);
  nand n75038(x75038, x68462, x75040);
  nand n75039(x75039, x75038, x73504);
  nand n75041(x75041, x68462, x75043);
  nand n75042(x75042, x75041, x73509);
  nand n75044(x75044, x68462, x75046);
  nand n75045(x75045, x75044, x73514);
  nand n75047(x75047, x68462, x75049);
  nand n75048(x75048, x75047, x73519);
  nand n75050(x75050, x68462, x75052);
  nand n75051(x75051, x75050, x73524);
  nand n75053(x75053, x68462, x75055);
  nand n75054(x75054, x75053, x73529);
  nand n75056(x75056, x68462, x75058);
  nand n75057(x75057, x75056, x73534);
  nand n75059(x75059, x68462, x75061);
  nand n75060(x75060, x75059, x73539);
  nand n75062(x75062, x68462, x75064);
  nand n75063(x75063, x75062, x73544);
  nand n75065(x75065, x68462, x75067);
  nand n75066(x75066, x75065, x73549);
  nand n75068(x75068, x68462, x75070);
  nand n75069(x75069, x75068, x73554);
  nand n75071(x75071, x68462, x75073);
  nand n75072(x75072, x75071, x73559);
  nand n75074(x75074, x68462, x75076);
  nand n75075(x75075, x75074, x73564);
  nand n75077(x75077, x68462, x75079);
  nand n75078(x75078, x75077, x73569);
  nand n75080(x75080, x68462, x75082);
  nand n75081(x75081, x75080, x73574);
  nand n75083(x75083, x68462, x75085);
  nand n75084(x75084, x75083, x73579);
  nand n75086(x75086, x68462, x75088);
  nand n75087(x75087, x75086, x73584);
  nand n75089(x75089, x68462, x75091);
  nand n75090(x75090, x75089, x73589);
  nand n75092(x75092, x68462, x75094);
  nand n75093(x75093, x75092, x73594);
  nand n75095(x75095, x68462, x75097);
  nand n75096(x75096, x75095, x73599);
  nand n75098(x75098, x68462, x75100);
  nand n75099(x75099, x75098, x73604);
  nand n75101(x75101, x68462, x75103);
  nand n75102(x75102, x75101, x73609);
  nand n75104(x75104, x68462, x75106);
  nand n75105(x75105, x75104, x73614);
  nand n75107(x75107, x68462, x75109);
  nand n75108(x75108, x75107, x73619);
  nand n75110(x75110, x68462, x75112);
  nand n75111(x75111, x75110, x73624);
  nand n75113(x75113, x68462, x75115);
  nand n75114(x75114, x75113, x73629);
  nand n75116(x75116, x68462, x75118);
  nand n75117(x75117, x75116, x73634);
  nand n75119(x75119, x68462, x75121);
  nand n75120(x75120, x75119, x73639);
  nand n75122(x75122, x68462, x75124);
  nand n75123(x75123, x75122, x73644);
  nand n75125(x75125, x68462, x75127);
  nand n75126(x75126, x75125, x73649);
  nand n75128(x75128, x68462, x75130);
  nand n75129(x75129, x75128, x73654);
  nand n75131(x75131, x68462, x75133);
  nand n75132(x75132, x75131, x73659);
  nand n75134(x75134, x68462, x75136);
  nand n75135(x75135, x75134, x73664);
  nand n75137(x75137, x68462, x75139);
  nand n75138(x75138, x75137, x73669);
  nand n75140(x75140, x68462, x75142);
  nand n75141(x75141, x75140, x73674);
  nand n75143(x75143, x68462, x75145);
  nand n75144(x75144, x75143, x73679);
  nand n75146(x75146, x68462, x75148);
  nand n75147(x75147, x75146, x73684);
  nand n75149(x75149, x68462, x75151);
  nand n75150(x75150, x75149, x73689);
  nand n75152(x75152, x68462, x75154);
  nand n75153(x75153, x75152, x73694);
  nand n75155(x75155, x68462, x75157);
  nand n75156(x75156, x75155, x73699);
  nand n75158(x75158, x68462, x75160);
  nand n75159(x75159, x75158, x73704);
  nand n75161(x75161, x68462, x75163);
  nand n75162(x75162, x75161, x73709);
  nand n75164(x75164, x68462, x75166);
  nand n75165(x75165, x75164, x73714);
  nand n75167(x75167, x68462, x75169);
  nand n75168(x75168, x75167, x73719);
  nand n75170(x75170, x68462, x75172);
  nand n75171(x75171, x75170, x73724);
  nand n75173(x75173, x68462, x75175);
  nand n75174(x75174, x75173, x73729);
  nand n75176(x75176, x68462, x75178);
  nand n75177(x75177, x75176, x73734);
  nand n75179(x75179, x68462, x75181);
  nand n75180(x75180, x75179, x73739);
  nand n75182(x75182, x68462, x75184);
  nand n75183(x75183, x75182, x73744);
  nand n75185(x75185, x68462, x75187);
  nand n75186(x75186, x75185, x73749);
  nand n75188(x75188, x68462, x75190);
  nand n75189(x75189, x75188, x73754);
  nand n75191(x75191, x68462, x75193);
  nand n75192(x75192, x75191, x73759);
  nand n75194(x75194, x68462, x75196);
  nand n75195(x75195, x75194, x73764);
  nand n75197(x75197, x68462, x75199);
  nand n75198(x75198, x75197, x73769);
  nand n75200(x75200, x68462, x75202);
  nand n75201(x75201, x75200, x73774);
  nand n75203(x75203, x68462, x75205);
  nand n75204(x75204, x75203, x73779);
  nand n75206(x75206, x68462, x75208);
  nand n75207(x75207, x75206, x73784);
  nand n75209(x75209, x68462, x75211);
  nand n75210(x75210, x75209, x73789);
  nand n75212(x75212, x68462, x75214);
  nand n75213(x75213, x75212, x73794);
  nand n75215(x75215, x68462, x75217);
  nand n75216(x75216, x75215, x73799);
  nand n75218(x75218, x68462, x75220);
  nand n75219(x75219, x75218, x73804);
  nand n75221(x75221, x68462, x75223);
  nand n75222(x75222, x75221, x73809);
  nand n75224(x75224, x68462, x75226);
  nand n75225(x75225, x75224, x73814);
  nand n75227(x75227, x68462, x75229);
  nand n75228(x75228, x75227, x73819);
  nand n75230(x75230, x68462, x75232);
  nand n75231(x75231, x75230, x73824);
  nand n75233(x75233, x68462, x75235);
  nand n75234(x75234, x75233, x73829);
  nand n75236(x75236, x68462, x75238);
  nand n75237(x75237, x75236, x73834);
  nand n75239(x75239, x68462, x75241);
  nand n75240(x75240, x75239, x73839);
  nand n75242(x75242, x68462, x75244);
  nand n75243(x75243, x75242, x73844);
  nand n75245(x75245, x68462, x75247);
  nand n75246(x75246, x75245, x73849);
  nand n75248(x75248, x68462, x75250);
  nand n75249(x75249, x75248, x73854);
  nand n75251(x75251, x68462, x75253);
  nand n75252(x75252, x75251, x73859);
  nand n75254(x75254, x68462, x75256);
  nand n75255(x75255, x75254, x73864);
  nand n75257(x75257, x68462, x75259);
  nand n75258(x75258, x75257, x73869);
  nand n75260(x75260, x68462, x75262);
  nand n75261(x75261, x75260, x73874);
  nand n75263(x75263, x68462, x75265);
  nand n75264(x75264, x75263, x73879);
  nand n75266(x75266, x68462, x75268);
  nand n75267(x75267, x75266, x73884);
  nand n75269(x75269, x68462, x75271);
  nand n75270(x75270, x75269, x73889);
  nand n75272(x75272, x68462, x75274);
  nand n75273(x75273, x75272, x73894);
  nand n75275(x75275, x68462, x75277);
  nand n75276(x75276, x75275, x73899);
  nand n75278(x75278, x68462, x75280);
  nand n75279(x75279, x75278, x73904);
  nand n75281(x75281, x68462, x75283);
  nand n75282(x75282, x75281, x73909);
  nand n75284(x75284, x68462, x75286);
  nand n75285(x75285, x75284, x73914);
  nand n75287(x75287, x68462, x75289);
  nand n75288(x75288, x75287, x73919);
  nand n75290(x75290, x68462, x75292);
  nand n75291(x75291, x75290, x73924);
  nand n75293(x75293, x68462, x75295);
  nand n75294(x75294, x75293, x73929);
  nand n75296(x75296, x68462, x75298);
  nand n75297(x75297, x75296, x73934);
  nand n75299(x75299, x68462, x75301);
  nand n75300(x75300, x75299, x73939);
  nand n75302(x75302, x68462, x75304);
  nand n75303(x75303, x75302, x73944);
  nand n75305(x75305, x68462, x75307);
  nand n75306(x75306, x75305, x73949);
  nand n75308(x75308, x68462, x75310);
  nand n75309(x75309, x75308, x73954);
  nand n75311(x75311, x68462, x75313);
  nand n75312(x75312, x75311, x73959);
  nand n75314(x75314, x68462, x75316);
  nand n75315(x75315, x75314, x73964);
  nand n75317(x75317, x68462, x75319);
  nand n75318(x75318, x75317, x73969);
  nand n75320(x75320, x68462, x75322);
  nand n75321(x75321, x75320, x73974);
  nand n75323(x75323, x68462, x75325);
  nand n75324(x75324, x75323, x73979);
  nand n75326(x75326, x68462, x75328);
  nand n75327(x75327, x75326, x73984);
  nand n75329(x75329, x68462, x75331);
  nand n75330(x75330, x75329, x73989);
  nand n75332(x75332, x68462, x75334);
  nand n75333(x75333, x75332, x73994);
  nand n75335(x75335, x68462, x75337);
  nand n75336(x75336, x75335, x73999);
  nand n75338(x75338, x68462, x75340);
  nand n75339(x75339, x75338, x71799);
  nand n75341(x75341, x68462, x75343);
  nand n75342(x75342, x75341, x71804);
  nand n75344(x75344, x68462, x75346);
  nand n75345(x75345, x75344, x71809);
  nand n75347(x75347, x68462, x75349);
  nand n75348(x75348, x75347, x71814);
  nand n75350(x75350, x68462, x75352);
  nand n75351(x75351, x75350, x71819);
  nand n75353(x75353, x68462, x75355);
  nand n75354(x75354, x75353, x71824);
  nand n75356(x75356, x68462, x75358);
  nand n75357(x75357, x75356, x71829);
  nand n75359(x75359, x68462, x75361);
  nand n75360(x75360, x75359, x71834);
  nand n75362(x75362, x68462, x75364);
  nand n75363(x75363, x75362, x71839);
  nand n75365(x75365, x68462, x75367);
  nand n75366(x75366, x75365, x71844);
  nand n75368(x75368, x68462, x75370);
  nand n75369(x75369, x75368, x71849);
  nand n75371(x75371, x68462, x75373);
  nand n75372(x75372, x75371, x71854);
  nand n75374(x75374, x68462, x75376);
  nand n75375(x75375, x75374, x71859);
  nand n75377(x75377, x68462, x75379);
  nand n75378(x75378, x75377, x71864);
  nand n75380(x75380, x68462, x75382);
  nand n75381(x75381, x75380, x71869);
  nand n75383(x75383, x68462, x75385);
  nand n75384(x75384, x75383, x71874);
  nand n75386(x75386, x68462, x75388);
  nand n75387(x75387, x75386, x71879);
  nand n75389(x75389, x68462, x75391);
  nand n75390(x75390, x75389, x71884);
  nand n75392(x75392, x68462, x75394);
  nand n75393(x75393, x75392, x71889);
  nand n75395(x75395, x68462, x75397);
  nand n75396(x75396, x75395, x71894);
  nand n75398(x75398, x68462, x75400);
  nand n75399(x75399, x75398, x71899);
  nand n75401(x75401, x68462, x75403);
  nand n75402(x75402, x75401, x71904);
  nand n75404(x75404, x68462, x75406);
  nand n75405(x75405, x75404, x71904);
  nand n75407(x75407, x68462, x75409);
  nand n75408(x75408, x75407, x71904);
  nand n75410(x75410, x68462, x75412);
  nand n75411(x75411, x75410, x71904);
  nand n75413(x75413, x68462, x75415);
  nand n75414(x75414, x75413, x71904);
  nand n75416(x75416, x68462, x75418);
  nand n75417(x75417, x75416, x71904);
  nand n75419(x75419, x68462, x75421);
  nand n75420(x75420, x75419, x71904);
  nand n75422(x75422, x68462, x75424);
  nand n75423(x75423, x75422, x71904);
  nand n75425(x75425, x68462, x75427);
  nand n75426(x75426, x75425, x71904);
  nand n75428(x75428, x68462, x75430);
  nand n75429(x75429, x75428, x71904);
  nand n75431(x75431, x68462, x75433);
  nand n75432(x75432, x75431, x71904);
  nand n75434(x75434, x68462, x75436);
  nand n75435(x75435, x75434, x71939);
  nand n75437(x75437, x68462, x75439);
  nand n75438(x75438, x75437, x71944);
  nand n75440(x75440, x68462, x75442);
  nand n75441(x75441, x75440, x71949);
  nand n75443(x75443, x68462, x75445);
  nand n75444(x75444, x75443, x71954);
  nand n75446(x75446, x68462, x75448);
  nand n75447(x75447, x75446, x71959);
  nand n75449(x75449, x68462, x75451);
  nand n75450(x75450, x75449, x71964);
  nand n75452(x75452, x68462, x75454);
  nand n75453(x75453, x75452, x71969);
  nand n75455(x75455, x68462, x75457);
  nand n75456(x75456, x75455, x71974);
  nand n75458(x75458, x68462, x75460);
  nand n75459(x75459, x75458, x71979);
  nand n75461(x75461, x68462, x75463);
  nand n75462(x75462, x75461, x71984);
  nand n75464(x75464, x68462, x75466);
  nand n75465(x75465, x75464, x71989);
  nand n75467(x75467, x68462, x75469);
  nand n75468(x75468, x75467, x71994);
  nand n75470(x75470, x68462, x75472);
  nand n75471(x75471, x75470, x71999);
  nand n75473(x75473, x68462, x75475);
  nand n75474(x75474, x75473, x72004);
  nand n75476(x75476, x68462, x75478);
  nand n75477(x75477, x75476, x72009);
  nand n75479(x75479, x68462, x75481);
  nand n75480(x75480, x75479, x72014);
  nand n75482(x75482, x68462, x75484);
  nand n75483(x75483, x75482, x72019);
  nand n75485(x75485, x68462, x75487);
  nand n75486(x75486, x75485, x72024);
  nand n75488(x75488, x68462, x75490);
  nand n75489(x75489, x75488, x72029);
  nand n75491(x75491, x68462, x75493);
  nand n75492(x75492, x75491, x72034);
  nand n75494(x75494, x68462, x75496);
  nand n75495(x75495, x75494, x72039);
  nand n75497(x75497, x68462, x75499);
  nand n75498(x75498, x75497, x72044);
  nand n75500(x75500, x68462, x75502);
  nand n75501(x75501, x75500, x72049);
  nand n75503(x75503, x68462, x75505);
  nand n75504(x75504, x75503, x72054);
  nand n75506(x75506, x68462, x75508);
  nand n75507(x75507, x75506, x72059);
  nand n75509(x75509, x68462, x75511);
  nand n75510(x75510, x75509, x72064);
  nand n75512(x75512, x68462, x75514);
  nand n75513(x75513, x75512, x72069);
  nand n75515(x75515, x68462, x75517);
  nand n75516(x75516, x75515, x72074);
  nand n75518(x75518, x68462, x75520);
  nand n75519(x75519, x75518, x72079);
  nand n75521(x75521, x68462, x75523);
  nand n75522(x75522, x75521, x72084);
  nand n75524(x75524, x68462, x75526);
  nand n75525(x75525, x75524, x72089);
  nand n75527(x75527, x68462, x75529);
  nand n75528(x75528, x75527, x72094);
  nand n75530(x75530, x68462, x75532);
  nand n75531(x75531, x75530, x72099);
  nand n75533(x75533, x68462, x75535);
  nand n75534(x75534, x75533, x72104);
  nand n75536(x75536, x68462, x75538);
  nand n75537(x75537, x75536, x72109);
  nand n75539(x75539, x68462, x75541);
  nand n75540(x75540, x75539, x72114);
  nand n75542(x75542, x68462, x75544);
  nand n75543(x75543, x75542, x72119);
  nand n75545(x75545, x68462, x75547);
  nand n75546(x75546, x75545, x72124);
  nand n75548(x75548, x68462, x75550);
  nand n75549(x75549, x75548, x72129);
  nand n75551(x75551, x68462, x75553);
  nand n75552(x75552, x75551, x72134);
  nand n75554(x75554, x68462, x75556);
  nand n75555(x75555, x75554, x72139);
  nand n75557(x75557, x68462, x75559);
  nand n75558(x75558, x75557, x72144);
  nand n75560(x75560, x68462, x75562);
  nand n75561(x75561, x75560, x72149);
  nand n75563(x75563, x68462, x75565);
  nand n75564(x75564, x75563, x72154);
  nand n75566(x75566, x68462, x75568);
  nand n75567(x75567, x75566, x72159);
  nand n75569(x75569, x68462, x75571);
  nand n75570(x75570, x75569, x72164);
  nand n75572(x75572, x68462, x75574);
  nand n75573(x75573, x75572, x72169);
  nand n75575(x75575, x68462, x75577);
  nand n75576(x75576, x75575, x72174);
  nand n75578(x75578, x68462, x75580);
  nand n75579(x75579, x75578, x72179);
  nand n75581(x75581, x68462, x75583);
  nand n75582(x75582, x75581, x72184);
  nand n75584(x75584, x68462, x75586);
  nand n75585(x75585, x75584, x72189);
  nand n75587(x75587, x68462, x75589);
  nand n75588(x75588, x75587, x72194);
  nand n75590(x75590, x68462, x75592);
  nand n75591(x75591, x75590, x72199);
  nand n75593(x75593, x68462, x75595);
  nand n75594(x75594, x75593, x72204);
  nand n75596(x75596, x68462, x75598);
  nand n75597(x75597, x75596, x72209);
  nand n75599(x75599, x68462, x75601);
  nand n75600(x75600, x75599, x72214);
  nand n75602(x75602, x68462, x75604);
  nand n75603(x75603, x75602, x72219);
  nand n75605(x75605, x68462, x75607);
  nand n75606(x75606, x75605, x72224);
  nand n75608(x75608, x68462, x75610);
  nand n75609(x75609, x75608, x72229);
  nand n75611(x75611, x68462, x75613);
  nand n75612(x75612, x75611, x72234);
  nand n75614(x75614, x68462, x75616);
  nand n75615(x75615, x75614, x72239);
  nand n75617(x75617, x68462, x75619);
  nand n75618(x75618, x75617, x72244);
  nand n75620(x75620, x68462, x75622);
  nand n75621(x75621, x75620, x72249);
  nand n75623(x75623, x68462, x75625);
  nand n75624(x75624, x75623, x72254);
  nand n75626(x75626, x68462, x75628);
  nand n75627(x75627, x75626, x72259);
  nand n75629(x75629, x68462, x75631);
  nand n75630(x75630, x75629, x72264);
  nand n75632(x75632, x68462, x75634);
  nand n75633(x75633, x75632, x72269);
  nand n75635(x75635, x68462, x75637);
  nand n75636(x75636, x75635, x72274);
  nand n75638(x75638, x68462, x75640);
  nand n75639(x75639, x75638, x72279);
  nand n75641(x75641, x68462, x75643);
  nand n75642(x75642, x75641, x72284);
  nand n75644(x75644, x68462, x75646);
  nand n75645(x75645, x75644, x72289);
  nand n75647(x75647, x68462, x75649);
  nand n75648(x75648, x75647, x72294);
  nand n75650(x75650, x68462, x75652);
  nand n75651(x75651, x75650, x72299);
  nand n75653(x75653, x68462, x75655);
  nand n75654(x75654, x75653, x72304);
  nand n75656(x75656, x68462, x75658);
  nand n75657(x75657, x75656, x72309);
  nand n75659(x75659, x68462, x75661);
  nand n75660(x75660, x75659, x72314);
  nand n75662(x75662, x68462, x75664);
  nand n75663(x75663, x75662, x72319);
  nand n75665(x75665, x68462, x75667);
  nand n75666(x75666, x75665, x72324);
  nand n75668(x75668, x68462, x75670);
  nand n75669(x75669, x75668, x72329);
  nand n75671(x75671, x68462, x75673);
  nand n75672(x75672, x75671, x72334);
  nand n75674(x75674, x68462, x75676);
  nand n75675(x75675, x75674, x72339);
  nand n75677(x75677, x68462, x75679);
  nand n75678(x75678, x75677, x72344);
  nand n75680(x75680, x68462, x75682);
  nand n75681(x75681, x75680, x72349);
  nand n75683(x75683, x68462, x75685);
  nand n75684(x75684, x75683, x72354);
  nand n75686(x75686, x68462, x75688);
  nand n75687(x75687, x75686, x72359);
  nand n75689(x75689, x68462, x75691);
  nand n75690(x75690, x75689, x72364);
  nand n75692(x75692, x68462, x75694);
  nand n75693(x75693, x75692, x72369);
  nand n75695(x75695, x68462, x75697);
  nand n75696(x75696, x75695, x72374);
  nand n75698(x75698, x68462, x75700);
  nand n75699(x75699, x75698, x72379);
  nand n75701(x75701, x68462, x75703);
  nand n75702(x75702, x75701, x72384);
  nand n75704(x75704, x68462, x75706);
  nand n75705(x75705, x75704, x72389);
  nand n75707(x75707, x68462, x75709);
  nand n75708(x75708, x75707, x72394);
  nand n75710(x75710, x68462, x75712);
  nand n75711(x75711, x75710, x72399);
  nand n75713(x75713, x68462, x75715);
  nand n75714(x75714, x75713, x72404);
  nand n75716(x75716, x68462, x75718);
  nand n75717(x75717, x75716, x72409);
  nand n75719(x75719, x68462, x75721);
  nand n75720(x75720, x75719, x72414);
  nand n75722(x75722, x68462, x75724);
  nand n75723(x75723, x75722, x72419);
  nand n75725(x75725, x68462, x75727);
  nand n75726(x75726, x75725, x72424);
  nand n75728(x75728, x68462, x75730);
  nand n75729(x75729, x75728, x72429);
  nand n75731(x75731, x68462, x75733);
  nand n75732(x75732, x75731, x72434);
  nand n75734(x75734, x68462, x75736);
  nand n75735(x75735, x75734, x72439);
  nand n75737(x75737, x68462, x75739);
  nand n75738(x75738, x75737, x72444);
  nand n75740(x75740, x68462, x75742);
  nand n75741(x75741, x75740, x72449);
  nand n75743(x75743, x68462, x75745);
  nand n75744(x75744, x75743, x72454);
  nand n75746(x75746, x68462, x75748);
  nand n75747(x75747, x75746, x72459);
  nand n75749(x75749, x68462, x75751);
  nand n75750(x75750, x75749, x72464);
  nand n75752(x75752, x68462, x75754);
  nand n75753(x75753, x75752, x72469);
  nand n75755(x75755, x68462, x75757);
  nand n75756(x75756, x75755, x72474);
  nand n75758(x75758, x68462, x75760);
  nand n75759(x75759, x75758, x72479);
  nand n75761(x75761, x68462, x75763);
  nand n75762(x75762, x75761, x72484);
  nand n75764(x75764, x68462, x75766);
  nand n75765(x75765, x75764, x72489);
  nand n75767(x75767, x68462, x75769);
  nand n75768(x75768, x75767, x72494);
  nand n75770(x75770, x68462, x75772);
  nand n75771(x75771, x75770, x72499);
  nand n75773(x75773, x68462, x75775);
  nand n75774(x75774, x75773, x72504);
  nand n75776(x75776, x68462, x75778);
  nand n75777(x75777, x75776, x72509);
  nand n75779(x75779, x68462, x75781);
  nand n75780(x75780, x75779, x72514);
  nand n75782(x75782, x68462, x75784);
  nand n75783(x75783, x75782, x72519);
  nand n75785(x75785, x68462, x75787);
  nand n75786(x75786, x75785, x72524);
  nand n75788(x75788, x68462, x75790);
  nand n75789(x75789, x75788, x72529);
  nand n75791(x75791, x68462, x75793);
  nand n75792(x75792, x75791, x72534);
  nand n75794(x75794, x68462, x75796);
  nand n75795(x75795, x75794, x72539);
  nand n75797(x75797, x68462, x75799);
  nand n75798(x75798, x75797, x72544);
  nand n75800(x75800, x68462, x75802);
  nand n75801(x75801, x75800, x72549);
  nand n75803(x75803, x68462, x75805);
  nand n75804(x75804, x75803, x72554);
  nand n75806(x75806, x68462, x75808);
  nand n75807(x75807, x75806, x72559);
  nand n75809(x75809, x68462, x75811);
  nand n75810(x75810, x75809, x72564);
  nand n75812(x75812, x68462, x75814);
  nand n75813(x75813, x75812, x72569);
  nand n75815(x75815, x68462, x75817);
  nand n75816(x75816, x75815, x72574);
  nand n75818(x75818, x68462, x75820);
  nand n75819(x75819, x75818, x72579);
  nand n75821(x75821, x68462, x75823);
  nand n75822(x75822, x75821, x72584);
  nand n75824(x75824, x68462, x75826);
  nand n75825(x75825, x75824, x72589);
  nand n75827(x75827, x68462, x75829);
  nand n75828(x75828, x75827, x72594);
  nand n75830(x75830, x68462, x75832);
  nand n75831(x75831, x75830, x72599);
  nand n75833(x75833, x68462, x75835);
  nand n75834(x75834, x75833, x72604);
  nand n75836(x75836, x68462, x75838);
  nand n75837(x75837, x75836, x72609);
  nand n75839(x75839, x68462, x75841);
  nand n75840(x75840, x75839, x72614);
  nand n75842(x75842, x68462, x75844);
  nand n75843(x75843, x75842, x72619);
  nand n75845(x75845, x68462, x75847);
  nand n75846(x75846, x75845, x72624);
  nand n75848(x75848, x68462, x75850);
  nand n75849(x75849, x75848, x72629);
  nand n75851(x75851, x68462, x75853);
  nand n75852(x75852, x75851, x72634);
  nand n75854(x75854, x68462, x75856);
  nand n75855(x75855, x75854, x72639);
  nand n75857(x75857, x68462, x75859);
  nand n75858(x75858, x75857, x72644);
  nand n75860(x75860, x68462, x75862);
  nand n75861(x75861, x75860, x72649);
  nand n75863(x75863, x68462, x75865);
  nand n75864(x75864, x75863, x72654);
  nand n75866(x75866, x68462, x75868);
  nand n75867(x75867, x75866, x72659);
  nand n75869(x75869, x68462, x75871);
  nand n75870(x75870, x75869, x72664);
  nand n75872(x75872, x68462, x75874);
  nand n75873(x75873, x75872, x72669);
  nand n75875(x75875, x68462, x75877);
  nand n75876(x75876, x75875, x72674);
  nand n75878(x75878, x68462, x75880);
  nand n75879(x75879, x75878, x72679);
  nand n75881(x75881, x68462, x75883);
  nand n75882(x75882, x75881, x72684);
  nand n75884(x75884, x68462, x75886);
  nand n75885(x75885, x75884, x72689);
  nand n75887(x75887, x68462, x75889);
  nand n75888(x75888, x75887, x72694);
  nand n75890(x75890, x68462, x75892);
  nand n75891(x75891, x75890, x72699);
  nand n75893(x75893, x68462, x75895);
  nand n75894(x75894, x75893, x72704);
  nand n75896(x75896, x68462, x75898);
  nand n75897(x75897, x75896, x72709);
  nand n75899(x75899, x68462, x75901);
  nand n75900(x75900, x75899, x72714);
  nand n75902(x75902, x68462, x75904);
  nand n75903(x75903, x75902, x72719);
  nand n75905(x75905, x68462, x75907);
  nand n75906(x75906, x75905, x72724);
  nand n75908(x75908, x68462, x75910);
  nand n75909(x75909, x75908, x72729);
  nand n75911(x75911, x68462, x75913);
  nand n75912(x75912, x75911, x72734);
  nand n75914(x75914, x68462, x75916);
  nand n75915(x75915, x75914, x72739);
  nand n75917(x75917, x68462, x75919);
  nand n75918(x75918, x75917, x72744);
  nand n75920(x75920, x68462, x75922);
  nand n75921(x75921, x75920, x72749);
  nand n75923(x75923, x68462, x75925);
  nand n75924(x75924, x75923, x72754);
  nand n75926(x75926, x68462, x75928);
  nand n75927(x75927, x75926, x72759);
  nand n75929(x75929, x68462, x75931);
  nand n75930(x75930, x75929, x72764);
  nand n75932(x75932, x68462, x75934);
  nand n75933(x75933, x75932, x72769);
  nand n75935(x75935, x68462, x75937);
  nand n75936(x75936, x75935, x72774);
  nand n75938(x75938, x68462, x75940);
  nand n75939(x75939, x75938, x72779);
  nand n75941(x75941, x68462, x75943);
  nand n75942(x75942, x75941, x72784);
  nand n75944(x75944, x68462, x75946);
  nand n75945(x75945, x75944, x72789);
  nand n75947(x75947, x68462, x75949);
  nand n75948(x75948, x75947, x72794);
  nand n75950(x75950, x68462, x75952);
  nand n75951(x75951, x75950, x72799);
  nand n75953(x75953, x68462, x75955);
  nand n75954(x75954, x75953, x72804);
  nand n75956(x75956, x68462, x75958);
  nand n75957(x75957, x75956, x72809);
  nand n75959(x75959, x68462, x75961);
  nand n75960(x75960, x75959, x72814);
  nand n75962(x75962, x68462, x75964);
  nand n75963(x75963, x75962, x72819);
  nand n75965(x75965, x68462, x75967);
  nand n75966(x75966, x75965, x72824);
  nand n75968(x75968, x68462, x75970);
  nand n75969(x75969, x75968, x72829);
  nand n75971(x75971, x68462, x75973);
  nand n75972(x75972, x75971, x72834);
  nand n75974(x75974, x68462, x75976);
  nand n75975(x75975, x75974, x72839);
  nand n75977(x75977, x68462, x75979);
  nand n75978(x75978, x75977, x72844);
  nand n75980(x75980, x68462, x75982);
  nand n75981(x75981, x75980, x72849);
  nand n75983(x75983, x68462, x75985);
  nand n75984(x75984, x75983, x72854);
  nand n75986(x75986, x68462, x75988);
  nand n75987(x75987, x75986, x72859);
  nand n75989(x75989, x68462, x75991);
  nand n75990(x75990, x75989, x72864);
  nand n75992(x75992, x68462, x75994);
  nand n75993(x75993, x75992, x72869);
  nand n75995(x75995, x68462, x75997);
  nand n75996(x75996, x75995, x72874);
  nand n75998(x75998, x68462, x76000);
  nand n75999(x75999, x75998, x72879);
  nand n76001(x76001, x68462, x76003);
  nand n76002(x76002, x76001, x72884);
  nand n76004(x76004, x68462, x76006);
  nand n76005(x76005, x76004, x72889);
  nand n76007(x76007, x68462, x76009);
  nand n76008(x76008, x76007, x72894);
  nand n76010(x76010, x68462, x76012);
  nand n76011(x76011, x76010, x72899);
  nand n76013(x76013, x68462, x76015);
  nand n76014(x76014, x76013, x72904);
  nand n76016(x76016, x68462, x76018);
  nand n76017(x76017, x76016, x72909);
  nand n76019(x76019, x68462, x76021);
  nand n76020(x76020, x76019, x72914);
  nand n76022(x76022, x68462, x76024);
  nand n76023(x76023, x76022, x72919);
  nand n76025(x76025, x68462, x76027);
  nand n76026(x76026, x76025, x72924);
  nand n76028(x76028, x68462, x76030);
  nand n76029(x76029, x76028, x72929);
  nand n76031(x76031, x68462, x76033);
  nand n76032(x76032, x76031, x72934);
  nand n76034(x76034, x68462, x76036);
  nand n76035(x76035, x76034, x72939);
  nand n76037(x76037, x68462, x76039);
  nand n76038(x76038, x76037, x72944);
  nand n76040(x76040, x68462, x76042);
  nand n76041(x76041, x76040, x72949);
  nand n76043(x76043, x68462, x76045);
  nand n76044(x76044, x76043, x72954);
  nand n76046(x76046, x68462, x76048);
  nand n76047(x76047, x76046, x72959);
  nand n76049(x76049, x68462, x76051);
  nand n76050(x76050, x76049, x72964);
  nand n76052(x76052, x68462, x76054);
  nand n76053(x76053, x76052, x72969);
  nand n76055(x76055, x68462, x76057);
  nand n76056(x76056, x76055, x72974);
  nand n76058(x76058, x68462, x76060);
  nand n76059(x76059, x76058, x72979);
  nand n76061(x76061, x68462, x76063);
  nand n76062(x76062, x76061, x72984);
  nand n76064(x76064, x68462, x76066);
  nand n76065(x76065, x76064, x72989);
  nand n76067(x76067, x68462, x76069);
  nand n76068(x76068, x76067, x72994);
  nand n76070(x76070, x68462, x76072);
  nand n76071(x76071, x76070, x72999);
  nand n76073(x76073, x68462, x76075);
  nand n76074(x76074, x76073, x73004);
  nand n76076(x76076, x68462, x76078);
  nand n76077(x76077, x76076, x73009);
  nand n76079(x76079, x68462, x76081);
  nand n76080(x76080, x76079, x73014);
  nand n76082(x76082, x68462, x76084);
  nand n76083(x76083, x76082, x73019);
  nand n76085(x76085, x68462, x76087);
  nand n76086(x76086, x76085, x73024);
  nand n76088(x76088, x68462, x76090);
  nand n76089(x76089, x76088, x73029);
  nand n76091(x76091, x68462, x76093);
  nand n76092(x76092, x76091, x73034);
  nand n76094(x76094, x68462, x76096);
  nand n76095(x76095, x76094, x73039);
  nand n76097(x76097, x68462, x76099);
  nand n76098(x76098, x76097, x73044);
  nand n76100(x76100, x68462, x76102);
  nand n76101(x76101, x76100, x73049);
  nand n76103(x76103, x68462, x76105);
  nand n76104(x76104, x76103, x73054);
  nand n76106(x76106, x68462, x76108);
  nand n76107(x76107, x76106, x73059);
  nand n76109(x76109, x68462, x76111);
  nand n76110(x76110, x76109, x73064);
  nand n76112(x76112, x68462, x76114);
  nand n76113(x76113, x76112, x73069);
  nand n76115(x76115, x68462, x76117);
  nand n76116(x76116, x76115, x73074);
  nand n76118(x76118, x68462, x76120);
  nand n76119(x76119, x76118, x73079);
  nand n76121(x76121, x68462, x76123);
  nand n76122(x76122, x76121, x73084);
  nand n76124(x76124, x68462, x76126);
  nand n76125(x76125, x76124, x73089);
  nand n76127(x76127, x68462, x76129);
  nand n76128(x76128, x76127, x73094);
  nand n76130(x76130, x68462, x76132);
  nand n76131(x76131, x76130, x73099);
  nand n76133(x76133, x68462, x76135);
  nand n76134(x76134, x76133, x73104);
  nand n76136(x76136, x68462, x76138);
  nand n76137(x76137, x76136, x73109);
  nand n76139(x76139, x68462, x76141);
  nand n76140(x76140, x76139, x73114);
  nand n76142(x76142, x68462, x76144);
  nand n76143(x76143, x76142, x73119);
  nand n76145(x76145, x68462, x76147);
  nand n76146(x76146, x76145, x73124);
  nand n76148(x76148, x68462, x76150);
  nand n76149(x76149, x76148, x73129);
  nand n76151(x76151, x68462, x76153);
  nand n76152(x76152, x76151, x73134);
  nand n76154(x76154, x68462, x76156);
  nand n76155(x76155, x76154, x73139);
  nand n76157(x76157, x68462, x76159);
  nand n76158(x76158, x76157, x73144);
  nand n76160(x76160, x68462, x76162);
  nand n76161(x76161, x76160, x73149);
  nand n76163(x76163, x68462, x76165);
  nand n76164(x76164, x76163, x73154);
  nand n76166(x76166, x68462, x76168);
  nand n76167(x76167, x76166, x73159);
  nand n76169(x76169, x68462, x76171);
  nand n76170(x76170, x76169, x73164);
  nand n76172(x76172, x68462, x76174);
  nand n76173(x76173, x76172, x73169);
  nand n76175(x76175, x68462, x76177);
  nand n76176(x76176, x76175, x73174);
  nand n76178(x76178, x68462, x76180);
  nand n76179(x76179, x76178, x73179);
  nand n76181(x76181, x68462, x76183);
  nand n76182(x76182, x76181, x73184);
  nand n76184(x76184, x68462, x76186);
  nand n76185(x76185, x76184, x73189);
  nand n76187(x76187, x68462, x76189);
  nand n76188(x76188, x76187, x73194);
  nand n76190(x76190, x68462, x76192);
  nand n76191(x76191, x76190, x73199);
  nand n76193(x76193, x68462, x76195);
  nand n76194(x76194, x76193, x73204);
  nand n76196(x76196, x68462, x76198);
  nand n76197(x76197, x76196, x73209);
  nand n76199(x76199, x68462, x76201);
  nand n76200(x76200, x76199, x73214);
  nand n76202(x76202, x68462, x76204);
  nand n76203(x76203, x76202, x73219);
  nand n76205(x76205, x68462, x76207);
  nand n76206(x76206, x76205, x73224);
  nand n76208(x76208, x68462, x76210);
  nand n76209(x76209, x76208, x73229);
  nand n76211(x76211, x68462, x76213);
  nand n76212(x76212, x76211, x73234);
  nand n76214(x76214, x68462, x76216);
  nand n76215(x76215, x76214, x73239);
  nand n76217(x76217, x68462, x76219);
  nand n76218(x76218, x76217, x73244);
  nand n76220(x76220, x68462, x76222);
  nand n76221(x76221, x76220, x73249);
  nand n76223(x76223, x68462, x76225);
  nand n76224(x76224, x76223, x73254);
  nand n76226(x76226, x68462, x76228);
  nand n76227(x76227, x76226, x73259);
  nand n76229(x76229, x68462, x76231);
  nand n76230(x76230, x76229, x73264);
  nand n76232(x76232, x68462, x76234);
  nand n76233(x76233, x76232, x73269);
  nand n76235(x76235, x68462, x76237);
  nand n76236(x76236, x76235, x73274);
  nand n76238(x76238, x68462, x76240);
  nand n76239(x76239, x76238, x73279);
  nand n76241(x76241, x68462, x76243);
  nand n76242(x76242, x76241, x73284);
  nand n76244(x76244, x68462, x76246);
  nand n76245(x76245, x76244, x73289);
  nand n76247(x76247, x68462, x76249);
  nand n76248(x76248, x76247, x73294);
  nand n76250(x76250, x68462, x76252);
  nand n76251(x76251, x76250, x73299);
  nand n76253(x76253, x68462, x76255);
  nand n76254(x76254, x76253, x73304);
  nand n76256(x76256, x68462, x76258);
  nand n76257(x76257, x76256, x73309);
  nand n76259(x76259, x68462, x76261);
  nand n76260(x76260, x76259, x73314);
  nand n76262(x76262, x68462, x76264);
  nand n76263(x76263, x76262, x73319);
  nand n76265(x76265, x68462, x76267);
  nand n76266(x76266, x76265, x73324);
  nand n76268(x76268, x68462, x76270);
  nand n76269(x76269, x76268, x73329);
  nand n76271(x76271, x68462, x76273);
  nand n76272(x76272, x76271, x73334);
  nand n76274(x76274, x68462, x76276);
  nand n76275(x76275, x76274, x73339);
  nand n76277(x76277, x68462, x76279);
  nand n76278(x76278, x76277, x73344);
  nand n76280(x76280, x68462, x76282);
  nand n76281(x76281, x76280, x73349);
  nand n76283(x76283, x68462, x76285);
  nand n76284(x76284, x76283, x73354);
  nand n76286(x76286, x68462, x76288);
  nand n76287(x76287, x76286, x73359);
  nand n76289(x76289, x68462, x76291);
  nand n76290(x76290, x76289, x73364);
  nand n76292(x76292, x68462, x76294);
  nand n76293(x76293, x76292, x73369);
  nand n76295(x76295, x68462, x76297);
  nand n76296(x76296, x76295, x73374);
  nand n76298(x76298, x68462, x76300);
  nand n76299(x76299, x76298, x73379);
  nand n76301(x76301, x68462, x76303);
  nand n76302(x76302, x76301, x73384);
  nand n76304(x76304, x68462, x76306);
  nand n76305(x76305, x76304, x73389);
  nand n76307(x76307, x68462, x76309);
  nand n76308(x76308, x76307, x73394);
  nand n76310(x76310, x68462, x76312);
  nand n76311(x76311, x76310, x73399);
  nand n76313(x76313, x68462, x76315);
  nand n76314(x76314, x76313, x73404);
  nand n76316(x76316, x68462, x76318);
  nand n76317(x76317, x76316, x73409);
  nand n76319(x76319, x68462, x76321);
  nand n76320(x76320, x76319, x73414);
  nand n76322(x76322, x68462, x76324);
  nand n76323(x76323, x76322, x73419);
  nand n76325(x76325, x68462, x76327);
  nand n76326(x76326, x76325, x73424);
  nand n76328(x76328, x68462, x76330);
  nand n76329(x76329, x76328, x73429);
  nand n76331(x76331, x68462, x76333);
  nand n76332(x76332, x76331, x73434);
  nand n76334(x76334, x68462, x76336);
  nand n76335(x76335, x76334, x73439);
  nand n76337(x76337, x68462, x76339);
  nand n76338(x76338, x76337, x73444);
  nand n76340(x76340, x68462, x76342);
  nand n76341(x76341, x76340, x73449);
  nand n76343(x76343, x68462, x76345);
  nand n76344(x76344, x76343, x73454);
  nand n76346(x76346, x68462, x76348);
  nand n76347(x76347, x76346, x73459);
  nand n76349(x76349, x68462, x76351);
  nand n76350(x76350, x76349, x73464);
  nand n76352(x76352, x68462, x76354);
  nand n76353(x76353, x76352, x73469);
  nand n76355(x76355, x68462, x76357);
  nand n76356(x76356, x76355, x73474);
  nand n76358(x76358, x68462, x76360);
  nand n76359(x76359, x76358, x73479);
  nand n76361(x76361, x68462, x76363);
  nand n76362(x76362, x76361, x73484);
  nand n76364(x76364, x68462, x76366);
  nand n76365(x76365, x76364, x73489);
  nand n76367(x76367, x68462, x76369);
  nand n76368(x76368, x76367, x73494);
  nand n76370(x76370, x68462, x76372);
  nand n76371(x76371, x76370, x73499);
  nand n76373(x76373, x68462, x76375);
  nand n76374(x76374, x76373, x73504);
  nand n76376(x76376, x68462, x76378);
  nand n76377(x76377, x76376, x73509);
  nand n76379(x76379, x68462, x76381);
  nand n76380(x76380, x76379, x73514);
  nand n76382(x76382, x68462, x76384);
  nand n76383(x76383, x76382, x73519);
  nand n76385(x76385, x68462, x76387);
  nand n76386(x76386, x76385, x73524);
  nand n76388(x76388, x68462, x76390);
  nand n76389(x76389, x76388, x73529);
  nand n76391(x76391, x68462, x76393);
  nand n76392(x76392, x76391, x73534);
  nand n76394(x76394, x68462, x76396);
  nand n76395(x76395, x76394, x73539);
  nand n76397(x76397, x68462, x76399);
  nand n76398(x76398, x76397, x73544);
  nand n76400(x76400, x68462, x76402);
  nand n76401(x76401, x76400, x73549);
  nand n76403(x76403, x68462, x76405);
  nand n76404(x76404, x76403, x73554);
  nand n76406(x76406, x68462, x76408);
  nand n76407(x76407, x76406, x73559);
  nand n76409(x76409, x68462, x76411);
  nand n76410(x76410, x76409, x73564);
  nand n76412(x76412, x68462, x76414);
  nand n76413(x76413, x76412, x73569);
  nand n76415(x76415, x68462, x76417);
  nand n76416(x76416, x76415, x73574);
  nand n76418(x76418, x68462, x76420);
  nand n76419(x76419, x76418, x73579);
  nand n76421(x76421, x68462, x76423);
  nand n76422(x76422, x76421, x73584);
  nand n76424(x76424, x68462, x76426);
  nand n76425(x76425, x76424, x73589);
  nand n76427(x76427, x68462, x76429);
  nand n76428(x76428, x76427, x73594);
  nand n76430(x76430, x68462, x76432);
  nand n76431(x76431, x76430, x73599);
  nand n76433(x76433, x68462, x76435);
  nand n76434(x76434, x76433, x73604);
  nand n76436(x76436, x68462, x76438);
  nand n76437(x76437, x76436, x73609);
  nand n76439(x76439, x68462, x76441);
  nand n76440(x76440, x76439, x73614);
  nand n76442(x76442, x68462, x76444);
  nand n76443(x76443, x76442, x73619);
  nand n76445(x76445, x68462, x76447);
  nand n76446(x76446, x76445, x73624);
  nand n76448(x76448, x68462, x76450);
  nand n76449(x76449, x76448, x73629);
  nand n76451(x76451, x68462, x76453);
  nand n76452(x76452, x76451, x73634);
  nand n76454(x76454, x68462, x76456);
  nand n76455(x76455, x76454, x73639);
  nand n76457(x76457, x68462, x76459);
  nand n76458(x76458, x76457, x73644);
  nand n76460(x76460, x68462, x76462);
  nand n76461(x76461, x76460, x73649);
  nand n76463(x76463, x68462, x76465);
  nand n76464(x76464, x76463, x73654);
  nand n76466(x76466, x68462, x76468);
  nand n76467(x76467, x76466, x73659);
  nand n76469(x76469, x68462, x76471);
  nand n76470(x76470, x76469, x73664);
  nand n76472(x76472, x68462, x76474);
  nand n76473(x76473, x76472, x73669);
  nand n76475(x76475, x68462, x76477);
  nand n76476(x76476, x76475, x73674);
  nand n76478(x76478, x68462, x76480);
  nand n76479(x76479, x76478, x73679);
  nand n76481(x76481, x68462, x76483);
  nand n76482(x76482, x76481, x73684);
  nand n76484(x76484, x68462, x76486);
  nand n76485(x76485, x76484, x73689);
  nand n76487(x76487, x68462, x76489);
  nand n76488(x76488, x76487, x73694);
  nand n76490(x76490, x68462, x76492);
  nand n76491(x76491, x76490, x73699);
  nand n76493(x76493, x68462, x76495);
  nand n76494(x76494, x76493, x73704);
  nand n76496(x76496, x68462, x76498);
  nand n76497(x76497, x76496, x73709);
  nand n76499(x76499, x68462, x76501);
  nand n76500(x76500, x76499, x73714);
  nand n76502(x76502, x68462, x76504);
  nand n76503(x76503, x76502, x73719);
  nand n76505(x76505, x68462, x76507);
  nand n76506(x76506, x76505, x73724);
  nand n76508(x76508, x68462, x76510);
  nand n76509(x76509, x76508, x73729);
  nand n76511(x76511, x68462, x76513);
  nand n76512(x76512, x76511, x73734);
  nand n76514(x76514, x68462, x76516);
  nand n76515(x76515, x76514, x73739);
  nand n76517(x76517, x68462, x76519);
  nand n76518(x76518, x76517, x73744);
  nand n76520(x76520, x68462, x76522);
  nand n76521(x76521, x76520, x73749);
  nand n76523(x76523, x68462, x76525);
  nand n76524(x76524, x76523, x73754);
  nand n76526(x76526, x68462, x76528);
  nand n76527(x76527, x76526, x73759);
  nand n76529(x76529, x68462, x76531);
  nand n76530(x76530, x76529, x73764);
  nand n76532(x76532, x68462, x76534);
  nand n76533(x76533, x76532, x73769);
  nand n76535(x76535, x68462, x76537);
  nand n76536(x76536, x76535, x73774);
  nand n76538(x76538, x68462, x76540);
  nand n76539(x76539, x76538, x73779);
  nand n76541(x76541, x68462, x76543);
  nand n76542(x76542, x76541, x73784);
  nand n76544(x76544, x68462, x76546);
  nand n76545(x76545, x76544, x73789);
  nand n76547(x76547, x68462, x76549);
  nand n76548(x76548, x76547, x73794);
  nand n76550(x76550, x68462, x76552);
  nand n76551(x76551, x76550, x73799);
  nand n76553(x76553, x68462, x76555);
  nand n76554(x76554, x76553, x73804);
  nand n76556(x76556, x68462, x76558);
  nand n76557(x76557, x76556, x73809);
  nand n76559(x76559, x68462, x76561);
  nand n76560(x76560, x76559, x73814);
  nand n76562(x76562, x68462, x76564);
  nand n76563(x76563, x76562, x73819);
  nand n76565(x76565, x68462, x76567);
  nand n76566(x76566, x76565, x73824);
  nand n76568(x76568, x68462, x76570);
  nand n76569(x76569, x76568, x73829);
  nand n76571(x76571, x68462, x76573);
  nand n76572(x76572, x76571, x73834);
  nand n76574(x76574, x68462, x76576);
  nand n76575(x76575, x76574, x73839);
  nand n76577(x76577, x68462, x76579);
  nand n76578(x76578, x76577, x73844);
  nand n76580(x76580, x68462, x76582);
  nand n76581(x76581, x76580, x73849);
  nand n76583(x76583, x68462, x76585);
  nand n76584(x76584, x76583, x73854);
  nand n76586(x76586, x68462, x76588);
  nand n76587(x76587, x76586, x73859);
  nand n76589(x76589, x68462, x76591);
  nand n76590(x76590, x76589, x73864);
  nand n76592(x76592, x68462, x76594);
  nand n76593(x76593, x76592, x73869);
  nand n76595(x76595, x68462, x76597);
  nand n76596(x76596, x76595, x73874);
  nand n76598(x76598, x68462, x76600);
  nand n76599(x76599, x76598, x73879);
  nand n76601(x76601, x68462, x76603);
  nand n76602(x76602, x76601, x73884);
  nand n76604(x76604, x68462, x76606);
  nand n76605(x76605, x76604, x73889);
  nand n76607(x76607, x68462, x76609);
  nand n76608(x76608, x76607, x73894);
  nand n76610(x76610, x68462, x76612);
  nand n76611(x76611, x76610, x73899);
  nand n76613(x76613, x68462, x76615);
  nand n76614(x76614, x76613, x73904);
  nand n76616(x76616, x68462, x76618);
  nand n76617(x76617, x76616, x73909);
  nand n76619(x76619, x68462, x76621);
  nand n76620(x76620, x76619, x73914);
  nand n76622(x76622, x68462, x76624);
  nand n76623(x76623, x76622, x73919);
  nand n76625(x76625, x68462, x76627);
  nand n76626(x76626, x76625, x73924);
  nand n76628(x76628, x68462, x76630);
  nand n76629(x76629, x76628, x73929);
  nand n76631(x76631, x68462, x76633);
  nand n76632(x76632, x76631, x73934);
  nand n76634(x76634, x68462, x76636);
  nand n76635(x76635, x76634, x73939);
  nand n76637(x76637, x68462, x76639);
  nand n76638(x76638, x76637, x73944);
  nand n76640(x76640, x68462, x76642);
  nand n76641(x76641, x76640, x73949);
  nand n76643(x76643, x68462, x76645);
  nand n76644(x76644, x76643, x73954);
  nand n76646(x76646, x68462, x76648);
  nand n76647(x76647, x76646, x73959);
  nand n76649(x76649, x68462, x76651);
  nand n76650(x76650, x76649, x73964);
  nand n76652(x76652, x68462, x76654);
  nand n76653(x76653, x76652, x73969);
  nand n76655(x76655, x68462, x76657);
  nand n76656(x76656, x76655, x73974);
  nand n76658(x76658, x68462, x76660);
  nand n76659(x76659, x76658, x73979);
  nand n76661(x76661, x68462, x76663);
  nand n76662(x76662, x76661, x73984);
  nand n76664(x76664, x68462, x76666);
  nand n76665(x76665, x76664, x73989);
  nand n76667(x76667, x68462, x76669);
  nand n76668(x76668, x76667, x73994);
  nand n76670(x76670, x68462, x76672);
  nand n76671(x76671, x76670, x73999);
  nand n76673(x76673, x68462, x76675);
  nand n76674(x76674, x76673, x71799);
  nand n76676(x76676, x68462, x76678);
  nand n76677(x76677, x76676, x71804);
  nand n76679(x76679, x68462, x76681);
  nand n76680(x76680, x76679, x71809);
  nand n76682(x76682, x68462, x76684);
  nand n76683(x76683, x76682, x71814);
  nand n76685(x76685, x68462, x76687);
  nand n76686(x76686, x76685, x71819);
  nand n76688(x76688, x68462, x76690);
  nand n76689(x76689, x76688, x71824);
  nand n76691(x76691, x68462, x76693);
  nand n76692(x76692, x76691, x71829);
  nand n76694(x76694, x68462, x76696);
  nand n76695(x76695, x76694, x71834);
  nand n76697(x76697, x68462, x76699);
  nand n76698(x76698, x76697, x71839);
  nand n76700(x76700, x68462, x76702);
  nand n76701(x76701, x76700, x71844);
  nand n76703(x76703, x68462, x76705);
  nand n76704(x76704, x76703, x71849);
  nand n76706(x76706, x68462, x76708);
  nand n76707(x76707, x76706, x71854);
  nand n76709(x76709, x68462, x76711);
  nand n76710(x76710, x76709, x71859);
  nand n76712(x76712, x68462, x76714);
  nand n76713(x76713, x76712, x71864);
  nand n76715(x76715, x68462, x76717);
  nand n76716(x76716, x76715, x71869);
  nand n76718(x76718, x68462, x76720);
  nand n76719(x76719, x76718, x71874);
  nand n76721(x76721, x68462, x76723);
  nand n76722(x76722, x76721, x71879);
  nand n76724(x76724, x68462, x76726);
  nand n76725(x76725, x76724, x71884);
  nand n76727(x76727, x68462, x76729);
  nand n76728(x76728, x76727, x71889);
  nand n76730(x76730, x68462, x76732);
  nand n76731(x76731, x76730, x71894);
  nand n76733(x76733, x68462, x76735);
  nand n76734(x76734, x76733, x71899);
  nand n76736(x76736, x68462, x76738);
  nand n76737(x76737, x76736, x71904);
  nand n76739(x76739, x68462, x76741);
  nand n76740(x76740, x76739, x71904);
  nand n76742(x76742, x68462, x76744);
  nand n76743(x76743, x76742, x71904);
  nand n76745(x76745, x68462, x76747);
  nand n76746(x76746, x76745, x71904);
  nand n76748(x76748, x68462, x76750);
  nand n76749(x76749, x76748, x71904);
  nand n76751(x76751, x68462, x76753);
  nand n76752(x76752, x76751, x71904);
  nand n76754(x76754, x68462, x76756);
  nand n76755(x76755, x76754, x71904);
  nand n76757(x76757, x68462, x76759);
  nand n76758(x76758, x76757, x71904);
  nand n76760(x76760, x68462, x76762);
  nand n76761(x76761, x76760, x71904);
  nand n76763(x76763, x68462, x76765);
  nand n76764(x76764, x76763, x71904);
  nand n76766(x76766, x68462, x76768);
  nand n76767(x76767, x76766, x71904);
  nand n76769(x76769, x68462, x76771);
  nand n76770(x76770, x76769, x71939);
  nand n76772(x76772, x68462, x76774);
  nand n76773(x76773, x76772, x71944);
  nand n76775(x76775, x68462, x76777);
  nand n76776(x76776, x76775, x71949);
  nand n76778(x76778, x68462, x76780);
  nand n76779(x76779, x76778, x71954);
  nand n76781(x76781, x68462, x76783);
  nand n76782(x76782, x76781, x71959);
  nand n76784(x76784, x68462, x76786);
  nand n76785(x76785, x76784, x71964);
  nand n76787(x76787, x68462, x76789);
  nand n76788(x76788, x76787, x71969);
  nand n76790(x76790, x68462, x76792);
  nand n76791(x76791, x76790, x71974);
  nand n76793(x76793, x68462, x76795);
  nand n76794(x76794, x76793, x71979);
  nand n76796(x76796, x68462, x76798);
  nand n76797(x76797, x76796, x71984);
  nand n76799(x76799, x68462, x76801);
  nand n76800(x76800, x76799, x71989);
  nand n76802(x76802, x68462, x76804);
  nand n76803(x76803, x76802, x71994);
  nand n76805(x76805, x68462, x76807);
  nand n76806(x76806, x76805, x71999);
  nand n76808(x76808, x68462, x76810);
  nand n76809(x76809, x76808, x72004);
  nand n76811(x76811, x68462, x76813);
  nand n76812(x76812, x76811, x72009);
  nand n76814(x76814, x68462, x76816);
  nand n76815(x76815, x76814, x72014);
  nand n76817(x76817, x68462, x76819);
  nand n76818(x76818, x76817, x72019);
  nand n76820(x76820, x68462, x76822);
  nand n76821(x76821, x76820, x72024);
  nand n76823(x76823, x68462, x76825);
  nand n76824(x76824, x76823, x72029);
  nand n76826(x76826, x68462, x76828);
  nand n76827(x76827, x76826, x72034);
  nand n76829(x76829, x68462, x76831);
  nand n76830(x76830, x76829, x72039);
  nand n76832(x76832, x68462, x76834);
  nand n76833(x76833, x76832, x72044);
  nand n76835(x76835, x68462, x76837);
  nand n76836(x76836, x76835, x72049);
  nand n76838(x76838, x68462, x76840);
  nand n76839(x76839, x76838, x72054);
  nand n76841(x76841, x68462, x76843);
  nand n76842(x76842, x76841, x72059);
  nand n76844(x76844, x68462, x76846);
  nand n76845(x76845, x76844, x72064);
  nand n76847(x76847, x68462, x76849);
  nand n76848(x76848, x76847, x72069);
  nand n76850(x76850, x68462, x76852);
  nand n76851(x76851, x76850, x72074);
  nand n76853(x76853, x68462, x76855);
  nand n76854(x76854, x76853, x72079);
  nand n76856(x76856, x68462, x76858);
  nand n76857(x76857, x76856, x72084);
  nand n76859(x76859, x68462, x76861);
  nand n76860(x76860, x76859, x72089);
  nand n76862(x76862, x68462, x76864);
  nand n76863(x76863, x76862, x72094);
  nand n76865(x76865, x68462, x76867);
  nand n76866(x76866, x76865, x72099);
  nand n76868(x76868, x68462, x76870);
  nand n76869(x76869, x76868, x72104);
  nand n76871(x76871, x68462, x76873);
  nand n76872(x76872, x76871, x72109);
  nand n76874(x76874, x68462, x76876);
  nand n76875(x76875, x76874, x72114);
  nand n76877(x76877, x68462, x76879);
  nand n76878(x76878, x76877, x72119);
  nand n76880(x76880, x68462, x76882);
  nand n76881(x76881, x76880, x72124);
  nand n76883(x76883, x68462, x76885);
  nand n76884(x76884, x76883, x72129);
  nand n76886(x76886, x68462, x76888);
  nand n76887(x76887, x76886, x72134);
  nand n76889(x76889, x68462, x76891);
  nand n76890(x76890, x76889, x72139);
  nand n76892(x76892, x68462, x76894);
  nand n76893(x76893, x76892, x72144);
  nand n76895(x76895, x68462, x76897);
  nand n76896(x76896, x76895, x72149);
  nand n76898(x76898, x68462, x76900);
  nand n76899(x76899, x76898, x72154);
  nand n76901(x76901, x68462, x76903);
  nand n76902(x76902, x76901, x72159);
  nand n76904(x76904, x68462, x76906);
  nand n76905(x76905, x76904, x72164);
  nand n76907(x76907, x68462, x76909);
  nand n76908(x76908, x76907, x72169);
  nand n76910(x76910, x68462, x76912);
  nand n76911(x76911, x76910, x72174);
  nand n76913(x76913, x68462, x76915);
  nand n76914(x76914, x76913, x72179);
  nand n76916(x76916, x68462, x76918);
  nand n76917(x76917, x76916, x72184);
  nand n76919(x76919, x68462, x76921);
  nand n76920(x76920, x76919, x72189);
  nand n76922(x76922, x68462, x76924);
  nand n76923(x76923, x76922, x72194);
  nand n76925(x76925, x68462, x76927);
  nand n76926(x76926, x76925, x72199);
  nand n76928(x76928, x68462, x76930);
  nand n76929(x76929, x76928, x72204);
  nand n76931(x76931, x68462, x76933);
  nand n76932(x76932, x76931, x72209);
  nand n76934(x76934, x68462, x76936);
  nand n76935(x76935, x76934, x72214);
  nand n76937(x76937, x68462, x76939);
  nand n76938(x76938, x76937, x72219);
  nand n76940(x76940, x68462, x76942);
  nand n76941(x76941, x76940, x72224);
  nand n76943(x76943, x68462, x76945);
  nand n76944(x76944, x76943, x72229);
  nand n76946(x76946, x68462, x76948);
  nand n76947(x76947, x76946, x72234);
  nand n76949(x76949, x68462, x76951);
  nand n76950(x76950, x76949, x72239);
  nand n76952(x76952, x68462, x76954);
  nand n76953(x76953, x76952, x72244);
  nand n76955(x76955, x68462, x76957);
  nand n76956(x76956, x76955, x72249);
  nand n76958(x76958, x68462, x76960);
  nand n76959(x76959, x76958, x72254);
  nand n76961(x76961, x68462, x76963);
  nand n76962(x76962, x76961, x72259);
  nand n76964(x76964, x68462, x76966);
  nand n76965(x76965, x76964, x72264);
  nand n76967(x76967, x68462, x76969);
  nand n76968(x76968, x76967, x72269);
  nand n76970(x76970, x68462, x76972);
  nand n76971(x76971, x76970, x72274);
  nand n76973(x76973, x68462, x76975);
  nand n76974(x76974, x76973, x72279);
  nand n76976(x76976, x68462, x76978);
  nand n76977(x76977, x76976, x72284);
  nand n76979(x76979, x68462, x76981);
  nand n76980(x76980, x76979, x72289);
  nand n76982(x76982, x68462, x76984);
  nand n76983(x76983, x76982, x72294);
  nand n76985(x76985, x68462, x76987);
  nand n76986(x76986, x76985, x72299);
  nand n76988(x76988, x68462, x76990);
  nand n76989(x76989, x76988, x72304);
  nand n76991(x76991, x68462, x76993);
  nand n76992(x76992, x76991, x72309);
  nand n76994(x76994, x68462, x76996);
  nand n76995(x76995, x76994, x72314);
  nand n76997(x76997, x68462, x76999);
  nand n76998(x76998, x76997, x72319);
  nand n77000(x77000, x68462, x77002);
  nand n77001(x77001, x77000, x72324);
  nand n77003(x77003, x68462, x77005);
  nand n77004(x77004, x77003, x72329);
  nand n77006(x77006, x68462, x77008);
  nand n77007(x77007, x77006, x72334);
  nand n77009(x77009, x68462, x77011);
  nand n77010(x77010, x77009, x72339);
  nand n77012(x77012, x68462, x77014);
  nand n77013(x77013, x77012, x72344);
  nand n77015(x77015, x68462, x77017);
  nand n77016(x77016, x77015, x72349);
  nand n77018(x77018, x68462, x77020);
  nand n77019(x77019, x77018, x72354);
  nand n77021(x77021, x68462, x77023);
  nand n77022(x77022, x77021, x72359);
  nand n77024(x77024, x68462, x77026);
  nand n77025(x77025, x77024, x72364);
  nand n77027(x77027, x68462, x77029);
  nand n77028(x77028, x77027, x72369);
  nand n77030(x77030, x68462, x77032);
  nand n77031(x77031, x77030, x72374);
  nand n77033(x77033, x68462, x77035);
  nand n77034(x77034, x77033, x72379);
  nand n77036(x77036, x68462, x77038);
  nand n77037(x77037, x77036, x72384);
  nand n77039(x77039, x68462, x77041);
  nand n77040(x77040, x77039, x72389);
  nand n77042(x77042, x68462, x77044);
  nand n77043(x77043, x77042, x72394);
  nand n77045(x77045, x68462, x77047);
  nand n77046(x77046, x77045, x72399);
  nand n77048(x77048, x68462, x77050);
  nand n77049(x77049, x77048, x72404);
  nand n77051(x77051, x68462, x77053);
  nand n77052(x77052, x77051, x72409);
  nand n77054(x77054, x68462, x77056);
  nand n77055(x77055, x77054, x72414);
  nand n77057(x77057, x68462, x77059);
  nand n77058(x77058, x77057, x72419);
  nand n77060(x77060, x68462, x77062);
  nand n77061(x77061, x77060, x72424);
  nand n77063(x77063, x68462, x77065);
  nand n77064(x77064, x77063, x72429);
  nand n77066(x77066, x68462, x77068);
  nand n77067(x77067, x77066, x72434);
  nand n77069(x77069, x68462, x77071);
  nand n77070(x77070, x77069, x72439);
  nand n77072(x77072, x68462, x77074);
  nand n77073(x77073, x77072, x72444);
  nand n77075(x77075, x68462, x77077);
  nand n77076(x77076, x77075, x72449);
  nand n77078(x77078, x68462, x77080);
  nand n77079(x77079, x77078, x72454);
  nand n77081(x77081, x68462, x77083);
  nand n77082(x77082, x77081, x72459);
  nand n77084(x77084, x68462, x77086);
  nand n77085(x77085, x77084, x72464);
  nand n77087(x77087, x68462, x77089);
  nand n77088(x77088, x77087, x72469);
  nand n77090(x77090, x68462, x77092);
  nand n77091(x77091, x77090, x72474);
  nand n77093(x77093, x68462, x77095);
  nand n77094(x77094, x77093, x72479);
  nand n77096(x77096, x68462, x77098);
  nand n77097(x77097, x77096, x72484);
  nand n77099(x77099, x68462, x77101);
  nand n77100(x77100, x77099, x72489);
  nand n77102(x77102, x68462, x77104);
  nand n77103(x77103, x77102, x72494);
  nand n77105(x77105, x68462, x77107);
  nand n77106(x77106, x77105, x72499);
  nand n77108(x77108, x68462, x77110);
  nand n77109(x77109, x77108, x72504);
  nand n77111(x77111, x68462, x77113);
  nand n77112(x77112, x77111, x72509);
  nand n77114(x77114, x68462, x77116);
  nand n77115(x77115, x77114, x72514);
  nand n77117(x77117, x68462, x77119);
  nand n77118(x77118, x77117, x72519);
  nand n77120(x77120, x68462, x77122);
  nand n77121(x77121, x77120, x72524);
  nand n77123(x77123, x68462, x77125);
  nand n77124(x77124, x77123, x72529);
  nand n77126(x77126, x68462, x77128);
  nand n77127(x77127, x77126, x72534);
  nand n77129(x77129, x68462, x77131);
  nand n77130(x77130, x77129, x72539);
  nand n77132(x77132, x68462, x77134);
  nand n77133(x77133, x77132, x72544);
  nand n77135(x77135, x68462, x77137);
  nand n77136(x77136, x77135, x72549);
  nand n77138(x77138, x68462, x77140);
  nand n77139(x77139, x77138, x72554);
  nand n77141(x77141, x68462, x77143);
  nand n77142(x77142, x77141, x72559);
  nand n77144(x77144, x68462, x77146);
  nand n77145(x77145, x77144, x72564);
  nand n77147(x77147, x68462, x77149);
  nand n77148(x77148, x77147, x72569);
  nand n77150(x77150, x68462, x77152);
  nand n77151(x77151, x77150, x72574);
  nand n77153(x77153, x68462, x77155);
  nand n77154(x77154, x77153, x72579);
  nand n77156(x77156, x68462, x77158);
  nand n77157(x77157, x77156, x72584);
  nand n77159(x77159, x68462, x77161);
  nand n77160(x77160, x77159, x72589);
  nand n77162(x77162, x68462, x77164);
  nand n77163(x77163, x77162, x72594);
  nand n77165(x77165, x68462, x77167);
  nand n77166(x77166, x77165, x72599);
  nand n77168(x77168, x68462, x77170);
  nand n77169(x77169, x77168, x72604);
  nand n77171(x77171, x68462, x77173);
  nand n77172(x77172, x77171, x72609);
  nand n77174(x77174, x68462, x77176);
  nand n77175(x77175, x77174, x72614);
  nand n77177(x77177, x68462, x77179);
  nand n77178(x77178, x77177, x72619);
  nand n77180(x77180, x68462, x77182);
  nand n77181(x77181, x77180, x72624);
  nand n77183(x77183, x68462, x77185);
  nand n77184(x77184, x77183, x72629);
  nand n77186(x77186, x68462, x77188);
  nand n77187(x77187, x77186, x72634);
  nand n77189(x77189, x68462, x77191);
  nand n77190(x77190, x77189, x72639);
  nand n77192(x77192, x68462, x77194);
  nand n77193(x77193, x77192, x72644);
  nand n77195(x77195, x68462, x77197);
  nand n77196(x77196, x77195, x72649);
  nand n77198(x77198, x68462, x77200);
  nand n77199(x77199, x77198, x72654);
  nand n77201(x77201, x68462, x77203);
  nand n77202(x77202, x77201, x72659);
  nand n77204(x77204, x68462, x77206);
  nand n77205(x77205, x77204, x72664);
  nand n77207(x77207, x68462, x77209);
  nand n77208(x77208, x77207, x72669);
  nand n77210(x77210, x68462, x77212);
  nand n77211(x77211, x77210, x72674);
  nand n77213(x77213, x68462, x77215);
  nand n77214(x77214, x77213, x72679);
  nand n77216(x77216, x68462, x77218);
  nand n77217(x77217, x77216, x72684);
  nand n77219(x77219, x68462, x77221);
  nand n77220(x77220, x77219, x72689);
  nand n77222(x77222, x68462, x77224);
  nand n77223(x77223, x77222, x72694);
  nand n77225(x77225, x68462, x77227);
  nand n77226(x77226, x77225, x72699);
  nand n77228(x77228, x68462, x77230);
  nand n77229(x77229, x77228, x72704);
  nand n77231(x77231, x68462, x77233);
  nand n77232(x77232, x77231, x72709);
  nand n77234(x77234, x68462, x77236);
  nand n77235(x77235, x77234, x72714);
  nand n77237(x77237, x68462, x77239);
  nand n77238(x77238, x77237, x72719);
  nand n77240(x77240, x68462, x77242);
  nand n77241(x77241, x77240, x72724);
  nand n77243(x77243, x68462, x77245);
  nand n77244(x77244, x77243, x72729);
  nand n77246(x77246, x68462, x77248);
  nand n77247(x77247, x77246, x72734);
  nand n77249(x77249, x68462, x77251);
  nand n77250(x77250, x77249, x72739);
  nand n77252(x77252, x68462, x77254);
  nand n77253(x77253, x77252, x72744);
  nand n77255(x77255, x68462, x77257);
  nand n77256(x77256, x77255, x72749);
  nand n77258(x77258, x68462, x77260);
  nand n77259(x77259, x77258, x72754);
  nand n77261(x77261, x68462, x77263);
  nand n77262(x77262, x77261, x72759);
  nand n77264(x77264, x68462, x77266);
  nand n77265(x77265, x77264, x72764);
  nand n77267(x77267, x68462, x77269);
  nand n77268(x77268, x77267, x72769);
  nand n77270(x77270, x68462, x77272);
  nand n77271(x77271, x77270, x72774);
  nand n77273(x77273, x68462, x77275);
  nand n77274(x77274, x77273, x72779);
  nand n77276(x77276, x68462, x77278);
  nand n77277(x77277, x77276, x72784);
  nand n77279(x77279, x68462, x77281);
  nand n77280(x77280, x77279, x72789);
  nand n77282(x77282, x68462, x77284);
  nand n77283(x77283, x77282, x72794);
  nand n77285(x77285, x68462, x77287);
  nand n77286(x77286, x77285, x72799);
  nand n77288(x77288, x68462, x77290);
  nand n77289(x77289, x77288, x72804);
  nand n77291(x77291, x68462, x77293);
  nand n77292(x77292, x77291, x72809);
  nand n77294(x77294, x68462, x77296);
  nand n77295(x77295, x77294, x72814);
  nand n77297(x77297, x68462, x77299);
  nand n77298(x77298, x77297, x72819);
  nand n77300(x77300, x68462, x77302);
  nand n77301(x77301, x77300, x72824);
  nand n77303(x77303, x68462, x77305);
  nand n77304(x77304, x77303, x72829);
  nand n77306(x77306, x68462, x77308);
  nand n77307(x77307, x77306, x72834);
  nand n77309(x77309, x68462, x77311);
  nand n77310(x77310, x77309, x72839);
  nand n77312(x77312, x68462, x77314);
  nand n77313(x77313, x77312, x72844);
  nand n77315(x77315, x68462, x77317);
  nand n77316(x77316, x77315, x72849);
  nand n77318(x77318, x68462, x77320);
  nand n77319(x77319, x77318, x72854);
  nand n77321(x77321, x68462, x77323);
  nand n77322(x77322, x77321, x72859);
  nand n77324(x77324, x68462, x77326);
  nand n77325(x77325, x77324, x72864);
  nand n77327(x77327, x68462, x77329);
  nand n77328(x77328, x77327, x72869);
  nand n77330(x77330, x68462, x77332);
  nand n77331(x77331, x77330, x72874);
  nand n77333(x77333, x68462, x77335);
  nand n77334(x77334, x77333, x72879);
  nand n77336(x77336, x68462, x77338);
  nand n77337(x77337, x77336, x72884);
  nand n77339(x77339, x68462, x77341);
  nand n77340(x77340, x77339, x72889);
  nand n77342(x77342, x68462, x77344);
  nand n77343(x77343, x77342, x72894);
  nand n77345(x77345, x68462, x77347);
  nand n77346(x77346, x77345, x72899);
  nand n77348(x77348, x68462, x77350);
  nand n77349(x77349, x77348, x72904);
  nand n77351(x77351, x68462, x77353);
  nand n77352(x77352, x77351, x72909);
  nand n77354(x77354, x68462, x77356);
  nand n77355(x77355, x77354, x72914);
  nand n77357(x77357, x68462, x77359);
  nand n77358(x77358, x77357, x72919);
  nand n77360(x77360, x68462, x77362);
  nand n77361(x77361, x77360, x72924);
  nand n77363(x77363, x68462, x77365);
  nand n77364(x77364, x77363, x72929);
  nand n77366(x77366, x68462, x77368);
  nand n77367(x77367, x77366, x72934);
  nand n77369(x77369, x68462, x77371);
  nand n77370(x77370, x77369, x72939);
  nand n77372(x77372, x68462, x77374);
  nand n77373(x77373, x77372, x72944);
  nand n77375(x77375, x68462, x77377);
  nand n77376(x77376, x77375, x72949);
  nand n77378(x77378, x68462, x77380);
  nand n77379(x77379, x77378, x72954);
  nand n77381(x77381, x68462, x77383);
  nand n77382(x77382, x77381, x72959);
  nand n77384(x77384, x68462, x77386);
  nand n77385(x77385, x77384, x72964);
  nand n77387(x77387, x68462, x77389);
  nand n77388(x77388, x77387, x72969);
  nand n77390(x77390, x68462, x77392);
  nand n77391(x77391, x77390, x72974);
  nand n77393(x77393, x68462, x77395);
  nand n77394(x77394, x77393, x72979);
  nand n77396(x77396, x68462, x77398);
  nand n77397(x77397, x77396, x72984);
  nand n77399(x77399, x68462, x77401);
  nand n77400(x77400, x77399, x72989);
  nand n77402(x77402, x68462, x77404);
  nand n77403(x77403, x77402, x72994);
  nand n77405(x77405, x68462, x77407);
  nand n77406(x77406, x77405, x72999);
  nand n77408(x77408, x68462, x77410);
  nand n77409(x77409, x77408, x73004);
  nand n77411(x77411, x68462, x77413);
  nand n77412(x77412, x77411, x73009);
  nand n77414(x77414, x68462, x77416);
  nand n77415(x77415, x77414, x73014);
  nand n77417(x77417, x68462, x77419);
  nand n77418(x77418, x77417, x73019);
  nand n77420(x77420, x68462, x77422);
  nand n77421(x77421, x77420, x73024);
  nand n77423(x77423, x68462, x77425);
  nand n77424(x77424, x77423, x73029);
  nand n77426(x77426, x68462, x77428);
  nand n77427(x77427, x77426, x73034);
  nand n77429(x77429, x68462, x77431);
  nand n77430(x77430, x77429, x73039);
  nand n77432(x77432, x68462, x77434);
  nand n77433(x77433, x77432, x73044);
  nand n77435(x77435, x68462, x77437);
  nand n77436(x77436, x77435, x73049);
  nand n77438(x77438, x68462, x77440);
  nand n77439(x77439, x77438, x73054);
  nand n77441(x77441, x68462, x77443);
  nand n77442(x77442, x77441, x73059);
  nand n77444(x77444, x68462, x77446);
  nand n77445(x77445, x77444, x73064);
  nand n77447(x77447, x68462, x77449);
  nand n77448(x77448, x77447, x73069);
  nand n77450(x77450, x68462, x77452);
  nand n77451(x77451, x77450, x73074);
  nand n77453(x77453, x68462, x77455);
  nand n77454(x77454, x77453, x73079);
  nand n77456(x77456, x68462, x77458);
  nand n77457(x77457, x77456, x73084);
  nand n77459(x77459, x68462, x77461);
  nand n77460(x77460, x77459, x73089);
  nand n77462(x77462, x68462, x77464);
  nand n77463(x77463, x77462, x73094);
  nand n77465(x77465, x68462, x77467);
  nand n77466(x77466, x77465, x73099);
  nand n77468(x77468, x68462, x77470);
  nand n77469(x77469, x77468, x73104);
  nand n77471(x77471, x68462, x77473);
  nand n77472(x77472, x77471, x73109);
  nand n77474(x77474, x68462, x77476);
  nand n77475(x77475, x77474, x73114);
  nand n77477(x77477, x68462, x77479);
  nand n77478(x77478, x77477, x73119);
  nand n77480(x77480, x68462, x77482);
  nand n77481(x77481, x77480, x73124);
  nand n77483(x77483, x68462, x77485);
  nand n77484(x77484, x77483, x73129);
  nand n77486(x77486, x68462, x77488);
  nand n77487(x77487, x77486, x73134);
  nand n77489(x77489, x68462, x77491);
  nand n77490(x77490, x77489, x73139);
  nand n77492(x77492, x68462, x77494);
  nand n77493(x77493, x77492, x73144);
  nand n77495(x77495, x68462, x77497);
  nand n77496(x77496, x77495, x73149);
  nand n77498(x77498, x68462, x77500);
  nand n77499(x77499, x77498, x73154);
  nand n77501(x77501, x68462, x77503);
  nand n77502(x77502, x77501, x73159);
  nand n77504(x77504, x68462, x77506);
  nand n77505(x77505, x77504, x73164);
  nand n77507(x77507, x68462, x77509);
  nand n77508(x77508, x77507, x73169);
  nand n77510(x77510, x68462, x77512);
  nand n77511(x77511, x77510, x73174);
  nand n77513(x77513, x68462, x77515);
  nand n77514(x77514, x77513, x73179);
  nand n77516(x77516, x68462, x77518);
  nand n77517(x77517, x77516, x73184);
  nand n77519(x77519, x68462, x77521);
  nand n77520(x77520, x77519, x73189);
  nand n77522(x77522, x68462, x77524);
  nand n77523(x77523, x77522, x73194);
  nand n77525(x77525, x68462, x77527);
  nand n77526(x77526, x77525, x73199);
  nand n77528(x77528, x68462, x77530);
  nand n77529(x77529, x77528, x73204);
  nand n77531(x77531, x68462, x77533);
  nand n77532(x77532, x77531, x73209);
  nand n77534(x77534, x68462, x77536);
  nand n77535(x77535, x77534, x73214);
  nand n77537(x77537, x68462, x77539);
  nand n77538(x77538, x77537, x73219);
  nand n77540(x77540, x68462, x77542);
  nand n77541(x77541, x77540, x73224);
  nand n77543(x77543, x68462, x77545);
  nand n77544(x77544, x77543, x73229);
  nand n77546(x77546, x68462, x77548);
  nand n77547(x77547, x77546, x73234);
  nand n77549(x77549, x68462, x77551);
  nand n77550(x77550, x77549, x73239);
  nand n77552(x77552, x68462, x77554);
  nand n77553(x77553, x77552, x73244);
  nand n77555(x77555, x68462, x77557);
  nand n77556(x77556, x77555, x73249);
  nand n77558(x77558, x68462, x77560);
  nand n77559(x77559, x77558, x73254);
  nand n77561(x77561, x68462, x77563);
  nand n77562(x77562, x77561, x73259);
  nand n77564(x77564, x68462, x77566);
  nand n77565(x77565, x77564, x73264);
  nand n77567(x77567, x68462, x77569);
  nand n77568(x77568, x77567, x73269);
  nand n77570(x77570, x68462, x77572);
  nand n77571(x77571, x77570, x73274);
  nand n77573(x77573, x68462, x77575);
  nand n77574(x77574, x77573, x73279);
  nand n77576(x77576, x68462, x77578);
  nand n77577(x77577, x77576, x73284);
  nand n77579(x77579, x68462, x77581);
  nand n77580(x77580, x77579, x73289);
  nand n77582(x77582, x68462, x77584);
  nand n77583(x77583, x77582, x73294);
  nand n77585(x77585, x68462, x77587);
  nand n77586(x77586, x77585, x73299);
  nand n77588(x77588, x68462, x77590);
  nand n77589(x77589, x77588, x73304);
  nand n77591(x77591, x68462, x77593);
  nand n77592(x77592, x77591, x73309);
  nand n77594(x77594, x68462, x77596);
  nand n77595(x77595, x77594, x73314);
  nand n77597(x77597, x68462, x77599);
  nand n77598(x77598, x77597, x73319);
  nand n77600(x77600, x68462, x77602);
  nand n77601(x77601, x77600, x73324);
  nand n77603(x77603, x68462, x77605);
  nand n77604(x77604, x77603, x73329);
  nand n77606(x77606, x68462, x77608);
  nand n77607(x77607, x77606, x73334);
  nand n77609(x77609, x68462, x77611);
  nand n77610(x77610, x77609, x73339);
  nand n77612(x77612, x68462, x77614);
  nand n77613(x77613, x77612, x73344);
  nand n77615(x77615, x68462, x77617);
  nand n77616(x77616, x77615, x73349);
  nand n77618(x77618, x68462, x77620);
  nand n77619(x77619, x77618, x73354);
  nand n77621(x77621, x68462, x77623);
  nand n77622(x77622, x77621, x73359);
  nand n77624(x77624, x68462, x77626);
  nand n77625(x77625, x77624, x73364);
  nand n77627(x77627, x68462, x77629);
  nand n77628(x77628, x77627, x73369);
  nand n77630(x77630, x68462, x77632);
  nand n77631(x77631, x77630, x73374);
  nand n77633(x77633, x68462, x77635);
  nand n77634(x77634, x77633, x73379);
  nand n77636(x77636, x68462, x77638);
  nand n77637(x77637, x77636, x73384);
  nand n77639(x77639, x68462, x77641);
  nand n77640(x77640, x77639, x73389);
  nand n77642(x77642, x68462, x77644);
  nand n77643(x77643, x77642, x73394);
  nand n77645(x77645, x68462, x77647);
  nand n77646(x77646, x77645, x73399);
  nand n77648(x77648, x68462, x77650);
  nand n77649(x77649, x77648, x73404);
  nand n77651(x77651, x68462, x77653);
  nand n77652(x77652, x77651, x73409);
  nand n77654(x77654, x68462, x77656);
  nand n77655(x77655, x77654, x73414);
  nand n77657(x77657, x68462, x77659);
  nand n77658(x77658, x77657, x73419);
  nand n77660(x77660, x68462, x77662);
  nand n77661(x77661, x77660, x73424);
  nand n77663(x77663, x68462, x77665);
  nand n77664(x77664, x77663, x73429);
  nand n77666(x77666, x68462, x77668);
  nand n77667(x77667, x77666, x73434);
  nand n77669(x77669, x68462, x77671);
  nand n77670(x77670, x77669, x73439);
  nand n77672(x77672, x68462, x77674);
  nand n77673(x77673, x77672, x73444);
  nand n77675(x77675, x68462, x77677);
  nand n77676(x77676, x77675, x73449);
  nand n77678(x77678, x68462, x77680);
  nand n77679(x77679, x77678, x73454);
  nand n77681(x77681, x68462, x77683);
  nand n77682(x77682, x77681, x73459);
  nand n77684(x77684, x68462, x77686);
  nand n77685(x77685, x77684, x73464);
  nand n77687(x77687, x68462, x77689);
  nand n77688(x77688, x77687, x73469);
  nand n77690(x77690, x68462, x77692);
  nand n77691(x77691, x77690, x73474);
  nand n77693(x77693, x68462, x77695);
  nand n77694(x77694, x77693, x73479);
  nand n77696(x77696, x68462, x77698);
  nand n77697(x77697, x77696, x73484);
  nand n77699(x77699, x68462, x77701);
  nand n77700(x77700, x77699, x73489);
  nand n77702(x77702, x68462, x77704);
  nand n77703(x77703, x77702, x73494);
  nand n77705(x77705, x68462, x77707);
  nand n77706(x77706, x77705, x73499);
  nand n77708(x77708, x68462, x77710);
  nand n77709(x77709, x77708, x73504);
  nand n77711(x77711, x68462, x77713);
  nand n77712(x77712, x77711, x73509);
  nand n77714(x77714, x68462, x77716);
  nand n77715(x77715, x77714, x73514);
  nand n77717(x77717, x68462, x77719);
  nand n77718(x77718, x77717, x73519);
  nand n77720(x77720, x68462, x77722);
  nand n77721(x77721, x77720, x73524);
  nand n77723(x77723, x68462, x77725);
  nand n77724(x77724, x77723, x73529);
  nand n77726(x77726, x68462, x77728);
  nand n77727(x77727, x77726, x73534);
  nand n77729(x77729, x68462, x77731);
  nand n77730(x77730, x77729, x73539);
  nand n77732(x77732, x68462, x77734);
  nand n77733(x77733, x77732, x73544);
  nand n77735(x77735, x68462, x77737);
  nand n77736(x77736, x77735, x73549);
  nand n77738(x77738, x68462, x77740);
  nand n77739(x77739, x77738, x73554);
  nand n77741(x77741, x68462, x77743);
  nand n77742(x77742, x77741, x73559);
  nand n77744(x77744, x68462, x77746);
  nand n77745(x77745, x77744, x73564);
  nand n77747(x77747, x68462, x77749);
  nand n77748(x77748, x77747, x73569);
  nand n77750(x77750, x68462, x77752);
  nand n77751(x77751, x77750, x73574);
  nand n77753(x77753, x68462, x77755);
  nand n77754(x77754, x77753, x73579);
  nand n77756(x77756, x68462, x77758);
  nand n77757(x77757, x77756, x73584);
  nand n77759(x77759, x68462, x77761);
  nand n77760(x77760, x77759, x73589);
  nand n77762(x77762, x68462, x77764);
  nand n77763(x77763, x77762, x73594);
  nand n77765(x77765, x68462, x77767);
  nand n77766(x77766, x77765, x73599);
  nand n77768(x77768, x68462, x77770);
  nand n77769(x77769, x77768, x73604);
  nand n77771(x77771, x68462, x77773);
  nand n77772(x77772, x77771, x73609);
  nand n77774(x77774, x68462, x77776);
  nand n77775(x77775, x77774, x73614);
  nand n77777(x77777, x68462, x77779);
  nand n77778(x77778, x77777, x73619);
  nand n77780(x77780, x68462, x77782);
  nand n77781(x77781, x77780, x73624);
  nand n77783(x77783, x68462, x77785);
  nand n77784(x77784, x77783, x73629);
  nand n77786(x77786, x68462, x77788);
  nand n77787(x77787, x77786, x73634);
  nand n77789(x77789, x68462, x77791);
  nand n77790(x77790, x77789, x73639);
  nand n77792(x77792, x68462, x77794);
  nand n77793(x77793, x77792, x73644);
  nand n77795(x77795, x68462, x77797);
  nand n77796(x77796, x77795, x73649);
  nand n77798(x77798, x68462, x77800);
  nand n77799(x77799, x77798, x73654);
  nand n77801(x77801, x68462, x77803);
  nand n77802(x77802, x77801, x73659);
  nand n77804(x77804, x68462, x77806);
  nand n77805(x77805, x77804, x73664);
  nand n77807(x77807, x68462, x77809);
  nand n77808(x77808, x77807, x73669);
  nand n77810(x77810, x68462, x77812);
  nand n77811(x77811, x77810, x73674);
  nand n77813(x77813, x68462, x77815);
  nand n77814(x77814, x77813, x73679);
  nand n77816(x77816, x68462, x77818);
  nand n77817(x77817, x77816, x73684);
  nand n77819(x77819, x68462, x77821);
  nand n77820(x77820, x77819, x73689);
  nand n77822(x77822, x68462, x77824);
  nand n77823(x77823, x77822, x73694);
  nand n77825(x77825, x68462, x77827);
  nand n77826(x77826, x77825, x73699);
  nand n77828(x77828, x68462, x77830);
  nand n77829(x77829, x77828, x73704);
  nand n77831(x77831, x68462, x77833);
  nand n77832(x77832, x77831, x73709);
  nand n77834(x77834, x68462, x77836);
  nand n77835(x77835, x77834, x73714);
  nand n77837(x77837, x68462, x77839);
  nand n77838(x77838, x77837, x73719);
  nand n77840(x77840, x68462, x77842);
  nand n77841(x77841, x77840, x73724);
  nand n77843(x77843, x68462, x77845);
  nand n77844(x77844, x77843, x73729);
  nand n77846(x77846, x68462, x77848);
  nand n77847(x77847, x77846, x73734);
  nand n77849(x77849, x68462, x77851);
  nand n77850(x77850, x77849, x73739);
  nand n77852(x77852, x68462, x77854);
  nand n77853(x77853, x77852, x73744);
  nand n77855(x77855, x68462, x77857);
  nand n77856(x77856, x77855, x73749);
  nand n77858(x77858, x68462, x77860);
  nand n77859(x77859, x77858, x73754);
  nand n77861(x77861, x68462, x77863);
  nand n77862(x77862, x77861, x73759);
  nand n77864(x77864, x68462, x77866);
  nand n77865(x77865, x77864, x73764);
  nand n77867(x77867, x68462, x77869);
  nand n77868(x77868, x77867, x73769);
  nand n77870(x77870, x68462, x77872);
  nand n77871(x77871, x77870, x73774);
  nand n77873(x77873, x68462, x77875);
  nand n77874(x77874, x77873, x73779);
  nand n77876(x77876, x68462, x77878);
  nand n77877(x77877, x77876, x73784);
  nand n77879(x77879, x68462, x77881);
  nand n77880(x77880, x77879, x73789);
  nand n77882(x77882, x68462, x77884);
  nand n77883(x77883, x77882, x73794);
  nand n77885(x77885, x68462, x77887);
  nand n77886(x77886, x77885, x73799);
  nand n77888(x77888, x68462, x77890);
  nand n77889(x77889, x77888, x73804);
  nand n77891(x77891, x68462, x77893);
  nand n77892(x77892, x77891, x73809);
  nand n77894(x77894, x68462, x77896);
  nand n77895(x77895, x77894, x73814);
  nand n77897(x77897, x68462, x77899);
  nand n77898(x77898, x77897, x73819);
  nand n77900(x77900, x68462, x77902);
  nand n77901(x77901, x77900, x73824);
  nand n77903(x77903, x68462, x77905);
  nand n77904(x77904, x77903, x73829);
  nand n77906(x77906, x68462, x77908);
  nand n77907(x77907, x77906, x73834);
  nand n77909(x77909, x68462, x77911);
  nand n77910(x77910, x77909, x73839);
  nand n77912(x77912, x68462, x77914);
  nand n77913(x77913, x77912, x73844);
  nand n77915(x77915, x68462, x77917);
  nand n77916(x77916, x77915, x73849);
  nand n77918(x77918, x68462, x77920);
  nand n77919(x77919, x77918, x73854);
  nand n77921(x77921, x68462, x77923);
  nand n77922(x77922, x77921, x73859);
  nand n77924(x77924, x68462, x77926);
  nand n77925(x77925, x77924, x73864);
  nand n77927(x77927, x68462, x77929);
  nand n77928(x77928, x77927, x73869);
  nand n77930(x77930, x68462, x77932);
  nand n77931(x77931, x77930, x73874);
  nand n77933(x77933, x68462, x77935);
  nand n77934(x77934, x77933, x73879);
  nand n77936(x77936, x68462, x77938);
  nand n77937(x77937, x77936, x73884);
  nand n77939(x77939, x68462, x77941);
  nand n77940(x77940, x77939, x73889);
  nand n77942(x77942, x68462, x77944);
  nand n77943(x77943, x77942, x73894);
  nand n77945(x77945, x68462, x77947);
  nand n77946(x77946, x77945, x73899);
  nand n77948(x77948, x68462, x77950);
  nand n77949(x77949, x77948, x73904);
  nand n77951(x77951, x68462, x77953);
  nand n77952(x77952, x77951, x73909);
  nand n77954(x77954, x68462, x77956);
  nand n77955(x77955, x77954, x73914);
  nand n77957(x77957, x68462, x77959);
  nand n77958(x77958, x77957, x73919);
  nand n77960(x77960, x68462, x77962);
  nand n77961(x77961, x77960, x73924);
  nand n77963(x77963, x68462, x77965);
  nand n77964(x77964, x77963, x73929);
  nand n77966(x77966, x68462, x77968);
  nand n77967(x77967, x77966, x73934);
  nand n77969(x77969, x68462, x77971);
  nand n77970(x77970, x77969, x73939);
  nand n77972(x77972, x68462, x77974);
  nand n77973(x77973, x77972, x73944);
  nand n77975(x77975, x68462, x77977);
  nand n77976(x77976, x77975, x73949);
  nand n77978(x77978, x68462, x77980);
  nand n77979(x77979, x77978, x73954);
  nand n77981(x77981, x68462, x77983);
  nand n77982(x77982, x77981, x73959);
  nand n77984(x77984, x68462, x77986);
  nand n77985(x77985, x77984, x73964);
  nand n77987(x77987, x68462, x77989);
  nand n77988(x77988, x77987, x73969);
  nand n77990(x77990, x68462, x77992);
  nand n77991(x77991, x77990, x73974);
  nand n77993(x77993, x68462, x77995);
  nand n77994(x77994, x77993, x73979);
  nand n77996(x77996, x68462, x77998);
  nand n77997(x77997, x77996, x73984);
  nand n77999(x77999, x68462, x78001);
  nand n78000(x78000, x77999, x73989);
  nand n78002(x78002, x68462, x78004);
  nand n78003(x78003, x78002, x73994);
  nand n78005(x78005, x68462, x78007);
  nand n78006(x78006, x78005, x73999);
  nand n78008(x78008, x68462, x78010);
  nand n78009(x78009, x78008, x71799);
  nand n78011(x78011, x68462, x78013);
  nand n78012(x78012, x78011, x71804);
  nand n78014(x78014, x68462, x78016);
  nand n78015(x78015, x78014, x71809);
  nand n78017(x78017, x68462, x78019);
  nand n78018(x78018, x78017, x71814);
  nand n78020(x78020, x68462, x78022);
  nand n78021(x78021, x78020, x71819);
  nand n78023(x78023, x68462, x78025);
  nand n78024(x78024, x78023, x71824);
  nand n78026(x78026, x68462, x78028);
  nand n78027(x78027, x78026, x71829);
  nand n78029(x78029, x68462, x78031);
  nand n78030(x78030, x78029, x71834);
  nand n78032(x78032, x68462, x78034);
  nand n78033(x78033, x78032, x71839);
  nand n78035(x78035, x68462, x78037);
  nand n78036(x78036, x78035, x71844);
  nand n78038(x78038, x68462, x78040);
  nand n78039(x78039, x78038, x71849);
  nand n78041(x78041, x68462, x78043);
  nand n78042(x78042, x78041, x71854);
  nand n78044(x78044, x68462, x78046);
  nand n78045(x78045, x78044, x71859);
  nand n78047(x78047, x68462, x78049);
  nand n78048(x78048, x78047, x71864);
  nand n78050(x78050, x68462, x78052);
  nand n78051(x78051, x78050, x71869);
  nand n78053(x78053, x68462, x78055);
  nand n78054(x78054, x78053, x71874);
  nand n78056(x78056, x68462, x78058);
  nand n78057(x78057, x78056, x71879);
  nand n78059(x78059, x68462, x78061);
  nand n78060(x78060, x78059, x71884);
  nand n78062(x78062, x68462, x78064);
  nand n78063(x78063, x78062, x71889);
  nand n78065(x78065, x68462, x78067);
  nand n78066(x78066, x78065, x71894);
  nand n78068(x78068, x68462, x78070);
  nand n78069(x78069, x78068, x71899);
  nand n78071(x78071, x68462, x78073);
  nand n78072(x78072, x78071, x71904);
  nand n78074(x78074, x68462, x78076);
  nand n78075(x78075, x78074, x71904);
  nand n78077(x78077, x68462, x78079);
  nand n78078(x78078, x78077, x71904);
  nand n78080(x78080, x68462, x78082);
  nand n78081(x78081, x78080, x71904);
  nand n78083(x78083, x68462, x78085);
  nand n78084(x78084, x78083, x71904);
  nand n78086(x78086, x68462, x78088);
  nand n78087(x78087, x78086, x71904);
  nand n78089(x78089, x68462, x78091);
  nand n78090(x78090, x78089, x71904);
  nand n78092(x78092, x68462, x78094);
  nand n78093(x78093, x78092, x71904);
  nand n78095(x78095, x68462, x78097);
  nand n78096(x78096, x78095, x71904);
  nand n78098(x78098, x68462, x78100);
  nand n78099(x78099, x78098, x71904);
  nand n78101(x78101, x68462, x78103);
  nand n78102(x78102, x78101, x71904);
  nand n78104(x78104, x68462, x78106);
  nand n78105(x78105, x78104, x71939);
  nand n78107(x78107, x68462, x78109);
  nand n78108(x78108, x78107, x71944);
  nand n78110(x78110, x68462, x78112);
  nand n78111(x78111, x78110, x71949);
  nand n78113(x78113, x68462, x78115);
  nand n78114(x78114, x78113, x71954);
  nand n78116(x78116, x68462, x78118);
  nand n78117(x78117, x78116, x71959);
  nand n78119(x78119, x68462, x78121);
  nand n78120(x78120, x78119, x71964);
  nand n78122(x78122, x68462, x78124);
  nand n78123(x78123, x78122, x71969);
  nand n78125(x78125, x68462, x78127);
  nand n78126(x78126, x78125, x71974);
  nand n78128(x78128, x68462, x78130);
  nand n78129(x78129, x78128, x71979);
  nand n78131(x78131, x68462, x78133);
  nand n78132(x78132, x78131, x71984);
  nand n78134(x78134, x68462, x78136);
  nand n78135(x78135, x78134, x71989);
  nand n78137(x78137, x68462, x78139);
  nand n78138(x78138, x78137, x71994);
  nand n78140(x78140, x68462, x78142);
  nand n78141(x78141, x78140, x71999);
  nand n78143(x78143, x68462, x78145);
  nand n78144(x78144, x78143, x72004);
  nand n78146(x78146, x68462, x78148);
  nand n78147(x78147, x78146, x72009);
  nand n78149(x78149, x68462, x78151);
  nand n78150(x78150, x78149, x72014);
  nand n78152(x78152, x68462, x78154);
  nand n78153(x78153, x78152, x72019);
  nand n78155(x78155, x68462, x78157);
  nand n78156(x78156, x78155, x72024);
  nand n78158(x78158, x68462, x78160);
  nand n78159(x78159, x78158, x72029);
  nand n78161(x78161, x68462, x78163);
  nand n78162(x78162, x78161, x72034);
  nand n78164(x78164, x68462, x78166);
  nand n78165(x78165, x78164, x72039);
  nand n78167(x78167, x68462, x78169);
  nand n78168(x78168, x78167, x72044);
  nand n78170(x78170, x68462, x78172);
  nand n78171(x78171, x78170, x72049);
  nand n78173(x78173, x68462, x78175);
  nand n78174(x78174, x78173, x72054);
  nand n78176(x78176, x68462, x78178);
  nand n78177(x78177, x78176, x72059);
  nand n78179(x78179, x68462, x78181);
  nand n78180(x78180, x78179, x72064);
  nand n78182(x78182, x68462, x78184);
  nand n78183(x78183, x78182, x72069);
  nand n78185(x78185, x68462, x78187);
  nand n78186(x78186, x78185, x72074);
  nand n78188(x78188, x68462, x78190);
  nand n78189(x78189, x78188, x72079);
  nand n78191(x78191, x68462, x78193);
  nand n78192(x78192, x78191, x72084);
  nand n78194(x78194, x68462, x78196);
  nand n78195(x78195, x78194, x72089);
  nand n78197(x78197, x68462, x78199);
  nand n78198(x78198, x78197, x72094);
  nand n78200(x78200, x68462, x78202);
  nand n78201(x78201, x78200, x72099);
  nand n78203(x78203, x68462, x78205);
  nand n78204(x78204, x78203, x72104);
  nand n78206(x78206, x68462, x78208);
  nand n78207(x78207, x78206, x72109);
  nand n78209(x78209, x68462, x78211);
  nand n78210(x78210, x78209, x72114);
  nand n78212(x78212, x68462, x78214);
  nand n78213(x78213, x78212, x72119);
  nand n78215(x78215, x68462, x78217);
  nand n78216(x78216, x78215, x72124);
  nand n78218(x78218, x68462, x78220);
  nand n78219(x78219, x78218, x72129);
  nand n78221(x78221, x68462, x78223);
  nand n78222(x78222, x78221, x72134);
  nand n78224(x78224, x68462, x78226);
  nand n78225(x78225, x78224, x72139);
  nand n78227(x78227, x68462, x78229);
  nand n78228(x78228, x78227, x72144);
  nand n78230(x78230, x68462, x78232);
  nand n78231(x78231, x78230, x72149);
  nand n78233(x78233, x68462, x78235);
  nand n78234(x78234, x78233, x72154);
  nand n78236(x78236, x68462, x78238);
  nand n78237(x78237, x78236, x72159);
  nand n78239(x78239, x68462, x78241);
  nand n78240(x78240, x78239, x72164);
  nand n78242(x78242, x68462, x78244);
  nand n78243(x78243, x78242, x72169);
  nand n78245(x78245, x68462, x78247);
  nand n78246(x78246, x78245, x72174);
  nand n78248(x78248, x68462, x78250);
  nand n78249(x78249, x78248, x72179);
  nand n78251(x78251, x68462, x78253);
  nand n78252(x78252, x78251, x72184);
  nand n78254(x78254, x68462, x78256);
  nand n78255(x78255, x78254, x72189);
  nand n78257(x78257, x68462, x78259);
  nand n78258(x78258, x78257, x72194);
  nand n78260(x78260, x68462, x78262);
  nand n78261(x78261, x78260, x72199);
  nand n78263(x78263, x68462, x78265);
  nand n78264(x78264, x78263, x72204);
  nand n78266(x78266, x68462, x78268);
  nand n78267(x78267, x78266, x72209);
  nand n78269(x78269, x68462, x78271);
  nand n78270(x78270, x78269, x72214);
  nand n78272(x78272, x68462, x78274);
  nand n78273(x78273, x78272, x72219);
  nand n78275(x78275, x68462, x78277);
  nand n78276(x78276, x78275, x72224);
  nand n78278(x78278, x68462, x78280);
  nand n78279(x78279, x78278, x72229);
  nand n78281(x78281, x68462, x78283);
  nand n78282(x78282, x78281, x72234);
  nand n78284(x78284, x68462, x78286);
  nand n78285(x78285, x78284, x72239);
  nand n78287(x78287, x68462, x78289);
  nand n78288(x78288, x78287, x72244);
  nand n78290(x78290, x68462, x78292);
  nand n78291(x78291, x78290, x72249);
  nand n78293(x78293, x68462, x78295);
  nand n78294(x78294, x78293, x72254);
  nand n78296(x78296, x68462, x78298);
  nand n78297(x78297, x78296, x72259);
  nand n78299(x78299, x68462, x78301);
  nand n78300(x78300, x78299, x72264);
  nand n78302(x78302, x68462, x78304);
  nand n78303(x78303, x78302, x72269);
  nand n78305(x78305, x68462, x78307);
  nand n78306(x78306, x78305, x72274);
  nand n78308(x78308, x68462, x78310);
  nand n78309(x78309, x78308, x72279);
  nand n78311(x78311, x68462, x78313);
  nand n78312(x78312, x78311, x72284);
  nand n78314(x78314, x68462, x78316);
  nand n78315(x78315, x78314, x72289);
  nand n78317(x78317, x68462, x78319);
  nand n78318(x78318, x78317, x72294);
  nand n78320(x78320, x68462, x78322);
  nand n78321(x78321, x78320, x72299);
  nand n78323(x78323, x68462, x78325);
  nand n78324(x78324, x78323, x72304);
  nand n78326(x78326, x68462, x78328);
  nand n78327(x78327, x78326, x72309);
  nand n78329(x78329, x68462, x78331);
  nand n78330(x78330, x78329, x72314);
  nand n78332(x78332, x68462, x78334);
  nand n78333(x78333, x78332, x72319);
  nand n78335(x78335, x68462, x78337);
  nand n78336(x78336, x78335, x72324);
  nand n78338(x78338, x68462, x78340);
  nand n78339(x78339, x78338, x72329);
  nand n78341(x78341, x68462, x78343);
  nand n78342(x78342, x78341, x72334);
  nand n78344(x78344, x68462, x78346);
  nand n78345(x78345, x78344, x72339);
  nand n78347(x78347, x68462, x78349);
  nand n78348(x78348, x78347, x72344);
  nand n78350(x78350, x68462, x78352);
  nand n78351(x78351, x78350, x72349);
  nand n78353(x78353, x68462, x78355);
  nand n78354(x78354, x78353, x72354);
  nand n78356(x78356, x68462, x78358);
  nand n78357(x78357, x78356, x72359);
  nand n78359(x78359, x68462, x78361);
  nand n78360(x78360, x78359, x72364);
  nand n78362(x78362, x68462, x78364);
  nand n78363(x78363, x78362, x72369);
  nand n78365(x78365, x68462, x78367);
  nand n78366(x78366, x78365, x72374);
  nand n78368(x78368, x68462, x78370);
  nand n78369(x78369, x78368, x72379);
  nand n78371(x78371, x68462, x78373);
  nand n78372(x78372, x78371, x72384);
  nand n78374(x78374, x68462, x78376);
  nand n78375(x78375, x78374, x72389);
  nand n78377(x78377, x68462, x78379);
  nand n78378(x78378, x78377, x72394);
  nand n78380(x78380, x68462, x78382);
  nand n78381(x78381, x78380, x72399);
  nand n78383(x78383, x68462, x78385);
  nand n78384(x78384, x78383, x72404);
  nand n78386(x78386, x68462, x78388);
  nand n78387(x78387, x78386, x72409);
  nand n78389(x78389, x68462, x78391);
  nand n78390(x78390, x78389, x72414);
  nand n78392(x78392, x68462, x78394);
  nand n78393(x78393, x78392, x72419);
  nand n78395(x78395, x68462, x78397);
  nand n78396(x78396, x78395, x72424);
  nand n78398(x78398, x68462, x78400);
  nand n78399(x78399, x78398, x72429);
  nand n78401(x78401, x68462, x78403);
  nand n78402(x78402, x78401, x72434);
  nand n78404(x78404, x68462, x78406);
  nand n78405(x78405, x78404, x72439);
  nand n78407(x78407, x68462, x78409);
  nand n78408(x78408, x78407, x72444);
  nand n78410(x78410, x68462, x78412);
  nand n78411(x78411, x78410, x72449);
  nand n78413(x78413, x68462, x78415);
  nand n78414(x78414, x78413, x72454);
  nand n78416(x78416, x68462, x78418);
  nand n78417(x78417, x78416, x72459);
  nand n78419(x78419, x68462, x78421);
  nand n78420(x78420, x78419, x72464);
  nand n78422(x78422, x68462, x78424);
  nand n78423(x78423, x78422, x72469);
  nand n78425(x78425, x68462, x78427);
  nand n78426(x78426, x78425, x72474);
  nand n78428(x78428, x68462, x78430);
  nand n78429(x78429, x78428, x72479);
  nand n78431(x78431, x68462, x78433);
  nand n78432(x78432, x78431, x72484);
  nand n78434(x78434, x68462, x78436);
  nand n78435(x78435, x78434, x72489);
  nand n78437(x78437, x68462, x78439);
  nand n78438(x78438, x78437, x72494);
  nand n78440(x78440, x68462, x78442);
  nand n78441(x78441, x78440, x72499);
  nand n78443(x78443, x68462, x78445);
  nand n78444(x78444, x78443, x72504);
  nand n78446(x78446, x68462, x78448);
  nand n78447(x78447, x78446, x72509);
  nand n78449(x78449, x68462, x78451);
  nand n78450(x78450, x78449, x72514);
  nand n78452(x78452, x68462, x78454);
  nand n78453(x78453, x78452, x72519);
  nand n78455(x78455, x68462, x78457);
  nand n78456(x78456, x78455, x72524);
  nand n78458(x78458, x68462, x78460);
  nand n78459(x78459, x78458, x72529);
  nand n78461(x78461, x68462, x78463);
  nand n78462(x78462, x78461, x72534);
  nand n78464(x78464, x68462, x78466);
  nand n78465(x78465, x78464, x72539);
  nand n78467(x78467, x68462, x78469);
  nand n78468(x78468, x78467, x72544);
  nand n78470(x78470, x68462, x78472);
  nand n78471(x78471, x78470, x72549);
  nand n78473(x78473, x68462, x78475);
  nand n78474(x78474, x78473, x72554);
  nand n78476(x78476, x68462, x78478);
  nand n78477(x78477, x78476, x72559);
  nand n78479(x78479, x68462, x78481);
  nand n78480(x78480, x78479, x72564);
  nand n78482(x78482, x68462, x78484);
  nand n78483(x78483, x78482, x72569);
  nand n78485(x78485, x68462, x78487);
  nand n78486(x78486, x78485, x72574);
  nand n78488(x78488, x68462, x78490);
  nand n78489(x78489, x78488, x72579);
  nand n78491(x78491, x68462, x78493);
  nand n78492(x78492, x78491, x72584);
  nand n78494(x78494, x68462, x78496);
  nand n78495(x78495, x78494, x72589);
  nand n78497(x78497, x68462, x78499);
  nand n78498(x78498, x78497, x72594);
  nand n78500(x78500, x68462, x78502);
  nand n78501(x78501, x78500, x72599);
  nand n78503(x78503, x68462, x78505);
  nand n78504(x78504, x78503, x72604);
  nand n78506(x78506, x68462, x78508);
  nand n78507(x78507, x78506, x72609);
  nand n78509(x78509, x68462, x78511);
  nand n78510(x78510, x78509, x72614);
  nand n78512(x78512, x68462, x78514);
  nand n78513(x78513, x78512, x72619);
  nand n78515(x78515, x68462, x78517);
  nand n78516(x78516, x78515, x72624);
  nand n78518(x78518, x68462, x78520);
  nand n78519(x78519, x78518, x72629);
  nand n78521(x78521, x68462, x78523);
  nand n78522(x78522, x78521, x72634);
  nand n78524(x78524, x68462, x78526);
  nand n78525(x78525, x78524, x72639);
  nand n78527(x78527, x68462, x78529);
  nand n78528(x78528, x78527, x72644);
  nand n78530(x78530, x68462, x78532);
  nand n78531(x78531, x78530, x72649);
  nand n78533(x78533, x68462, x78535);
  nand n78534(x78534, x78533, x72654);
  nand n78536(x78536, x68462, x78538);
  nand n78537(x78537, x78536, x72659);
  nand n78539(x78539, x68462, x78541);
  nand n78540(x78540, x78539, x72664);
  nand n78542(x78542, x68462, x78544);
  nand n78543(x78543, x78542, x72669);
  nand n78545(x78545, x68462, x78547);
  nand n78546(x78546, x78545, x72674);
  nand n78548(x78548, x68462, x78550);
  nand n78549(x78549, x78548, x72679);
  nand n78551(x78551, x68462, x78553);
  nand n78552(x78552, x78551, x72684);
  nand n78554(x78554, x68462, x78556);
  nand n78555(x78555, x78554, x72689);
  nand n78557(x78557, x68462, x78559);
  nand n78558(x78558, x78557, x72694);
  nand n78560(x78560, x68462, x78562);
  nand n78561(x78561, x78560, x72699);
  nand n78563(x78563, x68462, x78565);
  nand n78564(x78564, x78563, x72704);
  nand n78566(x78566, x68462, x78568);
  nand n78567(x78567, x78566, x72709);
  nand n78569(x78569, x68462, x78571);
  nand n78570(x78570, x78569, x72714);
  nand n78572(x78572, x68462, x78574);
  nand n78573(x78573, x78572, x72719);
  nand n78575(x78575, x68462, x78577);
  nand n78576(x78576, x78575, x72724);
  nand n78578(x78578, x68462, x78580);
  nand n78579(x78579, x78578, x72729);
  nand n78581(x78581, x68462, x78583);
  nand n78582(x78582, x78581, x72734);
  nand n78584(x78584, x68462, x78586);
  nand n78585(x78585, x78584, x72739);
  nand n78587(x78587, x68462, x78589);
  nand n78588(x78588, x78587, x72744);
  nand n78590(x78590, x68462, x78592);
  nand n78591(x78591, x78590, x72749);
  nand n78593(x78593, x68462, x78595);
  nand n78594(x78594, x78593, x72754);
  nand n78596(x78596, x68462, x78598);
  nand n78597(x78597, x78596, x72759);
  nand n78599(x78599, x68462, x78601);
  nand n78600(x78600, x78599, x72764);
  nand n78602(x78602, x68462, x78604);
  nand n78603(x78603, x78602, x72769);
  nand n78605(x78605, x68462, x78607);
  nand n78606(x78606, x78605, x72774);
  nand n78608(x78608, x68462, x78610);
  nand n78609(x78609, x78608, x72779);
  nand n78611(x78611, x68462, x78613);
  nand n78612(x78612, x78611, x72784);
  nand n78614(x78614, x68462, x78616);
  nand n78615(x78615, x78614, x72789);
  nand n78617(x78617, x68462, x78619);
  nand n78618(x78618, x78617, x72794);
  nand n78620(x78620, x68462, x78622);
  nand n78621(x78621, x78620, x72799);
  nand n78623(x78623, x68462, x78625);
  nand n78624(x78624, x78623, x72804);
  nand n78626(x78626, x68462, x78628);
  nand n78627(x78627, x78626, x72809);
  nand n78629(x78629, x68462, x78631);
  nand n78630(x78630, x78629, x72814);
  nand n78632(x78632, x68462, x78634);
  nand n78633(x78633, x78632, x72819);
  nand n78635(x78635, x68462, x78637);
  nand n78636(x78636, x78635, x72824);
  nand n78638(x78638, x68462, x78640);
  nand n78639(x78639, x78638, x72829);
  nand n78641(x78641, x68462, x78643);
  nand n78642(x78642, x78641, x72834);
  nand n78644(x78644, x68462, x78646);
  nand n78645(x78645, x78644, x72839);
  nand n78647(x78647, x68462, x78649);
  nand n78648(x78648, x78647, x72844);
  nand n78650(x78650, x68462, x78652);
  nand n78651(x78651, x78650, x72849);
  nand n78653(x78653, x68462, x78655);
  nand n78654(x78654, x78653, x72854);
  nand n78656(x78656, x68462, x78658);
  nand n78657(x78657, x78656, x72859);
  nand n78659(x78659, x68462, x78661);
  nand n78660(x78660, x78659, x72864);
  nand n78662(x78662, x68462, x78664);
  nand n78663(x78663, x78662, x72869);
  nand n78665(x78665, x68462, x78667);
  nand n78666(x78666, x78665, x72874);
  nand n78668(x78668, x68462, x78670);
  nand n78669(x78669, x78668, x72879);
  nand n78671(x78671, x68462, x78673);
  nand n78672(x78672, x78671, x72884);
  nand n78674(x78674, x68462, x78676);
  nand n78675(x78675, x78674, x72889);
  nand n78677(x78677, x68462, x78679);
  nand n78678(x78678, x78677, x72894);
  nand n78680(x78680, x68462, x78682);
  nand n78681(x78681, x78680, x72899);
  nand n78683(x78683, x68462, x78685);
  nand n78684(x78684, x78683, x72904);
  nand n78686(x78686, x68462, x78688);
  nand n78687(x78687, x78686, x72909);
  nand n78689(x78689, x68462, x78691);
  nand n78690(x78690, x78689, x72914);
  nand n78692(x78692, x68462, x78694);
  nand n78693(x78693, x78692, x72919);
  nand n78695(x78695, x68462, x78697);
  nand n78696(x78696, x78695, x72924);
  nand n78698(x78698, x68462, x78700);
  nand n78699(x78699, x78698, x72929);
  nand n78701(x78701, x68462, x78703);
  nand n78702(x78702, x78701, x72934);
  nand n78704(x78704, x68462, x78706);
  nand n78705(x78705, x78704, x72939);
  nand n78707(x78707, x68462, x78709);
  nand n78708(x78708, x78707, x72944);
  nand n78710(x78710, x68462, x78712);
  nand n78711(x78711, x78710, x72949);
  nand n78713(x78713, x68462, x78715);
  nand n78714(x78714, x78713, x72954);
  nand n78716(x78716, x68462, x78718);
  nand n78717(x78717, x78716, x72959);
  nand n78719(x78719, x68462, x78721);
  nand n78720(x78720, x78719, x72964);
  nand n78722(x78722, x68462, x78724);
  nand n78723(x78723, x78722, x72969);
  nand n78725(x78725, x68462, x78727);
  nand n78726(x78726, x78725, x72974);
  nand n78728(x78728, x68462, x78730);
  nand n78729(x78729, x78728, x72979);
  nand n78731(x78731, x68462, x78733);
  nand n78732(x78732, x78731, x72984);
  nand n78734(x78734, x68462, x78736);
  nand n78735(x78735, x78734, x72989);
  nand n78737(x78737, x68462, x78739);
  nand n78738(x78738, x78737, x72994);
  nand n78740(x78740, x68462, x78742);
  nand n78741(x78741, x78740, x72999);
  nand n78743(x78743, x68462, x78745);
  nand n78744(x78744, x78743, x73004);
  nand n78746(x78746, x68462, x78748);
  nand n78747(x78747, x78746, x73009);
  nand n78749(x78749, x68462, x78751);
  nand n78750(x78750, x78749, x73014);
  nand n78752(x78752, x68462, x78754);
  nand n78753(x78753, x78752, x73019);
  nand n78755(x78755, x68462, x78757);
  nand n78756(x78756, x78755, x73024);
  nand n78758(x78758, x68462, x78760);
  nand n78759(x78759, x78758, x73029);
  nand n78761(x78761, x68462, x78763);
  nand n78762(x78762, x78761, x73034);
  nand n78764(x78764, x68462, x78766);
  nand n78765(x78765, x78764, x73039);
  nand n78767(x78767, x68462, x78769);
  nand n78768(x78768, x78767, x73044);
  nand n78770(x78770, x68462, x78772);
  nand n78771(x78771, x78770, x73049);
  nand n78773(x78773, x68462, x78775);
  nand n78774(x78774, x78773, x73054);
  nand n78776(x78776, x68462, x78778);
  nand n78777(x78777, x78776, x73059);
  nand n78779(x78779, x68462, x78781);
  nand n78780(x78780, x78779, x73064);
  nand n78782(x78782, x68462, x78784);
  nand n78783(x78783, x78782, x73069);
  nand n78785(x78785, x68462, x78787);
  nand n78786(x78786, x78785, x73074);
  nand n78788(x78788, x68462, x78790);
  nand n78789(x78789, x78788, x73079);
  nand n78791(x78791, x68462, x78793);
  nand n78792(x78792, x78791, x73084);
  nand n78794(x78794, x68462, x78796);
  nand n78795(x78795, x78794, x73089);
  nand n78797(x78797, x68462, x78799);
  nand n78798(x78798, x78797, x73094);
  nand n78800(x78800, x68462, x78802);
  nand n78801(x78801, x78800, x73099);
  nand n78803(x78803, x68462, x78805);
  nand n78804(x78804, x78803, x73104);
  nand n78806(x78806, x68462, x78808);
  nand n78807(x78807, x78806, x73109);
  nand n78809(x78809, x68462, x78811);
  nand n78810(x78810, x78809, x73114);
  nand n78812(x78812, x68462, x78814);
  nand n78813(x78813, x78812, x73119);
  nand n78815(x78815, x68462, x78817);
  nand n78816(x78816, x78815, x73124);
  nand n78818(x78818, x68462, x78820);
  nand n78819(x78819, x78818, x73129);
  nand n78821(x78821, x68462, x78823);
  nand n78822(x78822, x78821, x73134);
  nand n78824(x78824, x68462, x78826);
  nand n78825(x78825, x78824, x73139);
  nand n78827(x78827, x68462, x78829);
  nand n78828(x78828, x78827, x73144);
  nand n78830(x78830, x68462, x78832);
  nand n78831(x78831, x78830, x73149);
  nand n78833(x78833, x68462, x78835);
  nand n78834(x78834, x78833, x73154);
  nand n78836(x78836, x68462, x78838);
  nand n78837(x78837, x78836, x73159);
  nand n78839(x78839, x68462, x78841);
  nand n78840(x78840, x78839, x73164);
  nand n78842(x78842, x68462, x78844);
  nand n78843(x78843, x78842, x73169);
  nand n78845(x78845, x68462, x78847);
  nand n78846(x78846, x78845, x73174);
  nand n78848(x78848, x68462, x78850);
  nand n78849(x78849, x78848, x73179);
  nand n78851(x78851, x68462, x78853);
  nand n78852(x78852, x78851, x73184);
  nand n78854(x78854, x68462, x78856);
  nand n78855(x78855, x78854, x73189);
  nand n78857(x78857, x68462, x78859);
  nand n78858(x78858, x78857, x73194);
  nand n78860(x78860, x68462, x78862);
  nand n78861(x78861, x78860, x73199);
  nand n78863(x78863, x68462, x78865);
  nand n78864(x78864, x78863, x73204);
  nand n78866(x78866, x68462, x78868);
  nand n78867(x78867, x78866, x73209);
  nand n78869(x78869, x68462, x78871);
  nand n78870(x78870, x78869, x73214);
  nand n78872(x78872, x68462, x78874);
  nand n78873(x78873, x78872, x73219);
  nand n78875(x78875, x68462, x78877);
  nand n78876(x78876, x78875, x73224);
  nand n78878(x78878, x68462, x78880);
  nand n78879(x78879, x78878, x73229);
  nand n78881(x78881, x68462, x78883);
  nand n78882(x78882, x78881, x73234);
  nand n78884(x78884, x68462, x78886);
  nand n78885(x78885, x78884, x73239);
  nand n78887(x78887, x68462, x78889);
  nand n78888(x78888, x78887, x73244);
  nand n78890(x78890, x68462, x78892);
  nand n78891(x78891, x78890, x73249);
  nand n78893(x78893, x68462, x78895);
  nand n78894(x78894, x78893, x73254);
  nand n78896(x78896, x68462, x78898);
  nand n78897(x78897, x78896, x73259);
  nand n78899(x78899, x68462, x78901);
  nand n78900(x78900, x78899, x73264);
  nand n78902(x78902, x68462, x78904);
  nand n78903(x78903, x78902, x73269);
  nand n78905(x78905, x68462, x78907);
  nand n78906(x78906, x78905, x73274);
  nand n78908(x78908, x68462, x78910);
  nand n78909(x78909, x78908, x73279);
  nand n78911(x78911, x68462, x78913);
  nand n78912(x78912, x78911, x73284);
  nand n78914(x78914, x68462, x78916);
  nand n78915(x78915, x78914, x73289);
  nand n78917(x78917, x68462, x78919);
  nand n78918(x78918, x78917, x73294);
  nand n78920(x78920, x68462, x78922);
  nand n78921(x78921, x78920, x73299);
  nand n78923(x78923, x68462, x78925);
  nand n78924(x78924, x78923, x73304);
  nand n78926(x78926, x68462, x78928);
  nand n78927(x78927, x78926, x73309);
  nand n78929(x78929, x68462, x78931);
  nand n78930(x78930, x78929, x73314);
  nand n78932(x78932, x68462, x78934);
  nand n78933(x78933, x78932, x73319);
  nand n78935(x78935, x68462, x78937);
  nand n78936(x78936, x78935, x73324);
  nand n78938(x78938, x68462, x78940);
  nand n78939(x78939, x78938, x73329);
  nand n78941(x78941, x68462, x78943);
  nand n78942(x78942, x78941, x73334);
  nand n78944(x78944, x68462, x78946);
  nand n78945(x78945, x78944, x73339);
  nand n78947(x78947, x68462, x78949);
  nand n78948(x78948, x78947, x73344);
  nand n78950(x78950, x68462, x78952);
  nand n78951(x78951, x78950, x73349);
  nand n78953(x78953, x68462, x78955);
  nand n78954(x78954, x78953, x73354);
  nand n78956(x78956, x68462, x78958);
  nand n78957(x78957, x78956, x73359);
  nand n78959(x78959, x68462, x78961);
  nand n78960(x78960, x78959, x73364);
  nand n78962(x78962, x68462, x78964);
  nand n78963(x78963, x78962, x73369);
  nand n78965(x78965, x68462, x78967);
  nand n78966(x78966, x78965, x73374);
  nand n78968(x78968, x68462, x78970);
  nand n78969(x78969, x78968, x73379);
  nand n78971(x78971, x68462, x78973);
  nand n78972(x78972, x78971, x73384);
  nand n78974(x78974, x68462, x78976);
  nand n78975(x78975, x78974, x73389);
  nand n78977(x78977, x68462, x78979);
  nand n78978(x78978, x78977, x73394);
  nand n78980(x78980, x68462, x78982);
  nand n78981(x78981, x78980, x73399);
  nand n78983(x78983, x68462, x78985);
  nand n78984(x78984, x78983, x73404);
  nand n78986(x78986, x68462, x78988);
  nand n78987(x78987, x78986, x73409);
  nand n78989(x78989, x68462, x78991);
  nand n78990(x78990, x78989, x73414);
  nand n78992(x78992, x68462, x78994);
  nand n78993(x78993, x78992, x73419);
  nand n78995(x78995, x68462, x78997);
  nand n78996(x78996, x78995, x73424);
  nand n78998(x78998, x68462, x79000);
  nand n78999(x78999, x78998, x73429);
  nand n79001(x79001, x68462, x79003);
  nand n79002(x79002, x79001, x73434);
  nand n79004(x79004, x68462, x79006);
  nand n79005(x79005, x79004, x73439);
  nand n79007(x79007, x68462, x79009);
  nand n79008(x79008, x79007, x73444);
  nand n79010(x79010, x68462, x79012);
  nand n79011(x79011, x79010, x73449);
  nand n79013(x79013, x68462, x79015);
  nand n79014(x79014, x79013, x73454);
  nand n79016(x79016, x68462, x79018);
  nand n79017(x79017, x79016, x73459);
  nand n79019(x79019, x68462, x79021);
  nand n79020(x79020, x79019, x73464);
  nand n79022(x79022, x68462, x79024);
  nand n79023(x79023, x79022, x73469);
  nand n79025(x79025, x68462, x79027);
  nand n79026(x79026, x79025, x73474);
  nand n79028(x79028, x68462, x79030);
  nand n79029(x79029, x79028, x73479);
  nand n79031(x79031, x68462, x79033);
  nand n79032(x79032, x79031, x73484);
  nand n79034(x79034, x68462, x79036);
  nand n79035(x79035, x79034, x73489);
  nand n79037(x79037, x68462, x79039);
  nand n79038(x79038, x79037, x73494);
  nand n79040(x79040, x68462, x79042);
  nand n79041(x79041, x79040, x73499);
  nand n79043(x79043, x68462, x79045);
  nand n79044(x79044, x79043, x73504);
  nand n79046(x79046, x68462, x79048);
  nand n79047(x79047, x79046, x73509);
  nand n79049(x79049, x68462, x79051);
  nand n79050(x79050, x79049, x73514);
  nand n79052(x79052, x68462, x79054);
  nand n79053(x79053, x79052, x73519);
  nand n79055(x79055, x68462, x79057);
  nand n79056(x79056, x79055, x73524);
  nand n79058(x79058, x68462, x79060);
  nand n79059(x79059, x79058, x73529);
  nand n79061(x79061, x68462, x79063);
  nand n79062(x79062, x79061, x73534);
  nand n79064(x79064, x68462, x79066);
  nand n79065(x79065, x79064, x73539);
  nand n79067(x79067, x68462, x79069);
  nand n79068(x79068, x79067, x73544);
  nand n79070(x79070, x68462, x79072);
  nand n79071(x79071, x79070, x73549);
  nand n79073(x79073, x68462, x79075);
  nand n79074(x79074, x79073, x73554);
  nand n79076(x79076, x68462, x79078);
  nand n79077(x79077, x79076, x73559);
  nand n79079(x79079, x68462, x79081);
  nand n79080(x79080, x79079, x73564);
  nand n79082(x79082, x68462, x79084);
  nand n79083(x79083, x79082, x73569);
  nand n79085(x79085, x68462, x79087);
  nand n79086(x79086, x79085, x73574);
  nand n79088(x79088, x68462, x79090);
  nand n79089(x79089, x79088, x73579);
  nand n79091(x79091, x68462, x79093);
  nand n79092(x79092, x79091, x73584);
  nand n79094(x79094, x68462, x79096);
  nand n79095(x79095, x79094, x73589);
  nand n79097(x79097, x68462, x79099);
  nand n79098(x79098, x79097, x73594);
  nand n79100(x79100, x68462, x79102);
  nand n79101(x79101, x79100, x73599);
  nand n79103(x79103, x68462, x79105);
  nand n79104(x79104, x79103, x73604);
  nand n79106(x79106, x68462, x79108);
  nand n79107(x79107, x79106, x73609);
  nand n79109(x79109, x68462, x79111);
  nand n79110(x79110, x79109, x73614);
  nand n79112(x79112, x68462, x79114);
  nand n79113(x79113, x79112, x73619);
  nand n79115(x79115, x68462, x79117);
  nand n79116(x79116, x79115, x73624);
  nand n79118(x79118, x68462, x79120);
  nand n79119(x79119, x79118, x73629);
  nand n79121(x79121, x68462, x79123);
  nand n79122(x79122, x79121, x73634);
  nand n79124(x79124, x68462, x79126);
  nand n79125(x79125, x79124, x73639);
  nand n79127(x79127, x68462, x79129);
  nand n79128(x79128, x79127, x73644);
  nand n79130(x79130, x68462, x79132);
  nand n79131(x79131, x79130, x73649);
  nand n79133(x79133, x68462, x79135);
  nand n79134(x79134, x79133, x73654);
  nand n79136(x79136, x68462, x79138);
  nand n79137(x79137, x79136, x73659);
  nand n79139(x79139, x68462, x79141);
  nand n79140(x79140, x79139, x73664);
  nand n79142(x79142, x68462, x79144);
  nand n79143(x79143, x79142, x73669);
  nand n79145(x79145, x68462, x79147);
  nand n79146(x79146, x79145, x73674);
  nand n79148(x79148, x68462, x79150);
  nand n79149(x79149, x79148, x73679);
  nand n79151(x79151, x68462, x79153);
  nand n79152(x79152, x79151, x73684);
  nand n79154(x79154, x68462, x79156);
  nand n79155(x79155, x79154, x73689);
  nand n79157(x79157, x68462, x79159);
  nand n79158(x79158, x79157, x73694);
  nand n79160(x79160, x68462, x79162);
  nand n79161(x79161, x79160, x73699);
  nand n79163(x79163, x68462, x79165);
  nand n79164(x79164, x79163, x73704);
  nand n79166(x79166, x68462, x79168);
  nand n79167(x79167, x79166, x73709);
  nand n79169(x79169, x68462, x79171);
  nand n79170(x79170, x79169, x73714);
  nand n79172(x79172, x68462, x79174);
  nand n79173(x79173, x79172, x73719);
  nand n79175(x79175, x68462, x79177);
  nand n79176(x79176, x79175, x73724);
  nand n79178(x79178, x68462, x79180);
  nand n79179(x79179, x79178, x73729);
  nand n79181(x79181, x68462, x79183);
  nand n79182(x79182, x79181, x73734);
  nand n79184(x79184, x68462, x79186);
  nand n79185(x79185, x79184, x73739);
  nand n79187(x79187, x68462, x79189);
  nand n79188(x79188, x79187, x73744);
  nand n79190(x79190, x68462, x79192);
  nand n79191(x79191, x79190, x73749);
  nand n79193(x79193, x68462, x79195);
  nand n79194(x79194, x79193, x73754);
  nand n79196(x79196, x68462, x79198);
  nand n79197(x79197, x79196, x73759);
  nand n79199(x79199, x68462, x79201);
  nand n79200(x79200, x79199, x73764);
  nand n79202(x79202, x68462, x79204);
  nand n79203(x79203, x79202, x73769);
  nand n79205(x79205, x68462, x79207);
  nand n79206(x79206, x79205, x73774);
  nand n79208(x79208, x68462, x79210);
  nand n79209(x79209, x79208, x73779);
  nand n79211(x79211, x68462, x79213);
  nand n79212(x79212, x79211, x73784);
  nand n79214(x79214, x68462, x79216);
  nand n79215(x79215, x79214, x73789);
  nand n79217(x79217, x68462, x79219);
  nand n79218(x79218, x79217, x73794);
  nand n79220(x79220, x68462, x79222);
  nand n79221(x79221, x79220, x73799);
  nand n79223(x79223, x68462, x79225);
  nand n79224(x79224, x79223, x73804);
  nand n79226(x79226, x68462, x79228);
  nand n79227(x79227, x79226, x73809);
  nand n79229(x79229, x68462, x79231);
  nand n79230(x79230, x79229, x73814);
  nand n79232(x79232, x68462, x79234);
  nand n79233(x79233, x79232, x73819);
  nand n79235(x79235, x68462, x79237);
  nand n79236(x79236, x79235, x73824);
  nand n79238(x79238, x68462, x79240);
  nand n79239(x79239, x79238, x73829);
  nand n79241(x79241, x68462, x79243);
  nand n79242(x79242, x79241, x73834);
  nand n79244(x79244, x68462, x79246);
  nand n79245(x79245, x79244, x73839);
  nand n79247(x79247, x68462, x79249);
  nand n79248(x79248, x79247, x73844);
  nand n79250(x79250, x68462, x79252);
  nand n79251(x79251, x79250, x73849);
  nand n79253(x79253, x68462, x79255);
  nand n79254(x79254, x79253, x73854);
  nand n79256(x79256, x68462, x79258);
  nand n79257(x79257, x79256, x73859);
  nand n79259(x79259, x68462, x79261);
  nand n79260(x79260, x79259, x73864);
  nand n79262(x79262, x68462, x79264);
  nand n79263(x79263, x79262, x73869);
  nand n79265(x79265, x68462, x79267);
  nand n79266(x79266, x79265, x73874);
  nand n79268(x79268, x68462, x79270);
  nand n79269(x79269, x79268, x73879);
  nand n79271(x79271, x68462, x79273);
  nand n79272(x79272, x79271, x73884);
  nand n79274(x79274, x68462, x79276);
  nand n79275(x79275, x79274, x73889);
  nand n79277(x79277, x68462, x79279);
  nand n79278(x79278, x79277, x73894);
  nand n79280(x79280, x68462, x79282);
  nand n79281(x79281, x79280, x73899);
  nand n79283(x79283, x68462, x79285);
  nand n79284(x79284, x79283, x73904);
  nand n79286(x79286, x68462, x79288);
  nand n79287(x79287, x79286, x73909);
  nand n79289(x79289, x68462, x79291);
  nand n79290(x79290, x79289, x73914);
  nand n79292(x79292, x68462, x79294);
  nand n79293(x79293, x79292, x73919);
  nand n79295(x79295, x68462, x79297);
  nand n79296(x79296, x79295, x73924);
  nand n79298(x79298, x68462, x79300);
  nand n79299(x79299, x79298, x73929);
  nand n79301(x79301, x68462, x79303);
  nand n79302(x79302, x79301, x73934);
  nand n79304(x79304, x68462, x79306);
  nand n79305(x79305, x79304, x73939);
  nand n79307(x79307, x68462, x79309);
  nand n79308(x79308, x79307, x73944);
  nand n79310(x79310, x68462, x79312);
  nand n79311(x79311, x79310, x73949);
  nand n79313(x79313, x68462, x79315);
  nand n79314(x79314, x79313, x73954);
  nand n79316(x79316, x68462, x79318);
  nand n79317(x79317, x79316, x73959);
  nand n79319(x79319, x68462, x79321);
  nand n79320(x79320, x79319, x73964);
  nand n79322(x79322, x68462, x79324);
  nand n79323(x79323, x79322, x73969);
  nand n79325(x79325, x68462, x79327);
  nand n79326(x79326, x79325, x73974);
  nand n79328(x79328, x68462, x79330);
  nand n79329(x79329, x79328, x73979);
  nand n79331(x79331, x68462, x79333);
  nand n79332(x79332, x79331, x73984);
  nand n79334(x79334, x68462, x79336);
  nand n79335(x79335, x79334, x73989);
  nand n79337(x79337, x68462, x79339);
  nand n79338(x79338, x79337, x73994);
  nand n79340(x79340, x68462, x79342);
  nand n79341(x79341, x79340, x73999);
  nand n79343(x79343, x68462, x79345);
  nand n79344(x79344, x79343, x71799);
  nand n79346(x79346, x68462, x79348);
  nand n79347(x79347, x79346, x71804);
  nand n79349(x79349, x68462, x79351);
  nand n79350(x79350, x79349, x71809);
  nand n79352(x79352, x68462, x79354);
  nand n79353(x79353, x79352, x71814);
  nand n79355(x79355, x68462, x79357);
  nand n79356(x79356, x79355, x71819);
  nand n79358(x79358, x68462, x79360);
  nand n79359(x79359, x79358, x71824);
  nand n79361(x79361, x68462, x79363);
  nand n79362(x79362, x79361, x71829);
  nand n79364(x79364, x68462, x79366);
  nand n79365(x79365, x79364, x71834);
  nand n79367(x79367, x68462, x79369);
  nand n79368(x79368, x79367, x71839);
  nand n79370(x79370, x68462, x79372);
  nand n79371(x79371, x79370, x71844);
  nand n79373(x79373, x68462, x79375);
  nand n79374(x79374, x79373, x71849);
  nand n79376(x79376, x68462, x79378);
  nand n79377(x79377, x79376, x71854);
  nand n79379(x79379, x68462, x79381);
  nand n79380(x79380, x79379, x71859);
  nand n79382(x79382, x68462, x79384);
  nand n79383(x79383, x79382, x71864);
  nand n79385(x79385, x68462, x79387);
  nand n79386(x79386, x79385, x71869);
  nand n79388(x79388, x68462, x79390);
  nand n79389(x79389, x79388, x71874);
  nand n79391(x79391, x68462, x79393);
  nand n79392(x79392, x79391, x71879);
  nand n79394(x79394, x68462, x79396);
  nand n79395(x79395, x79394, x71884);
  nand n79397(x79397, x68462, x79399);
  nand n79398(x79398, x79397, x71889);
  nand n79400(x79400, x68462, x79402);
  nand n79401(x79401, x79400, x71894);
  nand n79403(x79403, x68462, x79405);
  nand n79404(x79404, x79403, x71899);
  nand n79406(x79406, x68462, x79408);
  nand n79407(x79407, x79406, x71904);
  nand n79409(x79409, x68462, x79411);
  nand n79410(x79410, x79409, x71904);
  nand n79412(x79412, x68462, x79414);
  nand n79413(x79413, x79412, x71904);
  nand n79415(x79415, x68462, x79417);
  nand n79416(x79416, x79415, x71904);
  nand n79418(x79418, x68462, x79420);
  nand n79419(x79419, x79418, x71904);
  nand n79421(x79421, x68462, x79423);
  nand n79422(x79422, x79421, x71904);
  nand n79424(x79424, x68462, x79426);
  nand n79425(x79425, x79424, x71904);
  nand n79427(x79427, x68462, x79429);
  nand n79428(x79428, x79427, x71904);
  nand n79430(x79430, x68462, x79432);
  nand n79431(x79431, x79430, x71904);
  nand n79433(x79433, x68462, x79435);
  nand n79434(x79434, x79433, x71904);
  nand n79436(x79436, x68462, x79438);
  nand n79437(x79437, x79436, x71904);
  nand n79439(x79439, x68462, x79441);
  nand n79440(x79440, x79439, x71939);
  nand n79442(x79442, x68462, x79444);
  nand n79443(x79443, x79442, x71944);
  nand n79445(x79445, x68462, x79447);
  nand n79446(x79446, x79445, x71949);
  nand n79448(x79448, x68462, x79450);
  nand n79449(x79449, x79448, x71954);
  nand n79451(x79451, x68462, x79453);
  nand n79452(x79452, x79451, x71959);
  nand n79454(x79454, x68462, x79456);
  nand n79455(x79455, x79454, x71964);
  nand n79457(x79457, x68462, x79459);
  nand n79458(x79458, x79457, x71969);
  nand n79460(x79460, x68462, x79462);
  nand n79461(x79461, x79460, x71974);
  nand n79463(x79463, x68462, x79465);
  nand n79464(x79464, x79463, x71979);
  nand n79466(x79466, x68462, x79468);
  nand n79467(x79467, x79466, x71984);
  nand n79469(x79469, x68462, x79471);
  nand n79470(x79470, x79469, x71989);
  nand n79472(x79472, x68462, x79474);
  nand n79473(x79473, x79472, x71994);
  nand n79475(x79475, x68462, x79477);
  nand n79476(x79476, x79475, x71999);
  nand n79478(x79478, x68462, x79480);
  nand n79479(x79479, x79478, x72004);
  nand n79481(x79481, x68462, x79483);
  nand n79482(x79482, x79481, x72009);
  nand n79484(x79484, x68462, x79486);
  nand n79485(x79485, x79484, x72014);
  nand n79487(x79487, x68462, x79489);
  nand n79488(x79488, x79487, x72019);
  nand n79490(x79490, x68462, x79492);
  nand n79491(x79491, x79490, x72024);
  nand n79493(x79493, x68462, x79495);
  nand n79494(x79494, x79493, x72029);
  nand n79496(x79496, x68462, x79498);
  nand n79497(x79497, x79496, x72034);
  nand n79499(x79499, x68462, x79501);
  nand n79500(x79500, x79499, x72039);
  nand n79502(x79502, x68462, x79504);
  nand n79503(x79503, x79502, x72044);
  nand n79505(x79505, x68462, x79507);
  nand n79506(x79506, x79505, x72049);
  nand n79508(x79508, x68462, x79510);
  nand n79509(x79509, x79508, x72054);
  nand n79511(x79511, x68462, x79513);
  nand n79512(x79512, x79511, x72059);
  nand n79514(x79514, x68462, x79516);
  nand n79515(x79515, x79514, x72064);
  nand n79517(x79517, x68462, x79519);
  nand n79518(x79518, x79517, x72069);
  nand n79520(x79520, x68462, x79522);
  nand n79521(x79521, x79520, x72074);
  nand n79523(x79523, x68462, x79525);
  nand n79524(x79524, x79523, x72079);
  nand n79526(x79526, x68462, x79528);
  nand n79527(x79527, x79526, x72084);
  nand n79529(x79529, x68462, x79531);
  nand n79530(x79530, x79529, x72089);
  nand n79532(x79532, x68462, x79534);
  nand n79533(x79533, x79532, x72094);
  nand n79535(x79535, x68462, x79537);
  nand n79536(x79536, x79535, x72099);
  nand n79538(x79538, x68462, x79540);
  nand n79539(x79539, x79538, x72104);
  nand n79541(x79541, x68462, x79543);
  nand n79542(x79542, x79541, x72109);
  nand n79544(x79544, x68462, x79546);
  nand n79545(x79545, x79544, x72114);
  nand n79547(x79547, x68462, x79549);
  nand n79548(x79548, x79547, x72119);
  nand n79550(x79550, x68462, x79552);
  nand n79551(x79551, x79550, x72124);
  nand n79553(x79553, x68462, x79555);
  nand n79554(x79554, x79553, x72129);
  nand n79556(x79556, x68462, x79558);
  nand n79557(x79557, x79556, x72134);
  nand n79559(x79559, x68462, x79561);
  nand n79560(x79560, x79559, x72139);
  nand n79562(x79562, x68462, x79564);
  nand n79563(x79563, x79562, x72144);
  nand n79565(x79565, x68462, x79567);
  nand n79566(x79566, x79565, x72149);
  nand n79568(x79568, x68462, x79570);
  nand n79569(x79569, x79568, x72154);
  nand n79571(x79571, x68462, x79573);
  nand n79572(x79572, x79571, x72159);
  nand n79574(x79574, x68462, x79576);
  nand n79575(x79575, x79574, x72164);
  nand n79577(x79577, x68462, x79579);
  nand n79578(x79578, x79577, x72169);
  nand n79580(x79580, x68462, x79582);
  nand n79581(x79581, x79580, x72174);
  nand n79583(x79583, x68462, x79585);
  nand n79584(x79584, x79583, x72179);
  nand n79586(x79586, x68462, x79588);
  nand n79587(x79587, x79586, x72184);
  nand n79589(x79589, x68462, x79591);
  nand n79590(x79590, x79589, x72189);
  nand n79592(x79592, x68462, x79594);
  nand n79593(x79593, x79592, x72194);
  nand n79595(x79595, x68462, x79597);
  nand n79596(x79596, x79595, x72199);
  nand n79598(x79598, x68462, x79600);
  nand n79599(x79599, x79598, x72204);
  nand n79601(x79601, x68462, x79603);
  nand n79602(x79602, x79601, x72209);
  nand n79604(x79604, x68462, x79606);
  nand n79605(x79605, x79604, x72214);
  nand n79607(x79607, x68462, x79609);
  nand n79608(x79608, x79607, x72219);
  nand n79610(x79610, x68462, x79612);
  nand n79611(x79611, x79610, x72224);
  nand n79613(x79613, x68462, x79615);
  nand n79614(x79614, x79613, x72229);
  nand n79616(x79616, x68462, x79618);
  nand n79617(x79617, x79616, x72234);
  nand n79619(x79619, x68462, x79621);
  nand n79620(x79620, x79619, x72239);
  nand n79622(x79622, x68462, x79624);
  nand n79623(x79623, x79622, x72244);
  nand n79625(x79625, x68462, x79627);
  nand n79626(x79626, x79625, x72249);
  nand n79628(x79628, x68462, x79630);
  nand n79629(x79629, x79628, x72254);
  nand n79631(x79631, x68462, x79633);
  nand n79632(x79632, x79631, x72259);
  nand n79634(x79634, x68462, x79636);
  nand n79635(x79635, x79634, x72264);
  nand n79637(x79637, x68462, x79639);
  nand n79638(x79638, x79637, x72269);
  nand n79640(x79640, x68462, x79642);
  nand n79641(x79641, x79640, x72274);
  nand n79643(x79643, x68462, x79645);
  nand n79644(x79644, x79643, x72279);
  nand n79646(x79646, x68462, x79648);
  nand n79647(x79647, x79646, x72284);
  nand n79649(x79649, x68462, x79651);
  nand n79650(x79650, x79649, x72289);
  nand n79652(x79652, x68462, x79654);
  nand n79653(x79653, x79652, x72294);
  nand n79655(x79655, x68462, x79657);
  nand n79656(x79656, x79655, x72299);
  nand n79658(x79658, x68462, x79660);
  nand n79659(x79659, x79658, x72304);
  nand n79661(x79661, x68462, x79663);
  nand n79662(x79662, x79661, x72309);
  nand n79664(x79664, x68462, x79666);
  nand n79665(x79665, x79664, x72314);
  nand n79667(x79667, x68462, x79669);
  nand n79668(x79668, x79667, x72319);
  nand n79670(x79670, x68462, x79672);
  nand n79671(x79671, x79670, x72324);
  nand n79673(x79673, x68462, x79675);
  nand n79674(x79674, x79673, x72329);
  nand n79676(x79676, x68462, x79678);
  nand n79677(x79677, x79676, x72334);
  nand n79679(x79679, x68462, x79681);
  nand n79680(x79680, x79679, x72339);
  nand n79682(x79682, x68462, x79684);
  nand n79683(x79683, x79682, x72344);
  nand n79685(x79685, x68462, x79687);
  nand n79686(x79686, x79685, x72349);
  nand n79688(x79688, x68462, x79690);
  nand n79689(x79689, x79688, x72354);
  nand n79691(x79691, x68462, x79693);
  nand n79692(x79692, x79691, x72359);
  nand n79694(x79694, x68462, x79696);
  nand n79695(x79695, x79694, x72364);
  nand n79697(x79697, x68462, x79699);
  nand n79698(x79698, x79697, x72369);
  nand n79700(x79700, x68462, x79702);
  nand n79701(x79701, x79700, x72374);
  nand n79703(x79703, x68462, x79705);
  nand n79704(x79704, x79703, x72379);
  nand n79706(x79706, x68462, x79708);
  nand n79707(x79707, x79706, x72384);
  nand n79709(x79709, x68462, x79711);
  nand n79710(x79710, x79709, x72389);
  nand n79712(x79712, x68462, x79714);
  nand n79713(x79713, x79712, x72394);
  nand n79715(x79715, x68462, x79717);
  nand n79716(x79716, x79715, x72399);
  nand n79718(x79718, x68462, x79720);
  nand n79719(x79719, x79718, x72404);
  nand n79721(x79721, x68462, x79723);
  nand n79722(x79722, x79721, x72409);
  nand n79724(x79724, x68462, x79726);
  nand n79725(x79725, x79724, x72414);
  nand n79727(x79727, x68462, x79729);
  nand n79728(x79728, x79727, x72419);
  nand n79730(x79730, x68462, x79732);
  nand n79731(x79731, x79730, x72424);
  nand n79733(x79733, x68462, x79735);
  nand n79734(x79734, x79733, x72429);
  nand n79736(x79736, x68462, x79738);
  nand n79737(x79737, x79736, x72434);
  nand n79739(x79739, x68462, x79741);
  nand n79740(x79740, x79739, x72439);
  nand n79742(x79742, x68462, x79744);
  nand n79743(x79743, x79742, x72444);
  nand n79745(x79745, x68462, x79747);
  nand n79746(x79746, x79745, x72449);
  nand n79748(x79748, x68462, x79750);
  nand n79749(x79749, x79748, x72454);
  nand n79751(x79751, x68462, x79753);
  nand n79752(x79752, x79751, x72459);
  nand n79754(x79754, x68462, x79756);
  nand n79755(x79755, x79754, x72464);
  nand n79757(x79757, x68462, x79759);
  nand n79758(x79758, x79757, x72469);
  nand n79760(x79760, x68462, x79762);
  nand n79761(x79761, x79760, x72474);
  nand n79763(x79763, x68462, x79765);
  nand n79764(x79764, x79763, x72479);
  nand n79766(x79766, x68462, x79768);
  nand n79767(x79767, x79766, x72484);
  nand n79769(x79769, x68462, x79771);
  nand n79770(x79770, x79769, x72489);
  nand n79772(x79772, x68462, x79774);
  nand n79773(x79773, x79772, x72494);
  nand n79775(x79775, x68462, x79777);
  nand n79776(x79776, x79775, x72499);
  nand n79778(x79778, x68462, x79780);
  nand n79779(x79779, x79778, x72504);
  nand n79781(x79781, x68462, x79783);
  nand n79782(x79782, x79781, x72509);
  nand n79784(x79784, x68462, x79786);
  nand n79785(x79785, x79784, x72514);
  nand n79787(x79787, x68462, x79789);
  nand n79788(x79788, x79787, x72519);
  nand n79790(x79790, x68462, x79792);
  nand n79791(x79791, x79790, x72524);
  nand n79793(x79793, x68462, x79795);
  nand n79794(x79794, x79793, x72529);
  nand n79796(x79796, x68462, x79798);
  nand n79797(x79797, x79796, x72534);
  nand n79799(x79799, x68462, x79801);
  nand n79800(x79800, x79799, x72539);
  nand n79802(x79802, x68462, x79804);
  nand n79803(x79803, x79802, x72544);
  nand n79805(x79805, x68462, x79807);
  nand n79806(x79806, x79805, x72549);
  nand n79808(x79808, x68462, x79810);
  nand n79809(x79809, x79808, x72554);
  nand n79811(x79811, x68462, x79813);
  nand n79812(x79812, x79811, x72559);
  nand n79814(x79814, x68462, x79816);
  nand n79815(x79815, x79814, x72564);
  nand n79817(x79817, x68462, x79819);
  nand n79818(x79818, x79817, x72569);
  nand n79820(x79820, x68462, x79822);
  nand n79821(x79821, x79820, x72574);
  nand n79823(x79823, x68462, x79825);
  nand n79824(x79824, x79823, x72579);
  nand n79826(x79826, x68462, x79828);
  nand n79827(x79827, x79826, x72584);
  nand n79829(x79829, x68462, x79831);
  nand n79830(x79830, x79829, x72589);
  nand n79832(x79832, x68462, x79834);
  nand n79833(x79833, x79832, x72594);
  nand n79835(x79835, x68462, x79837);
  nand n79836(x79836, x79835, x72599);
  nand n79838(x79838, x68462, x79840);
  nand n79839(x79839, x79838, x72604);
  nand n79841(x79841, x68462, x79843);
  nand n79842(x79842, x79841, x72609);
  nand n79844(x79844, x68462, x79846);
  nand n79845(x79845, x79844, x72614);
  nand n79847(x79847, x68462, x79849);
  nand n79848(x79848, x79847, x72619);
  nand n79850(x79850, x68462, x79852);
  nand n79851(x79851, x79850, x72624);
  nand n79853(x79853, x68462, x79855);
  nand n79854(x79854, x79853, x72629);
  nand n79856(x79856, x68462, x79858);
  nand n79857(x79857, x79856, x72634);
  nand n79859(x79859, x68462, x79861);
  nand n79860(x79860, x79859, x72639);
  nand n79862(x79862, x68462, x79864);
  nand n79863(x79863, x79862, x72644);
  nand n79865(x79865, x68462, x79867);
  nand n79866(x79866, x79865, x72649);
  nand n79868(x79868, x68462, x79870);
  nand n79869(x79869, x79868, x72654);
  nand n79871(x79871, x68462, x79873);
  nand n79872(x79872, x79871, x72659);
  nand n79874(x79874, x68462, x79876);
  nand n79875(x79875, x79874, x72664);
  nand n79877(x79877, x68462, x79879);
  nand n79878(x79878, x79877, x72669);
  nand n79880(x79880, x68462, x79882);
  nand n79881(x79881, x79880, x72674);
  nand n79883(x79883, x68462, x79885);
  nand n79884(x79884, x79883, x72679);
  nand n79886(x79886, x68462, x79888);
  nand n79887(x79887, x79886, x72684);
  nand n79889(x79889, x68462, x79891);
  nand n79890(x79890, x79889, x72689);
  nand n79892(x79892, x68462, x79894);
  nand n79893(x79893, x79892, x72694);
  nand n79895(x79895, x68462, x79897);
  nand n79896(x79896, x79895, x72699);
  nand n79898(x79898, x68462, x79900);
  nand n79899(x79899, x79898, x72704);
  nand n79901(x79901, x68462, x79903);
  nand n79902(x79902, x79901, x72709);
  nand n79904(x79904, x68462, x79906);
  nand n79905(x79905, x79904, x72714);
  nand n79907(x79907, x68462, x79909);
  nand n79908(x79908, x79907, x72719);
  nand n79910(x79910, x68462, x79912);
  nand n79911(x79911, x79910, x72724);
  nand n79913(x79913, x68462, x79915);
  nand n79914(x79914, x79913, x72729);
  nand n79916(x79916, x68462, x79918);
  nand n79917(x79917, x79916, x72734);
  nand n79919(x79919, x68462, x79921);
  nand n79920(x79920, x79919, x72739);
  nand n79922(x79922, x68462, x79924);
  nand n79923(x79923, x79922, x72744);
  nand n79925(x79925, x68462, x79927);
  nand n79926(x79926, x79925, x72749);
  nand n79928(x79928, x68462, x79930);
  nand n79929(x79929, x79928, x72754);
  nand n79931(x79931, x68462, x79933);
  nand n79932(x79932, x79931, x72759);
  nand n79934(x79934, x68462, x79936);
  nand n79935(x79935, x79934, x72764);
  nand n79937(x79937, x68462, x79939);
  nand n79938(x79938, x79937, x72769);
  nand n79940(x79940, x68462, x79942);
  nand n79941(x79941, x79940, x72774);
  nand n79943(x79943, x68462, x79945);
  nand n79944(x79944, x79943, x72779);
  nand n79946(x79946, x68462, x79948);
  nand n79947(x79947, x79946, x72784);
  nand n79949(x79949, x68462, x79951);
  nand n79950(x79950, x79949, x72789);
  nand n79952(x79952, x68462, x79954);
  nand n79953(x79953, x79952, x72794);
  nand n79955(x79955, x68462, x79957);
  nand n79956(x79956, x79955, x72799);
  nand n79958(x79958, x68462, x79960);
  nand n79959(x79959, x79958, x72804);
  nand n79961(x79961, x68462, x79963);
  nand n79962(x79962, x79961, x72809);
  nand n79964(x79964, x68462, x79966);
  nand n79965(x79965, x79964, x72814);
  nand n79967(x79967, x68462, x79969);
  nand n79968(x79968, x79967, x72819);
  nand n79970(x79970, x68462, x79972);
  nand n79971(x79971, x79970, x72824);
  nand n79973(x79973, x68462, x79975);
  nand n79974(x79974, x79973, x72829);
  nand n79976(x79976, x68462, x79978);
  nand n79977(x79977, x79976, x72834);
  nand n79979(x79979, x68462, x79981);
  nand n79980(x79980, x79979, x72839);
  nand n79982(x79982, x68462, x79984);
  nand n79983(x79983, x79982, x72844);
  nand n79985(x79985, x68462, x79987);
  nand n79986(x79986, x79985, x72849);
  nand n79988(x79988, x68462, x79990);
  nand n79989(x79989, x79988, x72854);
  nand n79991(x79991, x68462, x79993);
  nand n79992(x79992, x79991, x72859);
  nand n79994(x79994, x68462, x79996);
  nand n79995(x79995, x79994, x72864);
  nand n79997(x79997, x68462, x79999);
  nand n79998(x79998, x79997, x72869);
  nand n80000(x80000, x68462, x80002);
  nand n80001(x80001, x80000, x72874);
  nand n80003(x80003, x68462, x80005);
  nand n80004(x80004, x80003, x72879);
  nand n80006(x80006, x68462, x80008);
  nand n80007(x80007, x80006, x72884);
  nand n80009(x80009, x68462, x80011);
  nand n80010(x80010, x80009, x72889);
  nand n80012(x80012, x68462, x80014);
  nand n80013(x80013, x80012, x72894);
  nand n80015(x80015, x68462, x80017);
  nand n80016(x80016, x80015, x72899);
  nand n80018(x80018, x68462, x80020);
  nand n80019(x80019, x80018, x72904);
  nand n80021(x80021, x68462, x80023);
  nand n80022(x80022, x80021, x72909);
  nand n80024(x80024, x68462, x80026);
  nand n80025(x80025, x80024, x72914);
  nand n80027(x80027, x68462, x80029);
  nand n80028(x80028, x80027, x72919);
  nand n80030(x80030, x68462, x80032);
  nand n80031(x80031, x80030, x72924);
  nand n80033(x80033, x68462, x80035);
  nand n80034(x80034, x80033, x72929);
  nand n80036(x80036, x68462, x80038);
  nand n80037(x80037, x80036, x72934);
  nand n80039(x80039, x68462, x80041);
  nand n80040(x80040, x80039, x72939);
  nand n80042(x80042, x68462, x80044);
  nand n80043(x80043, x80042, x72944);
  nand n80045(x80045, x68462, x80047);
  nand n80046(x80046, x80045, x72949);
  nand n80048(x80048, x68462, x80050);
  nand n80049(x80049, x80048, x72954);
  nand n80051(x80051, x68462, x80053);
  nand n80052(x80052, x80051, x72959);
  nand n80054(x80054, x68462, x80056);
  nand n80055(x80055, x80054, x72964);
  nand n80057(x80057, x68462, x80059);
  nand n80058(x80058, x80057, x72969);
  nand n80060(x80060, x68462, x80062);
  nand n80061(x80061, x80060, x72974);
  nand n80063(x80063, x68462, x80065);
  nand n80064(x80064, x80063, x72979);
  nand n80066(x80066, x68462, x80068);
  nand n80067(x80067, x80066, x72984);
  nand n80069(x80069, x68462, x80071);
  nand n80070(x80070, x80069, x72989);
  nand n80072(x80072, x68462, x80074);
  nand n80073(x80073, x80072, x72994);
  nand n80075(x80075, x68462, x80077);
  nand n80076(x80076, x80075, x72999);
  nand n80078(x80078, x68462, x80080);
  nand n80079(x80079, x80078, x73004);
  nand n80081(x80081, x68462, x80083);
  nand n80082(x80082, x80081, x73009);
  nand n80084(x80084, x68462, x80086);
  nand n80085(x80085, x80084, x73014);
  nand n80087(x80087, x68462, x80089);
  nand n80088(x80088, x80087, x73019);
  nand n80090(x80090, x68462, x80092);
  nand n80091(x80091, x80090, x73024);
  nand n80093(x80093, x68462, x80095);
  nand n80094(x80094, x80093, x73029);
  nand n80096(x80096, x68462, x80098);
  nand n80097(x80097, x80096, x73034);
  nand n80099(x80099, x68462, x80101);
  nand n80100(x80100, x80099, x73039);
  nand n80102(x80102, x68462, x80104);
  nand n80103(x80103, x80102, x73044);
  nand n80105(x80105, x68462, x80107);
  nand n80106(x80106, x80105, x73049);
  nand n80108(x80108, x68462, x80110);
  nand n80109(x80109, x80108, x73054);
  nand n80111(x80111, x68462, x80113);
  nand n80112(x80112, x80111, x73059);
  nand n80114(x80114, x68462, x80116);
  nand n80115(x80115, x80114, x73064);
  nand n80117(x80117, x68462, x80119);
  nand n80118(x80118, x80117, x73069);
  nand n80120(x80120, x68462, x80122);
  nand n80121(x80121, x80120, x73074);
  nand n80123(x80123, x68462, x80125);
  nand n80124(x80124, x80123, x73079);
  nand n80126(x80126, x68462, x80128);
  nand n80127(x80127, x80126, x73084);
  nand n80129(x80129, x68462, x80131);
  nand n80130(x80130, x80129, x73089);
  nand n80132(x80132, x68462, x80134);
  nand n80133(x80133, x80132, x73094);
  nand n80135(x80135, x68462, x80137);
  nand n80136(x80136, x80135, x73099);
  nand n80138(x80138, x68462, x80140);
  nand n80139(x80139, x80138, x73104);
  nand n80141(x80141, x68462, x80143);
  nand n80142(x80142, x80141, x73109);
  nand n80144(x80144, x68462, x80146);
  nand n80145(x80145, x80144, x73114);
  nand n80147(x80147, x68462, x80149);
  nand n80148(x80148, x80147, x73119);
  nand n80150(x80150, x68462, x80152);
  nand n80151(x80151, x80150, x73124);
  nand n80153(x80153, x68462, x80155);
  nand n80154(x80154, x80153, x73129);
  nand n80156(x80156, x68462, x80158);
  nand n80157(x80157, x80156, x73134);
  nand n80159(x80159, x68462, x80161);
  nand n80160(x80160, x80159, x73139);
  nand n80162(x80162, x68462, x80164);
  nand n80163(x80163, x80162, x73144);
  nand n80165(x80165, x68462, x80167);
  nand n80166(x80166, x80165, x73149);
  nand n80168(x80168, x68462, x80170);
  nand n80169(x80169, x80168, x73154);
  nand n80171(x80171, x68462, x80173);
  nand n80172(x80172, x80171, x73159);
  nand n80174(x80174, x68462, x80176);
  nand n80175(x80175, x80174, x73164);
  nand n80177(x80177, x68462, x80179);
  nand n80178(x80178, x80177, x73169);
  nand n80180(x80180, x68462, x80182);
  nand n80181(x80181, x80180, x73174);
  nand n80183(x80183, x68462, x80185);
  nand n80184(x80184, x80183, x73179);
  nand n80186(x80186, x68462, x80188);
  nand n80187(x80187, x80186, x73184);
  nand n80189(x80189, x68462, x80191);
  nand n80190(x80190, x80189, x73189);
  nand n80192(x80192, x68462, x80194);
  nand n80193(x80193, x80192, x73194);
  nand n80195(x80195, x68462, x80197);
  nand n80196(x80196, x80195, x73199);
  nand n80198(x80198, x68462, x80200);
  nand n80199(x80199, x80198, x73204);
  nand n80201(x80201, x68462, x80203);
  nand n80202(x80202, x80201, x73209);
  nand n80204(x80204, x68462, x80206);
  nand n80205(x80205, x80204, x73214);
  nand n80207(x80207, x68462, x80209);
  nand n80208(x80208, x80207, x73219);
  nand n80210(x80210, x68462, x80212);
  nand n80211(x80211, x80210, x73224);
  nand n80213(x80213, x68462, x80215);
  nand n80214(x80214, x80213, x73229);
  nand n80216(x80216, x68462, x80218);
  nand n80217(x80217, x80216, x73234);
  nand n80219(x80219, x68462, x80221);
  nand n80220(x80220, x80219, x73239);
  nand n80222(x80222, x68462, x80224);
  nand n80223(x80223, x80222, x73244);
  nand n80225(x80225, x68462, x80227);
  nand n80226(x80226, x80225, x73249);
  nand n80228(x80228, x68462, x80230);
  nand n80229(x80229, x80228, x73254);
  nand n80231(x80231, x68462, x80233);
  nand n80232(x80232, x80231, x73259);
  nand n80234(x80234, x68462, x80236);
  nand n80235(x80235, x80234, x73264);
  nand n80237(x80237, x68462, x80239);
  nand n80238(x80238, x80237, x73269);
  nand n80240(x80240, x68462, x80242);
  nand n80241(x80241, x80240, x73274);
  nand n80243(x80243, x68462, x80245);
  nand n80244(x80244, x80243, x73279);
  nand n80246(x80246, x68462, x80248);
  nand n80247(x80247, x80246, x73284);
  nand n80249(x80249, x68462, x80251);
  nand n80250(x80250, x80249, x73289);
  nand n80252(x80252, x68462, x80254);
  nand n80253(x80253, x80252, x73294);
  nand n80255(x80255, x68462, x80257);
  nand n80256(x80256, x80255, x73299);
  nand n80258(x80258, x68462, x80260);
  nand n80259(x80259, x80258, x73304);
  nand n80261(x80261, x68462, x80263);
  nand n80262(x80262, x80261, x73309);
  nand n80264(x80264, x68462, x80266);
  nand n80265(x80265, x80264, x73314);
  nand n80267(x80267, x68462, x80269);
  nand n80268(x80268, x80267, x73319);
  nand n80270(x80270, x68462, x80272);
  nand n80271(x80271, x80270, x73324);
  nand n80273(x80273, x68462, x80275);
  nand n80274(x80274, x80273, x73329);
  nand n80276(x80276, x68462, x80278);
  nand n80277(x80277, x80276, x73334);
  nand n80279(x80279, x68462, x80281);
  nand n80280(x80280, x80279, x73339);
  nand n80282(x80282, x68462, x80284);
  nand n80283(x80283, x80282, x73344);
  nand n80285(x80285, x68462, x80287);
  nand n80286(x80286, x80285, x73349);
  nand n80288(x80288, x68462, x80290);
  nand n80289(x80289, x80288, x73354);
  nand n80291(x80291, x68462, x80293);
  nand n80292(x80292, x80291, x73359);
  nand n80294(x80294, x68462, x80296);
  nand n80295(x80295, x80294, x73364);
  nand n80297(x80297, x68462, x80299);
  nand n80298(x80298, x80297, x73369);
  nand n80300(x80300, x68462, x80302);
  nand n80301(x80301, x80300, x73374);
  nand n80303(x80303, x68462, x80305);
  nand n80304(x80304, x80303, x73379);
  nand n80306(x80306, x68462, x80308);
  nand n80307(x80307, x80306, x73384);
  nand n80309(x80309, x68462, x80311);
  nand n80310(x80310, x80309, x73389);
  nand n80312(x80312, x68462, x80314);
  nand n80313(x80313, x80312, x73394);
  nand n80315(x80315, x68462, x80317);
  nand n80316(x80316, x80315, x73399);
  nand n80318(x80318, x68462, x80320);
  nand n80319(x80319, x80318, x73404);
  nand n80321(x80321, x68462, x80323);
  nand n80322(x80322, x80321, x73409);
  nand n80324(x80324, x68462, x80326);
  nand n80325(x80325, x80324, x73414);
  nand n80327(x80327, x68462, x80329);
  nand n80328(x80328, x80327, x73419);
  nand n80330(x80330, x68462, x80332);
  nand n80331(x80331, x80330, x73424);
  nand n80333(x80333, x68462, x80335);
  nand n80334(x80334, x80333, x73429);
  nand n80336(x80336, x68462, x80338);
  nand n80337(x80337, x80336, x73434);
  nand n80339(x80339, x68462, x80341);
  nand n80340(x80340, x80339, x73439);
  nand n80342(x80342, x68462, x80344);
  nand n80343(x80343, x80342, x73444);
  nand n80345(x80345, x68462, x80347);
  nand n80346(x80346, x80345, x73449);
  nand n80348(x80348, x68462, x80350);
  nand n80349(x80349, x80348, x73454);
  nand n80351(x80351, x68462, x80353);
  nand n80352(x80352, x80351, x73459);
  nand n80354(x80354, x68462, x80356);
  nand n80355(x80355, x80354, x73464);
  nand n80357(x80357, x68462, x80359);
  nand n80358(x80358, x80357, x73469);
  nand n80360(x80360, x68462, x80362);
  nand n80361(x80361, x80360, x73474);
  nand n80363(x80363, x68462, x80365);
  nand n80364(x80364, x80363, x73479);
  nand n80366(x80366, x68462, x80368);
  nand n80367(x80367, x80366, x73484);
  nand n80369(x80369, x68462, x80371);
  nand n80370(x80370, x80369, x73489);
  nand n80372(x80372, x68462, x80374);
  nand n80373(x80373, x80372, x73494);
  nand n80375(x80375, x68462, x80377);
  nand n80376(x80376, x80375, x73499);
  nand n80378(x80378, x68462, x80380);
  nand n80379(x80379, x80378, x73504);
  nand n80381(x80381, x68462, x80383);
  nand n80382(x80382, x80381, x73509);
  nand n80384(x80384, x68462, x80386);
  nand n80385(x80385, x80384, x73514);
  nand n80387(x80387, x68462, x80389);
  nand n80388(x80388, x80387, x73519);
  nand n80390(x80390, x68462, x80392);
  nand n80391(x80391, x80390, x73524);
  nand n80393(x80393, x68462, x80395);
  nand n80394(x80394, x80393, x73529);
  nand n80396(x80396, x68462, x80398);
  nand n80397(x80397, x80396, x73534);
  nand n80399(x80399, x68462, x80401);
  nand n80400(x80400, x80399, x73539);
  nand n80402(x80402, x68462, x80404);
  nand n80403(x80403, x80402, x73544);
  nand n80405(x80405, x68462, x80407);
  nand n80406(x80406, x80405, x73549);
  nand n80408(x80408, x68462, x80410);
  nand n80409(x80409, x80408, x73554);
  nand n80411(x80411, x68462, x80413);
  nand n80412(x80412, x80411, x73559);
  nand n80414(x80414, x68462, x80416);
  nand n80415(x80415, x80414, x73564);
  nand n80417(x80417, x68462, x80419);
  nand n80418(x80418, x80417, x73569);
  nand n80420(x80420, x68462, x80422);
  nand n80421(x80421, x80420, x73574);
  nand n80423(x80423, x68462, x80425);
  nand n80424(x80424, x80423, x73579);
  nand n80426(x80426, x68462, x80428);
  nand n80427(x80427, x80426, x73584);
  nand n80429(x80429, x68462, x80431);
  nand n80430(x80430, x80429, x73589);
  nand n80432(x80432, x68462, x80434);
  nand n80433(x80433, x80432, x73594);
  nand n80435(x80435, x68462, x80437);
  nand n80436(x80436, x80435, x73599);
  nand n80438(x80438, x68462, x80440);
  nand n80439(x80439, x80438, x73604);
  nand n80441(x80441, x68462, x80443);
  nand n80442(x80442, x80441, x73609);
  nand n80444(x80444, x68462, x80446);
  nand n80445(x80445, x80444, x73614);
  nand n80447(x80447, x68462, x80449);
  nand n80448(x80448, x80447, x73619);
  nand n80450(x80450, x68462, x80452);
  nand n80451(x80451, x80450, x73624);
  nand n80453(x80453, x68462, x80455);
  nand n80454(x80454, x80453, x73629);
  nand n80456(x80456, x68462, x80458);
  nand n80457(x80457, x80456, x73634);
  nand n80459(x80459, x68462, x80461);
  nand n80460(x80460, x80459, x73639);
  nand n80462(x80462, x68462, x80464);
  nand n80463(x80463, x80462, x73644);
  nand n80465(x80465, x68462, x80467);
  nand n80466(x80466, x80465, x73649);
  nand n80468(x80468, x68462, x80470);
  nand n80469(x80469, x80468, x73654);
  nand n80471(x80471, x68462, x80473);
  nand n80472(x80472, x80471, x73659);
  nand n80474(x80474, x68462, x80476);
  nand n80475(x80475, x80474, x73664);
  nand n80477(x80477, x68462, x80479);
  nand n80478(x80478, x80477, x73669);
  nand n80480(x80480, x68462, x80482);
  nand n80481(x80481, x80480, x73674);
  nand n80483(x80483, x68462, x80485);
  nand n80484(x80484, x80483, x73679);
  nand n80486(x80486, x68462, x80488);
  nand n80487(x80487, x80486, x73684);
  nand n80489(x80489, x68462, x80491);
  nand n80490(x80490, x80489, x73689);
  nand n80492(x80492, x68462, x80494);
  nand n80493(x80493, x80492, x73694);
  nand n80495(x80495, x68462, x80497);
  nand n80496(x80496, x80495, x73699);
  nand n80498(x80498, x68462, x80500);
  nand n80499(x80499, x80498, x73704);
  nand n80501(x80501, x68462, x80503);
  nand n80502(x80502, x80501, x73709);
  nand n80504(x80504, x68462, x80506);
  nand n80505(x80505, x80504, x73714);
  nand n80507(x80507, x68462, x80509);
  nand n80508(x80508, x80507, x73719);
  nand n80510(x80510, x68462, x80512);
  nand n80511(x80511, x80510, x73724);
  nand n80513(x80513, x68462, x80515);
  nand n80514(x80514, x80513, x73729);
  nand n80516(x80516, x68462, x80518);
  nand n80517(x80517, x80516, x73734);
  nand n80519(x80519, x68462, x80521);
  nand n80520(x80520, x80519, x73739);
  nand n80522(x80522, x68462, x80524);
  nand n80523(x80523, x80522, x73744);
  nand n80525(x80525, x68462, x80527);
  nand n80526(x80526, x80525, x73749);
  nand n80528(x80528, x68462, x80530);
  nand n80529(x80529, x80528, x73754);
  nand n80531(x80531, x68462, x80533);
  nand n80532(x80532, x80531, x73759);
  nand n80534(x80534, x68462, x80536);
  nand n80535(x80535, x80534, x73764);
  nand n80537(x80537, x68462, x80539);
  nand n80538(x80538, x80537, x73769);
  nand n80540(x80540, x68462, x80542);
  nand n80541(x80541, x80540, x73774);
  nand n80543(x80543, x68462, x80545);
  nand n80544(x80544, x80543, x73779);
  nand n80546(x80546, x68462, x80548);
  nand n80547(x80547, x80546, x73784);
  nand n80549(x80549, x68462, x80551);
  nand n80550(x80550, x80549, x73789);
  nand n80552(x80552, x68462, x80554);
  nand n80553(x80553, x80552, x73794);
  nand n80555(x80555, x68462, x80557);
  nand n80556(x80556, x80555, x73799);
  nand n80558(x80558, x68462, x80560);
  nand n80559(x80559, x80558, x73804);
  nand n80561(x80561, x68462, x80563);
  nand n80562(x80562, x80561, x73809);
  nand n80564(x80564, x68462, x80566);
  nand n80565(x80565, x80564, x73814);
  nand n80567(x80567, x68462, x80569);
  nand n80568(x80568, x80567, x73819);
  nand n80570(x80570, x68462, x80572);
  nand n80571(x80571, x80570, x73824);
  nand n80573(x80573, x68462, x80575);
  nand n80574(x80574, x80573, x73829);
  nand n80576(x80576, x68462, x80578);
  nand n80577(x80577, x80576, x73834);
  nand n80579(x80579, x68462, x80581);
  nand n80580(x80580, x80579, x73839);
  nand n80582(x80582, x68462, x80584);
  nand n80583(x80583, x80582, x73844);
  nand n80585(x80585, x68462, x80587);
  nand n80586(x80586, x80585, x73849);
  nand n80588(x80588, x68462, x80590);
  nand n80589(x80589, x80588, x73854);
  nand n80591(x80591, x68462, x80593);
  nand n80592(x80592, x80591, x73859);
  nand n80594(x80594, x68462, x80596);
  nand n80595(x80595, x80594, x73864);
  nand n80597(x80597, x68462, x80599);
  nand n80598(x80598, x80597, x73869);
  nand n80600(x80600, x68462, x80602);
  nand n80601(x80601, x80600, x73874);
  nand n80603(x80603, x68462, x80605);
  nand n80604(x80604, x80603, x73879);
  nand n80606(x80606, x68462, x80608);
  nand n80607(x80607, x80606, x73884);
  nand n80609(x80609, x68462, x80611);
  nand n80610(x80610, x80609, x73889);
  nand n80612(x80612, x68462, x80614);
  nand n80613(x80613, x80612, x73894);
  nand n80615(x80615, x68462, x80617);
  nand n80616(x80616, x80615, x73899);
  nand n80618(x80618, x68462, x80620);
  nand n80619(x80619, x80618, x73904);
  nand n80621(x80621, x68462, x80623);
  nand n80622(x80622, x80621, x73909);
  nand n80624(x80624, x68462, x80626);
  nand n80625(x80625, x80624, x73914);
  nand n80627(x80627, x68462, x80629);
  nand n80628(x80628, x80627, x73919);
  nand n80630(x80630, x68462, x80632);
  nand n80631(x80631, x80630, x73924);
  nand n80633(x80633, x68462, x80635);
  nand n80634(x80634, x80633, x73929);
  nand n80636(x80636, x68462, x80638);
  nand n80637(x80637, x80636, x73934);
  nand n80639(x80639, x68462, x80641);
  nand n80640(x80640, x80639, x73939);
  nand n80642(x80642, x68462, x80644);
  nand n80643(x80643, x80642, x73944);
  nand n80645(x80645, x68462, x80647);
  nand n80646(x80646, x80645, x73949);
  nand n80648(x80648, x68462, x80650);
  nand n80649(x80649, x80648, x73954);
  nand n80651(x80651, x68462, x80653);
  nand n80652(x80652, x80651, x73959);
  nand n80654(x80654, x68462, x80656);
  nand n80655(x80655, x80654, x73964);
  nand n80657(x80657, x68462, x80659);
  nand n80658(x80658, x80657, x73969);
  nand n80660(x80660, x68462, x80662);
  nand n80661(x80661, x80660, x73974);
  nand n80663(x80663, x68462, x80665);
  nand n80664(x80664, x80663, x73979);
  nand n80666(x80666, x68462, x80668);
  nand n80667(x80667, x80666, x73984);
  nand n80669(x80669, x68462, x80671);
  nand n80670(x80670, x80669, x73989);
  nand n80672(x80672, x68462, x80674);
  nand n80673(x80673, x80672, x73994);
  nand n80675(x80675, x68462, x80677);
  nand n80676(x80676, x80675, x73999);
  nand n80678(x80678, x68462, x80680);
  nand n80679(x80679, x80678, x71799);
  nand n80681(x80681, x68462, x80683);
  nand n80682(x80682, x80681, x71804);
  nand n80684(x80684, x68462, x80686);
  nand n80685(x80685, x80684, x71809);
  nand n80687(x80687, x68462, x80689);
  nand n80688(x80688, x80687, x71814);
  nand n80690(x80690, x68462, x80692);
  nand n80691(x80691, x80690, x71819);
  nand n80693(x80693, x68462, x80695);
  nand n80694(x80694, x80693, x71824);
  nand n80696(x80696, x68462, x80698);
  nand n80697(x80697, x80696, x71829);
  nand n80699(x80699, x68462, x80701);
  nand n80700(x80700, x80699, x71834);
  nand n80702(x80702, x68462, x80704);
  nand n80703(x80703, x80702, x71839);
  nand n80705(x80705, x68462, x80707);
  nand n80706(x80706, x80705, x71844);
  nand n80708(x80708, x68462, x80710);
  nand n80709(x80709, x80708, x71849);
  nand n80711(x80711, x68462, x80713);
  nand n80712(x80712, x80711, x71854);
  nand n80714(x80714, x68462, x80716);
  nand n80715(x80715, x80714, x71859);
  nand n80717(x80717, x68462, x80719);
  nand n80718(x80718, x80717, x71864);
  nand n80720(x80720, x68462, x80722);
  nand n80721(x80721, x80720, x71869);
  nand n80723(x80723, x68462, x80725);
  nand n80724(x80724, x80723, x71874);
  nand n80726(x80726, x68462, x80728);
  nand n80727(x80727, x80726, x71879);
  nand n80729(x80729, x68462, x80731);
  nand n80730(x80730, x80729, x71884);
  nand n80732(x80732, x68462, x80734);
  nand n80733(x80733, x80732, x71889);
  nand n80735(x80735, x68462, x80737);
  nand n80736(x80736, x80735, x71894);
  nand n80738(x80738, x68462, x80740);
  nand n80739(x80739, x80738, x71899);
  nand n80741(x80741, x68462, x80743);
  nand n80742(x80742, x80741, x71904);
  nand n80744(x80744, x68462, x80746);
  nand n80745(x80745, x80744, x71904);
  nand n80747(x80747, x68462, x80749);
  nand n80748(x80748, x80747, x71904);
  nand n80750(x80750, x68462, x80752);
  nand n80751(x80751, x80750, x71904);
  nand n80753(x80753, x68462, x80755);
  nand n80754(x80754, x80753, x71904);
  nand n80756(x80756, x68462, x80758);
  nand n80757(x80757, x80756, x71904);
  nand n80759(x80759, x68462, x80761);
  nand n80760(x80760, x80759, x71904);
  nand n80762(x80762, x68462, x80764);
  nand n80763(x80763, x80762, x71904);
  nand n80765(x80765, x68462, x80767);
  nand n80766(x80766, x80765, x71904);
  nand n80768(x80768, x68462, x80770);
  nand n80769(x80769, x80768, x71904);
  nand n80771(x80771, x68462, x80773);
  nand n80772(x80772, x80771, x71904);
  nand n80774(x80774, x68462, x80776);
  nand n80775(x80775, x80774, x71939);
  nand n80777(x80777, x68462, x80779);
  nand n80778(x80778, x80777, x71944);
  nand n80780(x80780, x68462, x80782);
  nand n80781(x80781, x80780, x71949);
  nand n80783(x80783, x68462, x80785);
  nand n80784(x80784, x80783, x71954);
  nand n80786(x80786, x68462, x80788);
  nand n80787(x80787, x80786, x71959);
  nand n80789(x80789, x68462, x80791);
  nand n80790(x80790, x80789, x71964);
  nand n80792(x80792, x68462, x80794);
  nand n80793(x80793, x80792, x71969);
  nand n80795(x80795, x68462, x80797);
  nand n80796(x80796, x80795, x71974);
  nand n80798(x80798, x68462, x80800);
  nand n80799(x80799, x80798, x71979);
  nand n80801(x80801, x68462, x80803);
  nand n80802(x80802, x80801, x71984);
  nand n80804(x80804, x68462, x80806);
  nand n80805(x80805, x80804, x71989);
  nand n80807(x80807, x68462, x80809);
  nand n80808(x80808, x80807, x71994);
  nand n80810(x80810, x68462, x80812);
  nand n80811(x80811, x80810, x71999);
  nand n80813(x80813, x68462, x80815);
  nand n80814(x80814, x80813, x72004);
  nand n80816(x80816, x68462, x80818);
  nand n80817(x80817, x80816, x72009);
  nand n80819(x80819, x68462, x80821);
  nand n80820(x80820, x80819, x72014);
  nand n80822(x80822, x68462, x80824);
  nand n80823(x80823, x80822, x72019);
  nand n80825(x80825, x68462, x80827);
  nand n80826(x80826, x80825, x72024);
  nand n80828(x80828, x68462, x80830);
  nand n80829(x80829, x80828, x72029);
  nand n80831(x80831, x68462, x80833);
  nand n80832(x80832, x80831, x72034);
  nand n80834(x80834, x68462, x80836);
  nand n80835(x80835, x80834, x72039);
  nand n80837(x80837, x68462, x80839);
  nand n80838(x80838, x80837, x72044);
  nand n80840(x80840, x68462, x80842);
  nand n80841(x80841, x80840, x72049);
  nand n80843(x80843, x68462, x80845);
  nand n80844(x80844, x80843, x72054);
  nand n80846(x80846, x68462, x80848);
  nand n80847(x80847, x80846, x72059);
  nand n80849(x80849, x68462, x80851);
  nand n80850(x80850, x80849, x72064);
  nand n80852(x80852, x68462, x80854);
  nand n80853(x80853, x80852, x72069);
  nand n80855(x80855, x68462, x80857);
  nand n80856(x80856, x80855, x72074);
  nand n80858(x80858, x68462, x80860);
  nand n80859(x80859, x80858, x72079);
  nand n80861(x80861, x68462, x80863);
  nand n80862(x80862, x80861, x72084);
  nand n80864(x80864, x68462, x80866);
  nand n80865(x80865, x80864, x72089);
  nand n80867(x80867, x68462, x80869);
  nand n80868(x80868, x80867, x72094);
  nand n80870(x80870, x68462, x80872);
  nand n80871(x80871, x80870, x72099);
  nand n80873(x80873, x68462, x80875);
  nand n80874(x80874, x80873, x72104);
  nand n80876(x80876, x68462, x80878);
  nand n80877(x80877, x80876, x72109);
  nand n80879(x80879, x68462, x80881);
  nand n80880(x80880, x80879, x72114);
  nand n80882(x80882, x68462, x80884);
  nand n80883(x80883, x80882, x72119);
  nand n80885(x80885, x68462, x80887);
  nand n80886(x80886, x80885, x72124);
  nand n80888(x80888, x68462, x80890);
  nand n80889(x80889, x80888, x72129);
  nand n80891(x80891, x68462, x80893);
  nand n80892(x80892, x80891, x72134);
  nand n80894(x80894, x68462, x80896);
  nand n80895(x80895, x80894, x72139);
  nand n80897(x80897, x68462, x80899);
  nand n80898(x80898, x80897, x72144);
  nand n80900(x80900, x68462, x80902);
  nand n80901(x80901, x80900, x72149);
  nand n80903(x80903, x68462, x80905);
  nand n80904(x80904, x80903, x72154);
  nand n80906(x80906, x68462, x80908);
  nand n80907(x80907, x80906, x72159);
  nand n80909(x80909, x68462, x80911);
  nand n80910(x80910, x80909, x72164);
  nand n80912(x80912, x68462, x80914);
  nand n80913(x80913, x80912, x72169);
  nand n80915(x80915, x68462, x80917);
  nand n80916(x80916, x80915, x72174);
  nand n80918(x80918, x68462, x80920);
  nand n80919(x80919, x80918, x72179);
  nand n80921(x80921, x68462, x80923);
  nand n80922(x80922, x80921, x72184);
  nand n80924(x80924, x68462, x80926);
  nand n80925(x80925, x80924, x72189);
  nand n80927(x80927, x68462, x80929);
  nand n80928(x80928, x80927, x72194);
  nand n80930(x80930, x68462, x80932);
  nand n80931(x80931, x80930, x72199);
  nand n80933(x80933, x68462, x80935);
  nand n80934(x80934, x80933, x72204);
  nand n80936(x80936, x68462, x80938);
  nand n80937(x80937, x80936, x72209);
  nand n80939(x80939, x68462, x80941);
  nand n80940(x80940, x80939, x72214);
  nand n80942(x80942, x68462, x80944);
  nand n80943(x80943, x80942, x72219);
  nand n80945(x80945, x68462, x80947);
  nand n80946(x80946, x80945, x72224);
  nand n80948(x80948, x68462, x80950);
  nand n80949(x80949, x80948, x72229);
  nand n80951(x80951, x68462, x80953);
  nand n80952(x80952, x80951, x72234);
  nand n80954(x80954, x68462, x80956);
  nand n80955(x80955, x80954, x72239);
  nand n80957(x80957, x68462, x80959);
  nand n80958(x80958, x80957, x72244);
  nand n80960(x80960, x68462, x80962);
  nand n80961(x80961, x80960, x72249);
  nand n80963(x80963, x68462, x80965);
  nand n80964(x80964, x80963, x72254);
  nand n80966(x80966, x68462, x80968);
  nand n80967(x80967, x80966, x72259);
  nand n80969(x80969, x68462, x80971);
  nand n80970(x80970, x80969, x72264);
  nand n80972(x80972, x68462, x80974);
  nand n80973(x80973, x80972, x72269);
  nand n80975(x80975, x68462, x80977);
  nand n80976(x80976, x80975, x72274);
  nand n80978(x80978, x68462, x80980);
  nand n80979(x80979, x80978, x72279);
  nand n80981(x80981, x68462, x80983);
  nand n80982(x80982, x80981, x72284);
  nand n80984(x80984, x68462, x80986);
  nand n80985(x80985, x80984, x72289);
  nand n80987(x80987, x68462, x80989);
  nand n80988(x80988, x80987, x72294);
  nand n80990(x80990, x68462, x80992);
  nand n80991(x80991, x80990, x72299);
  nand n80993(x80993, x68462, x80995);
  nand n80994(x80994, x80993, x72304);
  nand n80996(x80996, x68462, x80998);
  nand n80997(x80997, x80996, x72309);
  nand n80999(x80999, x68462, x81001);
  nand n81000(x81000, x80999, x72314);
  nand n81002(x81002, x68462, x81004);
  nand n81003(x81003, x81002, x72319);
  nand n81005(x81005, x68462, x81007);
  nand n81006(x81006, x81005, x72324);
  nand n81008(x81008, x68462, x81010);
  nand n81009(x81009, x81008, x72329);
  nand n81011(x81011, x68462, x81013);
  nand n81012(x81012, x81011, x72334);
  nand n81014(x81014, x68462, x81016);
  nand n81015(x81015, x81014, x72339);
  nand n81017(x81017, x68462, x81019);
  nand n81018(x81018, x81017, x72344);
  nand n81020(x81020, x68462, x81022);
  nand n81021(x81021, x81020, x72349);
  nand n81023(x81023, x68462, x81025);
  nand n81024(x81024, x81023, x72354);
  nand n81026(x81026, x68462, x81028);
  nand n81027(x81027, x81026, x72359);
  nand n81029(x81029, x68462, x81031);
  nand n81030(x81030, x81029, x72364);
  nand n81032(x81032, x68462, x81034);
  nand n81033(x81033, x81032, x72369);
  nand n81035(x81035, x68462, x81037);
  nand n81036(x81036, x81035, x72374);
  nand n81038(x81038, x68462, x81040);
  nand n81039(x81039, x81038, x72379);
  nand n81041(x81041, x68462, x81043);
  nand n81042(x81042, x81041, x72384);
  nand n81044(x81044, x68462, x81046);
  nand n81045(x81045, x81044, x72389);
  nand n81047(x81047, x68462, x81049);
  nand n81048(x81048, x81047, x72394);
  nand n81050(x81050, x68462, x81052);
  nand n81051(x81051, x81050, x72399);
  nand n81053(x81053, x68462, x81055);
  nand n81054(x81054, x81053, x72404);
  nand n81056(x81056, x68462, x81058);
  nand n81057(x81057, x81056, x72409);
  nand n81059(x81059, x68462, x81061);
  nand n81060(x81060, x81059, x72414);
  nand n81062(x81062, x68462, x81064);
  nand n81063(x81063, x81062, x72419);
  nand n81065(x81065, x68462, x81067);
  nand n81066(x81066, x81065, x72424);
  nand n81068(x81068, x68462, x81070);
  nand n81069(x81069, x81068, x72429);
  nand n81071(x81071, x68462, x81073);
  nand n81072(x81072, x81071, x72434);
  nand n81074(x81074, x68462, x81076);
  nand n81075(x81075, x81074, x72439);
  nand n81077(x81077, x68462, x81079);
  nand n81078(x81078, x81077, x72444);
  nand n81080(x81080, x68462, x81082);
  nand n81081(x81081, x81080, x72449);
  nand n81083(x81083, x68462, x81085);
  nand n81084(x81084, x81083, x72454);
  nand n81086(x81086, x68462, x81088);
  nand n81087(x81087, x81086, x72459);
  nand n81089(x81089, x68462, x81091);
  nand n81090(x81090, x81089, x72464);
  nand n81092(x81092, x68462, x81094);
  nand n81093(x81093, x81092, x72469);
  nand n81095(x81095, x68462, x81097);
  nand n81096(x81096, x81095, x72474);
  nand n81098(x81098, x68462, x81100);
  nand n81099(x81099, x81098, x72479);
  nand n81101(x81101, x68462, x81103);
  nand n81102(x81102, x81101, x72484);
  nand n81104(x81104, x68462, x81106);
  nand n81105(x81105, x81104, x72489);
  nand n81107(x81107, x68462, x81109);
  nand n81108(x81108, x81107, x72494);
  nand n81110(x81110, x68462, x81112);
  nand n81111(x81111, x81110, x72499);
  nand n81113(x81113, x68462, x81115);
  nand n81114(x81114, x81113, x72504);
  nand n81116(x81116, x68462, x81118);
  nand n81117(x81117, x81116, x72509);
  nand n81119(x81119, x68462, x81121);
  nand n81120(x81120, x81119, x72514);
  nand n81122(x81122, x68462, x81124);
  nand n81123(x81123, x81122, x72519);
  nand n81125(x81125, x68462, x81127);
  nand n81126(x81126, x81125, x72524);
  nand n81128(x81128, x68462, x81130);
  nand n81129(x81129, x81128, x72529);
  nand n81131(x81131, x68462, x81133);
  nand n81132(x81132, x81131, x72534);
  nand n81134(x81134, x68462, x81136);
  nand n81135(x81135, x81134, x72539);
  nand n81137(x81137, x68462, x81139);
  nand n81138(x81138, x81137, x72544);
  nand n81140(x81140, x68462, x81142);
  nand n81141(x81141, x81140, x72549);
  nand n81143(x81143, x68462, x81145);
  nand n81144(x81144, x81143, x72554);
  nand n81146(x81146, x68462, x81148);
  nand n81147(x81147, x81146, x72559);
  nand n81149(x81149, x68462, x81151);
  nand n81150(x81150, x81149, x72564);
  nand n81152(x81152, x68462, x81154);
  nand n81153(x81153, x81152, x72569);
  nand n81155(x81155, x68462, x81157);
  nand n81156(x81156, x81155, x72574);
  nand n81158(x81158, x68462, x81160);
  nand n81159(x81159, x81158, x72579);
  nand n81161(x81161, x68462, x81163);
  nand n81162(x81162, x81161, x72584);
  nand n81164(x81164, x68462, x81166);
  nand n81165(x81165, x81164, x72589);
  nand n81167(x81167, x68462, x81169);
  nand n81168(x81168, x81167, x72594);
  nand n81170(x81170, x68462, x81172);
  nand n81171(x81171, x81170, x72599);
  nand n81173(x81173, x68462, x81175);
  nand n81174(x81174, x81173, x72604);
  nand n81176(x81176, x68462, x81178);
  nand n81177(x81177, x81176, x72609);
  nand n81179(x81179, x68462, x81181);
  nand n81180(x81180, x81179, x72614);
  nand n81182(x81182, x68462, x81184);
  nand n81183(x81183, x81182, x72619);
  nand n81185(x81185, x68462, x81187);
  nand n81186(x81186, x81185, x72624);
  nand n81188(x81188, x68462, x81190);
  nand n81189(x81189, x81188, x72629);
  nand n81191(x81191, x68462, x81193);
  nand n81192(x81192, x81191, x72634);
  nand n81194(x81194, x68462, x81196);
  nand n81195(x81195, x81194, x72639);
  nand n81197(x81197, x68462, x81199);
  nand n81198(x81198, x81197, x72644);
  nand n81200(x81200, x68462, x81202);
  nand n81201(x81201, x81200, x72649);
  nand n81203(x81203, x68462, x81205);
  nand n81204(x81204, x81203, x72654);
  nand n81206(x81206, x68462, x81208);
  nand n81207(x81207, x81206, x72659);
  nand n81209(x81209, x68462, x81211);
  nand n81210(x81210, x81209, x72664);
  nand n81212(x81212, x68462, x81214);
  nand n81213(x81213, x81212, x72669);
  nand n81215(x81215, x68462, x81217);
  nand n81216(x81216, x81215, x72674);
  nand n81218(x81218, x68462, x81220);
  nand n81219(x81219, x81218, x72679);
  nand n81221(x81221, x68462, x81223);
  nand n81222(x81222, x81221, x72684);
  nand n81224(x81224, x68462, x81226);
  nand n81225(x81225, x81224, x72689);
  nand n81227(x81227, x68462, x81229);
  nand n81228(x81228, x81227, x72694);
  nand n81230(x81230, x68462, x81232);
  nand n81231(x81231, x81230, x72699);
  nand n81233(x81233, x68462, x81235);
  nand n81234(x81234, x81233, x72704);
  nand n81236(x81236, x68462, x81238);
  nand n81237(x81237, x81236, x72709);
  nand n81239(x81239, x68462, x81241);
  nand n81240(x81240, x81239, x72714);
  nand n81242(x81242, x68462, x81244);
  nand n81243(x81243, x81242, x72719);
  nand n81245(x81245, x68462, x81247);
  nand n81246(x81246, x81245, x72724);
  nand n81248(x81248, x68462, x81250);
  nand n81249(x81249, x81248, x72729);
  nand n81251(x81251, x68462, x81253);
  nand n81252(x81252, x81251, x72734);
  nand n81254(x81254, x68462, x81256);
  nand n81255(x81255, x81254, x72739);
  nand n81257(x81257, x68462, x81259);
  nand n81258(x81258, x81257, x72744);
  nand n81260(x81260, x68462, x81262);
  nand n81261(x81261, x81260, x72749);
  nand n81263(x81263, x68462, x81265);
  nand n81264(x81264, x81263, x72754);
  nand n81266(x81266, x68462, x81268);
  nand n81267(x81267, x81266, x72759);
  nand n81269(x81269, x68462, x81271);
  nand n81270(x81270, x81269, x72764);
  nand n81272(x81272, x68462, x81274);
  nand n81273(x81273, x81272, x72769);
  nand n81275(x81275, x68462, x81277);
  nand n81276(x81276, x81275, x72774);
  nand n81278(x81278, x68462, x81280);
  nand n81279(x81279, x81278, x72779);
  nand n81281(x81281, x68462, x81283);
  nand n81282(x81282, x81281, x72784);
  nand n81284(x81284, x68462, x81286);
  nand n81285(x81285, x81284, x72789);
  nand n81287(x81287, x68462, x81289);
  nand n81288(x81288, x81287, x72794);
  nand n81290(x81290, x68462, x81292);
  nand n81291(x81291, x81290, x72799);
  nand n81293(x81293, x68462, x81295);
  nand n81294(x81294, x81293, x72804);
  nand n81296(x81296, x68462, x81298);
  nand n81297(x81297, x81296, x72809);
  nand n81299(x81299, x68462, x81301);
  nand n81300(x81300, x81299, x72814);
  nand n81302(x81302, x68462, x81304);
  nand n81303(x81303, x81302, x72819);
  nand n81305(x81305, x68462, x81307);
  nand n81306(x81306, x81305, x72824);
  nand n81308(x81308, x68462, x81310);
  nand n81309(x81309, x81308, x72829);
  nand n81311(x81311, x68462, x81313);
  nand n81312(x81312, x81311, x72834);
  nand n81314(x81314, x68462, x81316);
  nand n81315(x81315, x81314, x72839);
  nand n81317(x81317, x68462, x81319);
  nand n81318(x81318, x81317, x72844);
  nand n81320(x81320, x68462, x81322);
  nand n81321(x81321, x81320, x72849);
  nand n81323(x81323, x68462, x81325);
  nand n81324(x81324, x81323, x72854);
  nand n81326(x81326, x68462, x81328);
  nand n81327(x81327, x81326, x72859);
  nand n81329(x81329, x68462, x81331);
  nand n81330(x81330, x81329, x72864);
  nand n81332(x81332, x68462, x81334);
  nand n81333(x81333, x81332, x72869);
  nand n81335(x81335, x68462, x81337);
  nand n81336(x81336, x81335, x72874);
  nand n81338(x81338, x68462, x81340);
  nand n81339(x81339, x81338, x72879);
  nand n81341(x81341, x68462, x81343);
  nand n81342(x81342, x81341, x72884);
  nand n81344(x81344, x68462, x81346);
  nand n81345(x81345, x81344, x72889);
  nand n81347(x81347, x68462, x81349);
  nand n81348(x81348, x81347, x72894);
  nand n81350(x81350, x68462, x81352);
  nand n81351(x81351, x81350, x72899);
  nand n81353(x81353, x68462, x81355);
  nand n81354(x81354, x81353, x72904);
  nand n81356(x81356, x68462, x81358);
  nand n81357(x81357, x81356, x72909);
  nand n81359(x81359, x68462, x81361);
  nand n81360(x81360, x81359, x72914);
  nand n81362(x81362, x68462, x81364);
  nand n81363(x81363, x81362, x72919);
  nand n81365(x81365, x68462, x81367);
  nand n81366(x81366, x81365, x72924);
  nand n81368(x81368, x68462, x81370);
  nand n81369(x81369, x81368, x72929);
  nand n81371(x81371, x68462, x81373);
  nand n81372(x81372, x81371, x72934);
  nand n81374(x81374, x68462, x81376);
  nand n81375(x81375, x81374, x72939);
  nand n81377(x81377, x68462, x81379);
  nand n81378(x81378, x81377, x72944);
  nand n81380(x81380, x68462, x81382);
  nand n81381(x81381, x81380, x72949);
  nand n81383(x81383, x68462, x81385);
  nand n81384(x81384, x81383, x72954);
  nand n81386(x81386, x68462, x81388);
  nand n81387(x81387, x81386, x72959);
  nand n81389(x81389, x68462, x81391);
  nand n81390(x81390, x81389, x72964);
  nand n81392(x81392, x68462, x81394);
  nand n81393(x81393, x81392, x72969);
  nand n81395(x81395, x68462, x81397);
  nand n81396(x81396, x81395, x72974);
  nand n81398(x81398, x68462, x81400);
  nand n81399(x81399, x81398, x72979);
  nand n81401(x81401, x68462, x81403);
  nand n81402(x81402, x81401, x72984);
  nand n81404(x81404, x68462, x81406);
  nand n81405(x81405, x81404, x72989);
  nand n81407(x81407, x68462, x81409);
  nand n81408(x81408, x81407, x72994);
  nand n81410(x81410, x68462, x81412);
  nand n81411(x81411, x81410, x72999);
  nand n81413(x81413, x68462, x81415);
  nand n81414(x81414, x81413, x73004);
  nand n81416(x81416, x68462, x81418);
  nand n81417(x81417, x81416, x73009);
  nand n81419(x81419, x68462, x81421);
  nand n81420(x81420, x81419, x73014);
  nand n81422(x81422, x68462, x81424);
  nand n81423(x81423, x81422, x73019);
  nand n81425(x81425, x68462, x81427);
  nand n81426(x81426, x81425, x73024);
  nand n81428(x81428, x68462, x81430);
  nand n81429(x81429, x81428, x73029);
  nand n81431(x81431, x68462, x81433);
  nand n81432(x81432, x81431, x73034);
  nand n81434(x81434, x68462, x81436);
  nand n81435(x81435, x81434, x73039);
  nand n81437(x81437, x68462, x81439);
  nand n81438(x81438, x81437, x73044);
  nand n81440(x81440, x68462, x81442);
  nand n81441(x81441, x81440, x73049);
  nand n81443(x81443, x68462, x81445);
  nand n81444(x81444, x81443, x73054);
  nand n81446(x81446, x68462, x81448);
  nand n81447(x81447, x81446, x73059);
  nand n81449(x81449, x68462, x81451);
  nand n81450(x81450, x81449, x73064);
  nand n81452(x81452, x68462, x81454);
  nand n81453(x81453, x81452, x73069);
  nand n81455(x81455, x68462, x81457);
  nand n81456(x81456, x81455, x73074);
  nand n81458(x81458, x68462, x81460);
  nand n81459(x81459, x81458, x73079);
  nand n81461(x81461, x68462, x81463);
  nand n81462(x81462, x81461, x73084);
  nand n81464(x81464, x68462, x81466);
  nand n81465(x81465, x81464, x73089);
  nand n81467(x81467, x68462, x81469);
  nand n81468(x81468, x81467, x73094);
  nand n81470(x81470, x68462, x81472);
  nand n81471(x81471, x81470, x73099);
  nand n81473(x81473, x68462, x81475);
  nand n81474(x81474, x81473, x73104);
  nand n81476(x81476, x68462, x81478);
  nand n81477(x81477, x81476, x73109);
  nand n81479(x81479, x68462, x81481);
  nand n81480(x81480, x81479, x73114);
  nand n81482(x81482, x68462, x81484);
  nand n81483(x81483, x81482, x73119);
  nand n81485(x81485, x68462, x81487);
  nand n81486(x81486, x81485, x73124);
  nand n81488(x81488, x68462, x81490);
  nand n81489(x81489, x81488, x73129);
  nand n81491(x81491, x68462, x81493);
  nand n81492(x81492, x81491, x73134);
  nand n81494(x81494, x68462, x81496);
  nand n81495(x81495, x81494, x73139);
  nand n81497(x81497, x68462, x81499);
  nand n81498(x81498, x81497, x73144);
  nand n81500(x81500, x68462, x81502);
  nand n81501(x81501, x81500, x73149);
  nand n81503(x81503, x68462, x81505);
  nand n81504(x81504, x81503, x73154);
  nand n81506(x81506, x68462, x81508);
  nand n81507(x81507, x81506, x73159);
  nand n81509(x81509, x68462, x81511);
  nand n81510(x81510, x81509, x73164);
  nand n81512(x81512, x68462, x81514);
  nand n81513(x81513, x81512, x73169);
  nand n81515(x81515, x68462, x81517);
  nand n81516(x81516, x81515, x73174);
  nand n81518(x81518, x68462, x81520);
  nand n81519(x81519, x81518, x73179);
  nand n81521(x81521, x68462, x81523);
  nand n81522(x81522, x81521, x73184);
  nand n81524(x81524, x68462, x81526);
  nand n81525(x81525, x81524, x73189);
  nand n81527(x81527, x68462, x81529);
  nand n81528(x81528, x81527, x73194);
  nand n81530(x81530, x68462, x81532);
  nand n81531(x81531, x81530, x73199);
  nand n81533(x81533, x68462, x81535);
  nand n81534(x81534, x81533, x73204);
  nand n81536(x81536, x68462, x81538);
  nand n81537(x81537, x81536, x73209);
  nand n81539(x81539, x68462, x81541);
  nand n81540(x81540, x81539, x73214);
  nand n81542(x81542, x68462, x81544);
  nand n81543(x81543, x81542, x73219);
  nand n81545(x81545, x68462, x81547);
  nand n81546(x81546, x81545, x73224);
  nand n81548(x81548, x68462, x81550);
  nand n81549(x81549, x81548, x73229);
  nand n81551(x81551, x68462, x81553);
  nand n81552(x81552, x81551, x73234);
  nand n81554(x81554, x68462, x81556);
  nand n81555(x81555, x81554, x73239);
  nand n81557(x81557, x68462, x81559);
  nand n81558(x81558, x81557, x73244);
  nand n81560(x81560, x68462, x81562);
  nand n81561(x81561, x81560, x73249);
  nand n81563(x81563, x68462, x81565);
  nand n81564(x81564, x81563, x73254);
  nand n81566(x81566, x68462, x81568);
  nand n81567(x81567, x81566, x73259);
  nand n81569(x81569, x68462, x81571);
  nand n81570(x81570, x81569, x73264);
  nand n81572(x81572, x68462, x81574);
  nand n81573(x81573, x81572, x73269);
  nand n81575(x81575, x68462, x81577);
  nand n81576(x81576, x81575, x73274);
  nand n81578(x81578, x68462, x81580);
  nand n81579(x81579, x81578, x73279);
  nand n81581(x81581, x68462, x81583);
  nand n81582(x81582, x81581, x73284);
  nand n81584(x81584, x68462, x81586);
  nand n81585(x81585, x81584, x73289);
  nand n81587(x81587, x68462, x81589);
  nand n81588(x81588, x81587, x73294);
  nand n81590(x81590, x68462, x81592);
  nand n81591(x81591, x81590, x73299);
  nand n81593(x81593, x68462, x81595);
  nand n81594(x81594, x81593, x73304);
  nand n81596(x81596, x68462, x81598);
  nand n81597(x81597, x81596, x73309);
  nand n81599(x81599, x68462, x81601);
  nand n81600(x81600, x81599, x73314);
  nand n81602(x81602, x68462, x81604);
  nand n81603(x81603, x81602, x73319);
  nand n81605(x81605, x68462, x81607);
  nand n81606(x81606, x81605, x73324);
  nand n81608(x81608, x68462, x81610);
  nand n81609(x81609, x81608, x73329);
  nand n81611(x81611, x68462, x81613);
  nand n81612(x81612, x81611, x73334);
  nand n81614(x81614, x68462, x81616);
  nand n81615(x81615, x81614, x73339);
  nand n81617(x81617, x68462, x81619);
  nand n81618(x81618, x81617, x73344);
  nand n81620(x81620, x68462, x81622);
  nand n81621(x81621, x81620, x73349);
  nand n81623(x81623, x68462, x81625);
  nand n81624(x81624, x81623, x73354);
  nand n81626(x81626, x68462, x81628);
  nand n81627(x81627, x81626, x73359);
  nand n81629(x81629, x68462, x81631);
  nand n81630(x81630, x81629, x73364);
  nand n81632(x81632, x68462, x81634);
  nand n81633(x81633, x81632, x73369);
  nand n81635(x81635, x68462, x81637);
  nand n81636(x81636, x81635, x73374);
  nand n81638(x81638, x68462, x81640);
  nand n81639(x81639, x81638, x73379);
  nand n81641(x81641, x68462, x81643);
  nand n81642(x81642, x81641, x73384);
  nand n81644(x81644, x68462, x81646);
  nand n81645(x81645, x81644, x73389);
  nand n81647(x81647, x68462, x81649);
  nand n81648(x81648, x81647, x73394);
  nand n81650(x81650, x68462, x81652);
  nand n81651(x81651, x81650, x73399);
  nand n81653(x81653, x68462, x81655);
  nand n81654(x81654, x81653, x73404);
  nand n81656(x81656, x68462, x81658);
  nand n81657(x81657, x81656, x73409);
  nand n81659(x81659, x68462, x81661);
  nand n81660(x81660, x81659, x73414);
  nand n81662(x81662, x68462, x81664);
  nand n81663(x81663, x81662, x73419);
  nand n81665(x81665, x68462, x81667);
  nand n81666(x81666, x81665, x73424);
  nand n81668(x81668, x68462, x81670);
  nand n81669(x81669, x81668, x73429);
  nand n81671(x81671, x68462, x81673);
  nand n81672(x81672, x81671, x73434);
  nand n81674(x81674, x68462, x81676);
  nand n81675(x81675, x81674, x73439);
  nand n81677(x81677, x68462, x81679);
  nand n81678(x81678, x81677, x73444);
  nand n81680(x81680, x68462, x81682);
  nand n81681(x81681, x81680, x73449);
  nand n81683(x81683, x68462, x81685);
  nand n81684(x81684, x81683, x73454);
  nand n81686(x81686, x68462, x81688);
  nand n81687(x81687, x81686, x73459);
  nand n81689(x81689, x68462, x81691);
  nand n81690(x81690, x81689, x73464);
  nand n81692(x81692, x68462, x81694);
  nand n81693(x81693, x81692, x73469);
  nand n81695(x81695, x68462, x81697);
  nand n81696(x81696, x81695, x73474);
  nand n81698(x81698, x68462, x81700);
  nand n81699(x81699, x81698, x73479);
  nand n81701(x81701, x68462, x81703);
  nand n81702(x81702, x81701, x73484);
  nand n81704(x81704, x68462, x81706);
  nand n81705(x81705, x81704, x73489);
  nand n81707(x81707, x68462, x81709);
  nand n81708(x81708, x81707, x73494);
  nand n81710(x81710, x68462, x81712);
  nand n81711(x81711, x81710, x73499);
  nand n81713(x81713, x68462, x81715);
  nand n81714(x81714, x81713, x73504);
  nand n81716(x81716, x68462, x81718);
  nand n81717(x81717, x81716, x73509);
  nand n81719(x81719, x68462, x81721);
  nand n81720(x81720, x81719, x73514);
  nand n81722(x81722, x68462, x81724);
  nand n81723(x81723, x81722, x73519);
  nand n81725(x81725, x68462, x81727);
  nand n81726(x81726, x81725, x73524);
  nand n81728(x81728, x68462, x81730);
  nand n81729(x81729, x81728, x73529);
  nand n81731(x81731, x68462, x81733);
  nand n81732(x81732, x81731, x73534);
  nand n81734(x81734, x68462, x81736);
  nand n81735(x81735, x81734, x73539);
  nand n81737(x81737, x68462, x81739);
  nand n81738(x81738, x81737, x73544);
  nand n81740(x81740, x68462, x81742);
  nand n81741(x81741, x81740, x73549);
  nand n81743(x81743, x68462, x81745);
  nand n81744(x81744, x81743, x73554);
  nand n81746(x81746, x68462, x81748);
  nand n81747(x81747, x81746, x73559);
  nand n81749(x81749, x68462, x81751);
  nand n81750(x81750, x81749, x73564);
  nand n81752(x81752, x68462, x81754);
  nand n81753(x81753, x81752, x73569);
  nand n81755(x81755, x68462, x81757);
  nand n81756(x81756, x81755, x73574);
  nand n81758(x81758, x68462, x81760);
  nand n81759(x81759, x81758, x73579);
  nand n81761(x81761, x68462, x81763);
  nand n81762(x81762, x81761, x73584);
  nand n81764(x81764, x68462, x81766);
  nand n81765(x81765, x81764, x73589);
  nand n81767(x81767, x68462, x81769);
  nand n81768(x81768, x81767, x73594);
  nand n81770(x81770, x68462, x81772);
  nand n81771(x81771, x81770, x73599);
  nand n81773(x81773, x68462, x81775);
  nand n81774(x81774, x81773, x73604);
  nand n81776(x81776, x68462, x81778);
  nand n81777(x81777, x81776, x73609);
  nand n81779(x81779, x68462, x81781);
  nand n81780(x81780, x81779, x73614);
  nand n81782(x81782, x68462, x81784);
  nand n81783(x81783, x81782, x73619);
  nand n81785(x81785, x68462, x81787);
  nand n81786(x81786, x81785, x73624);
  nand n81788(x81788, x68462, x81790);
  nand n81789(x81789, x81788, x73629);
  nand n81791(x81791, x68462, x81793);
  nand n81792(x81792, x81791, x73634);
  nand n81794(x81794, x68462, x81796);
  nand n81795(x81795, x81794, x73639);
  nand n81797(x81797, x68462, x81799);
  nand n81798(x81798, x81797, x73644);
  nand n81800(x81800, x68462, x81802);
  nand n81801(x81801, x81800, x73649);
  nand n81803(x81803, x68462, x81805);
  nand n81804(x81804, x81803, x73654);
  nand n81806(x81806, x68462, x81808);
  nand n81807(x81807, x81806, x73659);
  nand n81809(x81809, x68462, x81811);
  nand n81810(x81810, x81809, x73664);
  nand n81812(x81812, x68462, x81814);
  nand n81813(x81813, x81812, x73669);
  nand n81815(x81815, x68462, x81817);
  nand n81816(x81816, x81815, x73674);
  nand n81818(x81818, x68462, x81820);
  nand n81819(x81819, x81818, x73679);
  nand n81821(x81821, x68462, x81823);
  nand n81822(x81822, x81821, x73684);
  nand n81824(x81824, x68462, x81826);
  nand n81825(x81825, x81824, x73689);
  nand n81827(x81827, x68462, x81829);
  nand n81828(x81828, x81827, x73694);
  nand n81830(x81830, x68462, x81832);
  nand n81831(x81831, x81830, x73699);
  nand n81833(x81833, x68462, x81835);
  nand n81834(x81834, x81833, x73704);
  nand n81836(x81836, x68462, x81838);
  nand n81837(x81837, x81836, x73709);
  nand n81839(x81839, x68462, x81841);
  nand n81840(x81840, x81839, x73714);
  nand n81842(x81842, x68462, x81844);
  nand n81843(x81843, x81842, x73719);
  nand n81845(x81845, x68462, x81847);
  nand n81846(x81846, x81845, x73724);
  nand n81848(x81848, x68462, x81850);
  nand n81849(x81849, x81848, x73729);
  nand n81851(x81851, x68462, x81853);
  nand n81852(x81852, x81851, x73734);
  nand n81854(x81854, x68462, x81856);
  nand n81855(x81855, x81854, x73739);
  nand n81857(x81857, x68462, x81859);
  nand n81858(x81858, x81857, x73744);
  nand n81860(x81860, x68462, x81862);
  nand n81861(x81861, x81860, x73749);
  nand n81863(x81863, x68462, x81865);
  nand n81864(x81864, x81863, x73754);
  nand n81866(x81866, x68462, x81868);
  nand n81867(x81867, x81866, x73759);
  nand n81869(x81869, x68462, x81871);
  nand n81870(x81870, x81869, x73764);
  nand n81872(x81872, x68462, x81874);
  nand n81873(x81873, x81872, x73769);
  nand n81875(x81875, x68462, x81877);
  nand n81876(x81876, x81875, x73774);
  nand n81878(x81878, x68462, x81880);
  nand n81879(x81879, x81878, x73779);
  nand n81881(x81881, x68462, x81883);
  nand n81882(x81882, x81881, x73784);
  nand n81884(x81884, x68462, x81886);
  nand n81885(x81885, x81884, x73789);
  nand n81887(x81887, x68462, x81889);
  nand n81888(x81888, x81887, x73794);
  nand n81890(x81890, x68462, x81892);
  nand n81891(x81891, x81890, x73799);
  nand n81893(x81893, x68462, x81895);
  nand n81894(x81894, x81893, x73804);
  nand n81896(x81896, x68462, x81898);
  nand n81897(x81897, x81896, x73809);
  nand n81899(x81899, x68462, x81901);
  nand n81900(x81900, x81899, x73814);
  nand n81902(x81902, x68462, x81904);
  nand n81903(x81903, x81902, x73819);
  nand n81905(x81905, x68462, x81907);
  nand n81906(x81906, x81905, x73824);
  nand n81908(x81908, x68462, x81910);
  nand n81909(x81909, x81908, x73829);
  nand n81911(x81911, x68462, x81913);
  nand n81912(x81912, x81911, x73834);
  nand n81914(x81914, x68462, x81916);
  nand n81915(x81915, x81914, x73839);
  nand n81917(x81917, x68462, x81919);
  nand n81918(x81918, x81917, x73844);
  nand n81920(x81920, x68462, x81922);
  nand n81921(x81921, x81920, x73849);
  nand n81923(x81923, x68462, x81925);
  nand n81924(x81924, x81923, x73854);
  nand n81926(x81926, x68462, x81928);
  nand n81927(x81927, x81926, x73859);
  nand n81929(x81929, x68462, x81931);
  nand n81930(x81930, x81929, x73864);
  nand n81932(x81932, x68462, x81934);
  nand n81933(x81933, x81932, x73869);
  nand n81935(x81935, x68462, x81937);
  nand n81936(x81936, x81935, x73874);
  nand n81938(x81938, x68462, x81940);
  nand n81939(x81939, x81938, x73879);
  nand n81941(x81941, x68462, x81943);
  nand n81942(x81942, x81941, x73884);
  nand n81944(x81944, x68462, x81946);
  nand n81945(x81945, x81944, x73889);
  nand n81947(x81947, x68462, x81949);
  nand n81948(x81948, x81947, x73894);
  nand n81950(x81950, x68462, x81952);
  nand n81951(x81951, x81950, x73899);
  nand n81953(x81953, x68462, x81955);
  nand n81954(x81954, x81953, x73904);
  nand n81956(x81956, x68462, x81958);
  nand n81957(x81957, x81956, x73909);
  nand n81959(x81959, x68462, x81961);
  nand n81960(x81960, x81959, x73914);
  nand n81962(x81962, x68462, x81964);
  nand n81963(x81963, x81962, x73919);
  nand n81965(x81965, x68462, x81967);
  nand n81966(x81966, x81965, x73924);
  nand n81968(x81968, x68462, x81970);
  nand n81969(x81969, x81968, x73929);
  nand n81971(x81971, x68462, x81973);
  nand n81972(x81972, x81971, x73934);
  nand n81974(x81974, x68462, x81976);
  nand n81975(x81975, x81974, x73939);
  nand n81977(x81977, x68462, x81979);
  nand n81978(x81978, x81977, x73944);
  nand n81980(x81980, x68462, x81982);
  nand n81981(x81981, x81980, x73949);
  nand n81983(x81983, x68462, x81985);
  nand n81984(x81984, x81983, x73954);
  nand n81986(x81986, x68462, x81988);
  nand n81987(x81987, x81986, x73959);
  nand n81989(x81989, x68462, x81991);
  nand n81990(x81990, x81989, x73964);
  nand n81992(x81992, x68462, x81994);
  nand n81993(x81993, x81992, x73969);
  nand n81995(x81995, x68462, x81997);
  nand n81996(x81996, x81995, x73974);
  nand n81998(x81998, x68462, x82000);
  nand n81999(x81999, x81998, x73979);
  nand n82001(x82001, x68462, x82003);
  nand n82002(x82002, x82001, x73984);
  nand n82004(x82004, x68462, x82006);
  nand n82005(x82005, x82004, x73989);
  nand n82007(x82007, x68462, x82009);
  nand n82008(x82008, x82007, x73994);
  nand n82010(x82010, x68462, x82012);
  nand n82011(x82011, x82010, x73999);
  nand n82013(x82013, x68462, x82015);
  nand n82014(x82014, x82013, x71799);
  nand n82016(x82016, x68462, x82018);
  nand n82017(x82017, x82016, x71804);
  nand n82019(x82019, x68462, x82021);
  nand n82020(x82020, x82019, x71809);
  nand n82022(x82022, x68462, x82024);
  nand n82023(x82023, x82022, x71814);
  nand n82025(x82025, x68462, x82027);
  nand n82026(x82026, x82025, x71819);
  nand n82028(x82028, x68462, x82030);
  nand n82029(x82029, x82028, x71824);
  nand n82031(x82031, x68462, x82033);
  nand n82032(x82032, x82031, x71829);
  nand n82034(x82034, x68462, x82036);
  nand n82035(x82035, x82034, x71834);
  nand n82037(x82037, x68462, x82039);
  nand n82038(x82038, x82037, x71839);
  nand n82040(x82040, x68462, x82042);
  nand n82041(x82041, x82040, x71844);
  nand n82043(x82043, x68462, x82045);
  nand n82044(x82044, x82043, x71849);
  nand n82046(x82046, x68462, x82048);
  nand n82047(x82047, x82046, x71854);
  nand n82049(x82049, x68462, x82051);
  nand n82050(x82050, x82049, x71859);
  nand n82052(x82052, x68462, x82054);
  nand n82053(x82053, x82052, x71864);
  nand n82055(x82055, x68462, x82057);
  nand n82056(x82056, x82055, x71869);
  nand n82058(x82058, x68462, x82060);
  nand n82059(x82059, x82058, x71874);
  nand n82061(x82061, x68462, x82063);
  nand n82062(x82062, x82061, x71879);
  nand n82064(x82064, x68462, x82066);
  nand n82065(x82065, x82064, x71884);
  nand n82067(x82067, x68462, x82069);
  nand n82068(x82068, x82067, x71889);
  nand n82070(x82070, x68462, x82072);
  nand n82071(x82071, x82070, x71894);
  nand n82073(x82073, x68462, x82075);
  nand n82074(x82074, x82073, x71899);
  nand n82076(x82076, x68462, x82078);
  nand n82077(x82077, x82076, x71904);
  nand n82079(x82079, x68462, x82081);
  nand n82080(x82080, x82079, x71904);
  nand n82082(x82082, x68462, x82084);
  nand n82083(x82083, x82082, x71904);
  nand n82085(x82085, x68462, x82087);
  nand n82086(x82086, x82085, x71904);
  nand n82088(x82088, x68462, x82090);
  nand n82089(x82089, x82088, x71904);
  nand n82091(x82091, x68462, x82093);
  nand n82092(x82092, x82091, x71904);
  nand n82094(x82094, x68462, x82096);
  nand n82095(x82095, x82094, x71904);
  nand n82097(x82097, x68462, x82099);
  nand n82098(x82098, x82097, x71904);
  nand n82100(x82100, x68462, x82102);
  nand n82101(x82101, x82100, x71904);
  nand n82103(x82103, x68462, x82105);
  nand n82104(x82104, x82103, x71904);
  nand n82106(x82106, x68462, x82108);
  nand n82107(x82107, x82106, x71904);
  nand n82109(x82109, x68462, x82111);
  nand n82110(x82110, x82109, x71939);
  nand n82112(x82112, x68462, x82114);
  nand n82113(x82113, x82112, x71944);
  nand n82115(x82115, x68462, x82117);
  nand n82116(x82116, x82115, x71949);
  nand n82118(x82118, x68462, x82120);
  nand n82119(x82119, x82118, x71954);
  nand n82121(x82121, x68462, x82123);
  nand n82122(x82122, x82121, x71959);
  nand n82124(x82124, x68462, x82126);
  nand n82125(x82125, x82124, x71964);
  nand n82127(x82127, x68462, x82129);
  nand n82128(x82128, x82127, x71969);
  nand n82130(x82130, x68462, x82132);
  nand n82131(x82131, x82130, x71974);
  nand n82133(x82133, x68462, x82135);
  nand n82134(x82134, x82133, x71979);
  nand n82136(x82136, x68462, x82138);
  nand n82137(x82137, x82136, x71984);
  nand n82139(x82139, x68462, x82141);
  nand n82140(x82140, x82139, x71989);
  nand n82142(x82142, x68462, x82144);
  nand n82143(x82143, x82142, x71994);
  nand n82145(x82145, x68462, x82147);
  nand n82146(x82146, x82145, x71999);
  nand n82148(x82148, x68462, x82150);
  nand n82149(x82149, x82148, x72004);
  nand n82151(x82151, x68462, x82153);
  nand n82152(x82152, x82151, x72009);
  nand n82154(x82154, x68462, x82156);
  nand n82155(x82155, x82154, x72014);
  nand n82157(x82157, x68462, x82159);
  nand n82158(x82158, x82157, x72019);
  nand n82160(x82160, x68462, x82162);
  nand n82161(x82161, x82160, x72024);
  nand n82163(x82163, x68462, x82165);
  nand n82164(x82164, x82163, x72029);
  nand n82166(x82166, x68462, x82168);
  nand n82167(x82167, x82166, x72034);
  nand n82169(x82169, x68462, x82171);
  nand n82170(x82170, x82169, x72039);
  nand n82172(x82172, x68462, x82174);
  nand n82173(x82173, x82172, x72044);
  nand n82175(x82175, x68462, x82177);
  nand n82176(x82176, x82175, x72049);
  nand n82178(x82178, x68462, x82180);
  nand n82179(x82179, x82178, x72054);
  nand n82181(x82181, x68462, x82183);
  nand n82182(x82182, x82181, x72059);
  nand n82184(x82184, x68462, x82186);
  nand n82185(x82185, x82184, x72064);
  nand n82187(x82187, x68462, x82189);
  nand n82188(x82188, x82187, x72069);
  nand n82190(x82190, x68462, x82192);
  nand n82191(x82191, x82190, x72074);
  nand n82193(x82193, x68462, x82195);
  nand n82194(x82194, x82193, x72079);
  nand n82196(x82196, x68462, x82198);
  nand n82197(x82197, x82196, x72084);
  nand n82199(x82199, x68462, x82201);
  nand n82200(x82200, x82199, x72089);
  nand n82202(x82202, x68462, x82204);
  nand n82203(x82203, x82202, x72094);
  nand n82205(x82205, x68462, x82207);
  nand n82206(x82206, x82205, x72099);
  nand n82208(x82208, x68462, x82210);
  nand n82209(x82209, x82208, x72104);
  nand n82211(x82211, x68462, x82213);
  nand n82212(x82212, x82211, x72109);
  nand n82214(x82214, x68462, x82216);
  nand n82215(x82215, x82214, x72114);
  nand n82217(x82217, x68462, x82219);
  nand n82218(x82218, x82217, x72119);
  nand n82220(x82220, x68462, x82222);
  nand n82221(x82221, x82220, x72124);
  nand n82223(x82223, x68462, x82225);
  nand n82224(x82224, x82223, x72129);
  nand n82226(x82226, x68462, x82228);
  nand n82227(x82227, x82226, x72134);
  nand n82229(x82229, x68462, x82231);
  nand n82230(x82230, x82229, x72139);
  nand n82232(x82232, x68462, x82234);
  nand n82233(x82233, x82232, x72144);
  nand n82235(x82235, x68462, x82237);
  nand n82236(x82236, x82235, x72149);
  nand n82238(x82238, x68462, x82240);
  nand n82239(x82239, x82238, x72154);
  nand n82241(x82241, x68462, x82243);
  nand n82242(x82242, x82241, x72159);
  nand n82244(x82244, x68462, x82246);
  nand n82245(x82245, x82244, x72164);
  nand n82247(x82247, x68462, x82249);
  nand n82248(x82248, x82247, x72169);
  nand n82250(x82250, x68462, x82252);
  nand n82251(x82251, x82250, x72174);
  nand n82253(x82253, x68462, x82255);
  nand n82254(x82254, x82253, x72179);
  nand n82256(x82256, x68462, x82258);
  nand n82257(x82257, x82256, x72184);
  nand n82259(x82259, x68462, x82261);
  nand n82260(x82260, x82259, x72189);
  nand n82262(x82262, x68462, x82264);
  nand n82263(x82263, x82262, x72194);
  nand n82265(x82265, x68462, x82267);
  nand n82266(x82266, x82265, x72199);
  nand n82268(x82268, x68462, x82270);
  nand n82269(x82269, x82268, x72204);
  nand n82271(x82271, x68462, x82273);
  nand n82272(x82272, x82271, x72209);
  nand n82274(x82274, x68462, x82276);
  nand n82275(x82275, x82274, x72214);
  nand n82277(x82277, x68462, x82279);
  nand n82278(x82278, x82277, x72219);
  nand n82280(x82280, x68462, x82282);
  nand n82281(x82281, x82280, x72224);
  nand n82283(x82283, x68462, x82285);
  nand n82284(x82284, x82283, x72229);
  nand n82286(x82286, x68462, x82288);
  nand n82287(x82287, x82286, x72234);
  nand n82289(x82289, x68462, x82291);
  nand n82290(x82290, x82289, x72239);
  nand n82292(x82292, x68462, x82294);
  nand n82293(x82293, x82292, x72244);
  nand n82295(x82295, x68462, x82297);
  nand n82296(x82296, x82295, x72249);
  nand n82298(x82298, x68462, x82300);
  nand n82299(x82299, x82298, x72254);
  nand n82301(x82301, x68462, x82303);
  nand n82302(x82302, x82301, x72259);
  nand n82304(x82304, x68462, x82306);
  nand n82305(x82305, x82304, x72264);
  nand n82307(x82307, x68462, x82309);
  nand n82308(x82308, x82307, x72269);
  nand n82310(x82310, x68462, x82312);
  nand n82311(x82311, x82310, x72274);
  nand n82313(x82313, x68462, x82315);
  nand n82314(x82314, x82313, x72279);
  nand n82316(x82316, x68462, x82318);
  nand n82317(x82317, x82316, x72284);
  nand n82319(x82319, x68462, x82321);
  nand n82320(x82320, x82319, x72289);
  nand n82322(x82322, x68462, x82324);
  nand n82323(x82323, x82322, x72294);
  nand n82325(x82325, x68462, x82327);
  nand n82326(x82326, x82325, x72299);
  nand n82328(x82328, x68462, x82330);
  nand n82329(x82329, x82328, x72304);
  nand n82331(x82331, x68462, x82333);
  nand n82332(x82332, x82331, x72309);
  nand n82334(x82334, x68462, x82336);
  nand n82335(x82335, x82334, x72314);
  nand n82337(x82337, x68462, x82339);
  nand n82338(x82338, x82337, x72319);
  nand n82340(x82340, x68462, x82342);
  nand n82341(x82341, x82340, x72324);
  nand n82343(x82343, x68462, x82345);
  nand n82344(x82344, x82343, x72329);
  nand n82346(x82346, x68462, x82348);
  nand n82347(x82347, x82346, x72334);
  nand n82349(x82349, x68462, x82351);
  nand n82350(x82350, x82349, x72339);
  nand n82352(x82352, x68462, x82354);
  nand n82353(x82353, x82352, x72344);
  nand n82355(x82355, x68462, x82357);
  nand n82356(x82356, x82355, x72349);
  nand n82358(x82358, x68462, x82360);
  nand n82359(x82359, x82358, x72354);
  nand n82361(x82361, x68462, x82363);
  nand n82362(x82362, x82361, x72359);
  nand n82364(x82364, x68462, x82366);
  nand n82365(x82365, x82364, x72364);
  nand n82367(x82367, x68462, x82369);
  nand n82368(x82368, x82367, x72369);
  nand n82370(x82370, x68462, x82372);
  nand n82371(x82371, x82370, x72374);
  nand n82373(x82373, x68462, x82375);
  nand n82374(x82374, x82373, x72379);
  nand n82376(x82376, x68462, x82378);
  nand n82377(x82377, x82376, x72384);
  nand n82379(x82379, x68462, x82381);
  nand n82380(x82380, x82379, x72389);
  nand n82382(x82382, x68462, x82384);
  nand n82383(x82383, x82382, x72394);
  nand n82385(x82385, x68462, x82387);
  nand n82386(x82386, x82385, x72399);
  nand n82388(x82388, x68462, x82390);
  nand n82389(x82389, x82388, x72404);
  nand n82391(x82391, x68462, x82393);
  nand n82392(x82392, x82391, x72409);
  nand n82394(x82394, x68462, x82396);
  nand n82395(x82395, x82394, x72414);
  nand n82397(x82397, x68462, x82399);
  nand n82398(x82398, x82397, x72419);
  nand n82400(x82400, x68462, x82402);
  nand n82401(x82401, x82400, x72424);
  nand n82403(x82403, x68462, x82405);
  nand n82404(x82404, x82403, x72429);
  nand n82406(x82406, x68462, x82408);
  nand n82407(x82407, x82406, x72434);
  nand n82409(x82409, x68462, x82411);
  nand n82410(x82410, x82409, x72439);
  nand n82412(x82412, x68462, x82414);
  nand n82413(x82413, x82412, x72444);
  nand n82415(x82415, x68462, x82417);
  nand n82416(x82416, x82415, x72449);
  nand n82418(x82418, x68462, x82420);
  nand n82419(x82419, x82418, x72454);
  nand n82421(x82421, x68462, x82423);
  nand n82422(x82422, x82421, x72459);
  nand n82424(x82424, x68462, x82426);
  nand n82425(x82425, x82424, x72464);
  nand n82427(x82427, x68462, x82429);
  nand n82428(x82428, x82427, x72469);
  nand n82430(x82430, x68462, x82432);
  nand n82431(x82431, x82430, x72474);
  nand n82433(x82433, x68462, x82435);
  nand n82434(x82434, x82433, x72479);
  nand n82436(x82436, x68462, x82438);
  nand n82437(x82437, x82436, x72484);
  nand n82439(x82439, x68462, x82441);
  nand n82440(x82440, x82439, x72489);
  nand n82442(x82442, x68462, x82444);
  nand n82443(x82443, x82442, x72494);
  nand n82445(x82445, x68462, x82447);
  nand n82446(x82446, x82445, x72499);
  nand n82448(x82448, x68462, x82450);
  nand n82449(x82449, x82448, x72504);
  nand n82451(x82451, x68462, x82453);
  nand n82452(x82452, x82451, x72509);
  nand n82454(x82454, x68462, x82456);
  nand n82455(x82455, x82454, x72514);
  nand n82457(x82457, x68462, x82459);
  nand n82458(x82458, x82457, x72519);
  nand n82460(x82460, x68462, x82462);
  nand n82461(x82461, x82460, x72524);
  nand n82463(x82463, x68462, x82465);
  nand n82464(x82464, x82463, x72529);
  nand n82466(x82466, x68462, x82468);
  nand n82467(x82467, x82466, x72534);
  nand n82469(x82469, x68462, x82471);
  nand n82470(x82470, x82469, x72539);
  nand n82472(x82472, x68462, x82474);
  nand n82473(x82473, x82472, x72544);
  nand n82475(x82475, x68462, x82477);
  nand n82476(x82476, x82475, x72549);
  nand n82478(x82478, x68462, x82480);
  nand n82479(x82479, x82478, x72554);
  nand n82481(x82481, x68462, x82483);
  nand n82482(x82482, x82481, x72559);
  nand n82484(x82484, x68462, x82486);
  nand n82485(x82485, x82484, x72564);
  nand n82487(x82487, x68462, x82489);
  nand n82488(x82488, x82487, x72569);
  nand n82490(x82490, x68462, x82492);
  nand n82491(x82491, x82490, x72574);
  nand n82493(x82493, x68462, x82495);
  nand n82494(x82494, x82493, x72579);
  nand n82496(x82496, x68462, x82498);
  nand n82497(x82497, x82496, x72584);
  nand n82499(x82499, x68462, x82501);
  nand n82500(x82500, x82499, x72589);
  nand n82502(x82502, x68462, x82504);
  nand n82503(x82503, x82502, x72594);
  nand n82505(x82505, x68462, x82507);
  nand n82506(x82506, x82505, x72599);
  nand n82508(x82508, x68462, x82510);
  nand n82509(x82509, x82508, x72604);
  nand n82511(x82511, x68462, x82513);
  nand n82512(x82512, x82511, x72609);
  nand n82514(x82514, x68462, x82516);
  nand n82515(x82515, x82514, x72614);
  nand n82517(x82517, x68462, x82519);
  nand n82518(x82518, x82517, x72619);
  nand n82520(x82520, x68462, x82522);
  nand n82521(x82521, x82520, x72624);
  nand n82523(x82523, x68462, x82525);
  nand n82524(x82524, x82523, x72629);
  nand n82526(x82526, x68462, x82528);
  nand n82527(x82527, x82526, x72634);
  nand n82529(x82529, x68462, x82531);
  nand n82530(x82530, x82529, x72639);
  nand n82532(x82532, x68462, x82534);
  nand n82533(x82533, x82532, x72644);
  nand n82535(x82535, x68462, x82537);
  nand n82536(x82536, x82535, x72649);
  nand n82538(x82538, x68462, x82540);
  nand n82539(x82539, x82538, x72654);
  nand n82541(x82541, x68462, x82543);
  nand n82542(x82542, x82541, x72659);
  nand n82544(x82544, x68462, x82546);
  nand n82545(x82545, x82544, x72664);
  nand n82547(x82547, x68462, x82549);
  nand n82548(x82548, x82547, x72669);
  nand n82550(x82550, x68462, x82552);
  nand n82551(x82551, x82550, x72674);
  nand n82553(x82553, x68462, x82555);
  nand n82554(x82554, x82553, x72679);
  nand n82556(x82556, x68462, x82558);
  nand n82557(x82557, x82556, x72684);
  nand n82559(x82559, x68462, x82561);
  nand n82560(x82560, x82559, x72689);
  nand n82562(x82562, x68462, x82564);
  nand n82563(x82563, x82562, x72694);
  nand n82565(x82565, x68462, x82567);
  nand n82566(x82566, x82565, x72699);
  nand n82568(x82568, x68462, x82570);
  nand n82569(x82569, x82568, x72704);
  nand n82571(x82571, x68462, x82573);
  nand n82572(x82572, x82571, x72709);
  nand n82574(x82574, x68462, x82576);
  nand n82575(x82575, x82574, x72714);
  nand n82577(x82577, x68462, x82579);
  nand n82578(x82578, x82577, x72719);
  nand n82580(x82580, x68462, x82582);
  nand n82581(x82581, x82580, x72724);
  nand n82583(x82583, x68462, x82585);
  nand n82584(x82584, x82583, x72729);
  nand n82586(x82586, x68462, x82588);
  nand n82587(x82587, x82586, x72734);
  nand n82589(x82589, x68462, x82591);
  nand n82590(x82590, x82589, x72739);
  nand n82592(x82592, x68462, x82594);
  nand n82593(x82593, x82592, x72744);
  nand n82595(x82595, x68462, x82597);
  nand n82596(x82596, x82595, x72749);
  nand n82598(x82598, x68462, x82600);
  nand n82599(x82599, x82598, x72754);
  nand n82601(x82601, x68462, x82603);
  nand n82602(x82602, x82601, x72759);
  nand n82604(x82604, x68462, x82606);
  nand n82605(x82605, x82604, x72764);
  nand n82607(x82607, x68462, x82609);
  nand n82608(x82608, x82607, x72769);
  nand n82610(x82610, x68462, x82612);
  nand n82611(x82611, x82610, x72774);
  nand n82613(x82613, x68462, x82615);
  nand n82614(x82614, x82613, x72779);
  nand n82616(x82616, x68462, x82618);
  nand n82617(x82617, x82616, x72784);
  nand n82619(x82619, x68462, x82621);
  nand n82620(x82620, x82619, x72789);
  nand n82622(x82622, x68462, x82624);
  nand n82623(x82623, x82622, x72794);
  nand n82625(x82625, x68462, x82627);
  nand n82626(x82626, x82625, x72799);
  nand n82628(x82628, x68462, x82630);
  nand n82629(x82629, x82628, x72804);
  nand n82631(x82631, x68462, x82633);
  nand n82632(x82632, x82631, x72809);
  nand n82634(x82634, x68462, x82636);
  nand n82635(x82635, x82634, x72814);
  nand n82637(x82637, x68462, x82639);
  nand n82638(x82638, x82637, x72819);
  nand n82640(x82640, x68462, x82642);
  nand n82641(x82641, x82640, x72824);
  nand n82643(x82643, x68462, x82645);
  nand n82644(x82644, x82643, x72829);
  nand n82646(x82646, x68462, x82648);
  nand n82647(x82647, x82646, x72834);
  nand n82649(x82649, x68462, x82651);
  nand n82650(x82650, x82649, x72839);
  nand n82652(x82652, x68462, x82654);
  nand n82653(x82653, x82652, x72844);
  nand n82655(x82655, x68462, x82657);
  nand n82656(x82656, x82655, x72849);
  nand n82658(x82658, x68462, x82660);
  nand n82659(x82659, x82658, x72854);
  nand n82661(x82661, x68462, x82663);
  nand n82662(x82662, x82661, x72859);
  nand n82664(x82664, x68462, x82666);
  nand n82665(x82665, x82664, x72864);
  nand n82667(x82667, x68462, x82669);
  nand n82668(x82668, x82667, x72869);
  nand n82670(x82670, x68462, x82672);
  nand n82671(x82671, x82670, x72874);
  nand n82673(x82673, x68462, x82675);
  nand n82674(x82674, x82673, x72879);
  nand n82676(x82676, x68462, x82678);
  nand n82677(x82677, x82676, x72884);
  nand n82679(x82679, x68462, x82681);
  nand n82680(x82680, x82679, x72889);
  nand n82682(x82682, x68462, x82684);
  nand n82683(x82683, x82682, x72894);
  nand n82685(x82685, x68462, x82687);
  nand n82686(x82686, x82685, x72899);
  nand n82688(x82688, x68462, x82690);
  nand n82689(x82689, x82688, x72904);
  nand n82691(x82691, x68462, x82693);
  nand n82692(x82692, x82691, x72909);
  nand n82694(x82694, x68462, x82696);
  nand n82695(x82695, x82694, x72914);
  nand n82697(x82697, x68462, x82699);
  nand n82698(x82698, x82697, x72919);
  nand n82700(x82700, x68462, x82702);
  nand n82701(x82701, x82700, x72924);
  nand n82703(x82703, x68462, x82705);
  nand n82704(x82704, x82703, x72929);
  nand n82706(x82706, x68462, x82708);
  nand n82707(x82707, x82706, x72934);
  nand n82709(x82709, x68462, x82711);
  nand n82710(x82710, x82709, x72939);
  nand n82712(x82712, x68462, x82714);
  nand n82713(x82713, x82712, x72944);
  nand n82715(x82715, x68462, x82717);
  nand n82716(x82716, x82715, x72949);
  nand n82718(x82718, x68462, x82720);
  nand n82719(x82719, x82718, x72954);
  nand n82721(x82721, x68462, x82723);
  nand n82722(x82722, x82721, x72959);
  nand n82724(x82724, x68462, x82726);
  nand n82725(x82725, x82724, x72964);
  nand n82727(x82727, x68462, x82729);
  nand n82728(x82728, x82727, x72969);
  nand n82730(x82730, x68462, x82732);
  nand n82731(x82731, x82730, x72974);
  nand n82733(x82733, x68462, x82735);
  nand n82734(x82734, x82733, x72979);
  nand n82736(x82736, x68462, x82738);
  nand n82737(x82737, x82736, x72984);
  nand n82739(x82739, x68462, x82741);
  nand n82740(x82740, x82739, x72989);
  nand n82742(x82742, x68462, x82744);
  nand n82743(x82743, x82742, x72994);
  nand n82745(x82745, x68462, x82747);
  nand n82746(x82746, x82745, x72999);
  nand n82748(x82748, x68462, x82750);
  nand n82749(x82749, x82748, x73004);
  nand n82751(x82751, x68462, x82753);
  nand n82752(x82752, x82751, x73009);
  nand n82754(x82754, x68462, x82756);
  nand n82755(x82755, x82754, x73014);
  nand n82757(x82757, x68462, x82759);
  nand n82758(x82758, x82757, x73019);
  nand n82760(x82760, x68462, x82762);
  nand n82761(x82761, x82760, x73024);
  nand n82763(x82763, x68462, x82765);
  nand n82764(x82764, x82763, x73029);
  nand n82766(x82766, x68462, x82768);
  nand n82767(x82767, x82766, x73034);
  nand n82769(x82769, x68462, x82771);
  nand n82770(x82770, x82769, x73039);
  nand n82772(x82772, x68462, x82774);
  nand n82773(x82773, x82772, x73044);
  nand n82775(x82775, x68462, x82777);
  nand n82776(x82776, x82775, x73049);
  nand n82778(x82778, x68462, x82780);
  nand n82779(x82779, x82778, x73054);
  nand n82781(x82781, x68462, x82783);
  nand n82782(x82782, x82781, x73059);
  nand n82784(x82784, x68462, x82786);
  nand n82785(x82785, x82784, x73064);
  nand n82787(x82787, x68462, x82789);
  nand n82788(x82788, x82787, x73069);
  nand n82790(x82790, x68462, x82792);
  nand n82791(x82791, x82790, x73074);
  nand n82793(x82793, x68462, x82795);
  nand n82794(x82794, x82793, x73079);
  nand n82796(x82796, x68462, x82798);
  nand n82797(x82797, x82796, x73084);
  nand n82799(x82799, x68462, x82801);
  nand n82800(x82800, x82799, x73089);
  nand n82802(x82802, x68462, x82804);
  nand n82803(x82803, x82802, x73094);
  nand n82805(x82805, x68462, x82807);
  nand n82806(x82806, x82805, x73099);
  nand n82808(x82808, x68462, x82810);
  nand n82809(x82809, x82808, x73104);
  nand n82811(x82811, x68462, x82813);
  nand n82812(x82812, x82811, x73109);
  nand n82814(x82814, x68462, x82816);
  nand n82815(x82815, x82814, x73114);
  nand n82817(x82817, x68462, x82819);
  nand n82818(x82818, x82817, x73119);
  nand n82820(x82820, x68462, x82822);
  nand n82821(x82821, x82820, x73124);
  nand n82823(x82823, x68462, x82825);
  nand n82824(x82824, x82823, x73129);
  nand n82826(x82826, x68462, x82828);
  nand n82827(x82827, x82826, x73134);
  nand n82829(x82829, x68462, x82831);
  nand n82830(x82830, x82829, x73139);
  nand n82832(x82832, x68462, x82834);
  nand n82833(x82833, x82832, x73144);
  nand n82835(x82835, x68462, x82837);
  nand n82836(x82836, x82835, x73149);
  nand n82838(x82838, x68462, x82840);
  nand n82839(x82839, x82838, x73154);
  nand n82841(x82841, x68462, x82843);
  nand n82842(x82842, x82841, x73159);
  nand n82844(x82844, x68462, x82846);
  nand n82845(x82845, x82844, x73164);
  nand n82847(x82847, x68462, x82849);
  nand n82848(x82848, x82847, x73169);
  nand n82850(x82850, x68462, x82852);
  nand n82851(x82851, x82850, x73174);
  nand n82853(x82853, x68462, x82855);
  nand n82854(x82854, x82853, x73179);
  nand n82856(x82856, x68462, x82858);
  nand n82857(x82857, x82856, x73184);
  nand n82859(x82859, x68462, x82861);
  nand n82860(x82860, x82859, x73189);
  nand n82862(x82862, x68462, x82864);
  nand n82863(x82863, x82862, x73194);
  nand n82865(x82865, x68462, x82867);
  nand n82866(x82866, x82865, x73199);
  nand n82868(x82868, x68462, x82870);
  nand n82869(x82869, x82868, x73204);
  nand n82871(x82871, x68462, x82873);
  nand n82872(x82872, x82871, x73209);
  nand n82874(x82874, x68462, x82876);
  nand n82875(x82875, x82874, x73214);
  nand n82877(x82877, x68462, x82879);
  nand n82878(x82878, x82877, x73219);
  nand n82880(x82880, x68462, x82882);
  nand n82881(x82881, x82880, x73224);
  nand n82883(x82883, x68462, x82885);
  nand n82884(x82884, x82883, x73229);
  nand n82886(x82886, x68462, x82888);
  nand n82887(x82887, x82886, x73234);
  nand n82889(x82889, x68462, x82891);
  nand n82890(x82890, x82889, x73239);
  nand n82892(x82892, x68462, x82894);
  nand n82893(x82893, x82892, x73244);
  nand n82895(x82895, x68462, x82897);
  nand n82896(x82896, x82895, x73249);
  nand n82898(x82898, x68462, x82900);
  nand n82899(x82899, x82898, x73254);
  nand n82901(x82901, x68462, x82903);
  nand n82902(x82902, x82901, x73259);
  nand n82904(x82904, x68462, x82906);
  nand n82905(x82905, x82904, x73264);
  nand n82907(x82907, x68462, x82909);
  nand n82908(x82908, x82907, x73269);
  nand n82910(x82910, x68462, x82912);
  nand n82911(x82911, x82910, x73274);
  nand n82913(x82913, x68462, x82915);
  nand n82914(x82914, x82913, x73279);
  nand n82916(x82916, x68462, x82918);
  nand n82917(x82917, x82916, x73284);
  nand n82919(x82919, x68462, x82921);
  nand n82920(x82920, x82919, x73289);
  nand n82922(x82922, x68462, x82924);
  nand n82923(x82923, x82922, x73294);
  nand n82925(x82925, x68462, x82927);
  nand n82926(x82926, x82925, x73299);
  nand n82928(x82928, x68462, x82930);
  nand n82929(x82929, x82928, x73304);
  nand n82931(x82931, x68462, x82933);
  nand n82932(x82932, x82931, x73309);
  nand n82934(x82934, x68462, x82936);
  nand n82935(x82935, x82934, x73314);
  nand n82937(x82937, x68462, x82939);
  nand n82938(x82938, x82937, x73319);
  nand n82940(x82940, x68462, x82942);
  nand n82941(x82941, x82940, x73324);
  nand n82943(x82943, x68462, x82945);
  nand n82944(x82944, x82943, x73329);
  nand n82946(x82946, x68462, x82948);
  nand n82947(x82947, x82946, x73334);
  nand n82949(x82949, x68462, x82951);
  nand n82950(x82950, x82949, x73339);
  nand n82952(x82952, x68462, x82954);
  nand n82953(x82953, x82952, x73344);
  nand n82955(x82955, x68462, x82957);
  nand n82956(x82956, x82955, x73349);
  nand n82958(x82958, x68462, x82960);
  nand n82959(x82959, x82958, x73354);
  nand n82961(x82961, x68462, x82963);
  nand n82962(x82962, x82961, x73359);
  nand n82964(x82964, x68462, x82966);
  nand n82965(x82965, x82964, x73364);
  nand n82967(x82967, x68462, x82969);
  nand n82968(x82968, x82967, x73369);
  nand n82970(x82970, x68462, x82972);
  nand n82971(x82971, x82970, x73374);
  nand n82973(x82973, x68462, x82975);
  nand n82974(x82974, x82973, x73379);
  nand n82976(x82976, x68462, x82978);
  nand n82977(x82977, x82976, x73384);
  nand n82979(x82979, x68462, x82981);
  nand n82980(x82980, x82979, x73389);
  nand n82982(x82982, x68462, x82984);
  nand n82983(x82983, x82982, x73394);
  nand n82985(x82985, x68462, x82987);
  nand n82986(x82986, x82985, x73399);
  nand n82988(x82988, x68462, x82990);
  nand n82989(x82989, x82988, x73404);
  nand n82991(x82991, x68462, x82993);
  nand n82992(x82992, x82991, x73409);
  nand n82994(x82994, x68462, x82996);
  nand n82995(x82995, x82994, x73414);
  nand n82997(x82997, x68462, x82999);
  nand n82998(x82998, x82997, x73419);
  nand n83000(x83000, x68462, x83002);
  nand n83001(x83001, x83000, x73424);
  nand n83003(x83003, x68462, x83005);
  nand n83004(x83004, x83003, x73429);
  nand n83006(x83006, x68462, x83008);
  nand n83007(x83007, x83006, x73434);
  nand n83009(x83009, x68462, x83011);
  nand n83010(x83010, x83009, x73439);
  nand n83012(x83012, x68462, x83014);
  nand n83013(x83013, x83012, x73444);
  nand n83015(x83015, x68462, x83017);
  nand n83016(x83016, x83015, x73449);
  nand n83018(x83018, x68462, x83020);
  nand n83019(x83019, x83018, x73454);
  nand n83021(x83021, x68462, x83023);
  nand n83022(x83022, x83021, x73459);
  nand n83024(x83024, x68462, x83026);
  nand n83025(x83025, x83024, x73464);
  nand n83027(x83027, x68462, x83029);
  nand n83028(x83028, x83027, x73469);
  nand n83030(x83030, x68462, x83032);
  nand n83031(x83031, x83030, x73474);
  nand n83033(x83033, x68462, x83035);
  nand n83034(x83034, x83033, x73479);
  nand n83036(x83036, x68462, x83038);
  nand n83037(x83037, x83036, x73484);
  nand n83039(x83039, x68462, x83041);
  nand n83040(x83040, x83039, x73489);
  nand n83042(x83042, x68462, x83044);
  nand n83043(x83043, x83042, x73494);
  nand n83045(x83045, x68462, x83047);
  nand n83046(x83046, x83045, x73499);
  nand n83048(x83048, x68462, x83050);
  nand n83049(x83049, x83048, x73504);
  nand n83051(x83051, x68462, x83053);
  nand n83052(x83052, x83051, x73509);
  nand n83054(x83054, x68462, x83056);
  nand n83055(x83055, x83054, x73514);
  nand n83057(x83057, x68462, x83059);
  nand n83058(x83058, x83057, x73519);
  nand n83060(x83060, x68462, x83062);
  nand n83061(x83061, x83060, x73524);
  nand n83063(x83063, x68462, x83065);
  nand n83064(x83064, x83063, x73529);
  nand n83066(x83066, x68462, x83068);
  nand n83067(x83067, x83066, x73534);
  nand n83069(x83069, x68462, x83071);
  nand n83070(x83070, x83069, x73539);
  nand n83072(x83072, x68462, x83074);
  nand n83073(x83073, x83072, x73544);
  nand n83075(x83075, x68462, x83077);
  nand n83076(x83076, x83075, x73549);
  nand n83078(x83078, x68462, x83080);
  nand n83079(x83079, x83078, x73554);
  nand n83081(x83081, x68462, x83083);
  nand n83082(x83082, x83081, x73559);
  nand n83084(x83084, x68462, x83086);
  nand n83085(x83085, x83084, x73564);
  nand n83087(x83087, x68462, x83089);
  nand n83088(x83088, x83087, x73569);
  nand n83090(x83090, x68462, x83092);
  nand n83091(x83091, x83090, x73574);
  nand n83093(x83093, x68462, x83095);
  nand n83094(x83094, x83093, x73579);
  nand n83096(x83096, x68462, x83098);
  nand n83097(x83097, x83096, x73584);
  nand n83099(x83099, x68462, x83101);
  nand n83100(x83100, x83099, x73589);
  nand n83102(x83102, x68462, x83104);
  nand n83103(x83103, x83102, x73594);
  nand n83105(x83105, x68462, x83107);
  nand n83106(x83106, x83105, x73599);
  nand n83108(x83108, x68462, x83110);
  nand n83109(x83109, x83108, x73604);
  nand n83111(x83111, x68462, x83113);
  nand n83112(x83112, x83111, x73609);
  nand n83114(x83114, x68462, x83116);
  nand n83115(x83115, x83114, x73614);
  nand n83117(x83117, x68462, x83119);
  nand n83118(x83118, x83117, x73619);
  nand n83120(x83120, x68462, x83122);
  nand n83121(x83121, x83120, x73624);
  nand n83123(x83123, x68462, x83125);
  nand n83124(x83124, x83123, x73629);
  nand n83126(x83126, x68462, x83128);
  nand n83127(x83127, x83126, x73634);
  nand n83129(x83129, x68462, x83131);
  nand n83130(x83130, x83129, x73639);
  nand n83132(x83132, x68462, x83134);
  nand n83133(x83133, x83132, x73644);
  nand n83135(x83135, x68462, x83137);
  nand n83136(x83136, x83135, x73649);
  nand n83138(x83138, x68462, x83140);
  nand n83139(x83139, x83138, x73654);
  nand n83141(x83141, x68462, x83143);
  nand n83142(x83142, x83141, x73659);
  nand n83144(x83144, x68462, x83146);
  nand n83145(x83145, x83144, x73664);
  nand n83147(x83147, x68462, x83149);
  nand n83148(x83148, x83147, x73669);
  nand n83150(x83150, x68462, x83152);
  nand n83151(x83151, x83150, x73674);
  nand n83153(x83153, x68462, x83155);
  nand n83154(x83154, x83153, x73679);
  nand n83156(x83156, x68462, x83158);
  nand n83157(x83157, x83156, x73684);
  nand n83159(x83159, x68462, x83161);
  nand n83160(x83160, x83159, x73689);
  nand n83162(x83162, x68462, x83164);
  nand n83163(x83163, x83162, x73694);
  nand n83165(x83165, x68462, x83167);
  nand n83166(x83166, x83165, x73699);
  nand n83168(x83168, x68462, x83170);
  nand n83169(x83169, x83168, x73704);
  nand n83171(x83171, x68462, x83173);
  nand n83172(x83172, x83171, x73709);
  nand n83174(x83174, x68462, x83176);
  nand n83175(x83175, x83174, x73714);
  nand n83177(x83177, x68462, x83179);
  nand n83178(x83178, x83177, x73719);
  nand n83180(x83180, x68462, x83182);
  nand n83181(x83181, x83180, x73724);
  nand n83183(x83183, x68462, x83185);
  nand n83184(x83184, x83183, x73729);
  nand n83186(x83186, x68462, x83188);
  nand n83187(x83187, x83186, x73734);
  nand n83189(x83189, x68462, x83191);
  nand n83190(x83190, x83189, x73739);
  nand n83192(x83192, x68462, x83194);
  nand n83193(x83193, x83192, x73744);
  nand n83195(x83195, x68462, x83197);
  nand n83196(x83196, x83195, x73749);
  nand n83198(x83198, x68462, x83200);
  nand n83199(x83199, x83198, x73754);
  nand n83201(x83201, x68462, x83203);
  nand n83202(x83202, x83201, x73759);
  nand n83204(x83204, x68462, x83206);
  nand n83205(x83205, x83204, x73764);
  nand n83207(x83207, x68462, x83209);
  nand n83208(x83208, x83207, x73769);
  nand n83210(x83210, x68462, x83212);
  nand n83211(x83211, x83210, x73774);
  nand n83213(x83213, x68462, x83215);
  nand n83214(x83214, x83213, x73779);
  nand n83216(x83216, x68462, x83218);
  nand n83217(x83217, x83216, x73784);
  nand n83219(x83219, x68462, x83221);
  nand n83220(x83220, x83219, x73789);
  nand n83222(x83222, x68462, x83224);
  nand n83223(x83223, x83222, x73794);
  nand n83225(x83225, x68462, x83227);
  nand n83226(x83226, x83225, x73799);
  nand n83228(x83228, x68462, x83230);
  nand n83229(x83229, x83228, x73804);
  nand n83231(x83231, x68462, x83233);
  nand n83232(x83232, x83231, x73809);
  nand n83234(x83234, x68462, x83236);
  nand n83235(x83235, x83234, x73814);
  nand n83237(x83237, x68462, x83239);
  nand n83238(x83238, x83237, x73819);
  nand n83240(x83240, x68462, x83242);
  nand n83241(x83241, x83240, x73824);
  nand n83243(x83243, x68462, x83245);
  nand n83244(x83244, x83243, x73829);
  nand n83246(x83246, x68462, x83248);
  nand n83247(x83247, x83246, x73834);
  nand n83249(x83249, x68462, x83251);
  nand n83250(x83250, x83249, x73839);
  nand n83252(x83252, x68462, x83254);
  nand n83253(x83253, x83252, x73844);
  nand n83255(x83255, x68462, x83257);
  nand n83256(x83256, x83255, x73849);
  nand n83258(x83258, x68462, x83260);
  nand n83259(x83259, x83258, x73854);
  nand n83261(x83261, x68462, x83263);
  nand n83262(x83262, x83261, x73859);
  nand n83264(x83264, x68462, x83266);
  nand n83265(x83265, x83264, x73864);
  nand n83267(x83267, x68462, x83269);
  nand n83268(x83268, x83267, x73869);
  nand n83270(x83270, x68462, x83272);
  nand n83271(x83271, x83270, x73874);
  nand n83273(x83273, x68462, x83275);
  nand n83274(x83274, x83273, x73879);
  nand n83276(x83276, x68462, x83278);
  nand n83277(x83277, x83276, x73884);
  nand n83279(x83279, x68462, x83281);
  nand n83280(x83280, x83279, x73889);
  nand n83282(x83282, x68462, x83284);
  nand n83283(x83283, x83282, x73894);
  nand n83285(x83285, x68462, x83287);
  nand n83286(x83286, x83285, x73899);
  nand n83288(x83288, x68462, x83290);
  nand n83289(x83289, x83288, x73904);
  nand n83291(x83291, x68462, x83293);
  nand n83292(x83292, x83291, x73909);
  nand n83294(x83294, x68462, x83296);
  nand n83295(x83295, x83294, x73914);
  nand n83297(x83297, x68462, x83299);
  nand n83298(x83298, x83297, x73919);
  nand n83300(x83300, x68462, x83302);
  nand n83301(x83301, x83300, x73924);
  nand n83303(x83303, x68462, x83305);
  nand n83304(x83304, x83303, x73929);
  nand n83306(x83306, x68462, x83308);
  nand n83307(x83307, x83306, x73934);
  nand n83309(x83309, x68462, x83311);
  nand n83310(x83310, x83309, x73939);
  nand n83312(x83312, x68462, x83314);
  nand n83313(x83313, x83312, x73944);
  nand n83315(x83315, x68462, x83317);
  nand n83316(x83316, x83315, x73949);
  nand n83318(x83318, x68462, x83320);
  nand n83319(x83319, x83318, x73954);
  nand n83321(x83321, x68462, x83323);
  nand n83322(x83322, x83321, x73959);
  nand n83324(x83324, x68462, x83326);
  nand n83325(x83325, x83324, x73964);
  nand n83327(x83327, x68462, x83329);
  nand n83328(x83328, x83327, x73969);
  nand n83330(x83330, x68462, x83332);
  nand n83331(x83331, x83330, x73974);
  nand n83333(x83333, x68462, x83335);
  nand n83334(x83334, x83333, x73979);
  nand n83336(x83336, x68462, x83338);
  nand n83337(x83337, x83336, x73984);
  nand n83339(x83339, x68462, x83341);
  nand n83340(x83340, x83339, x73989);
  nand n83342(x83342, x68462, x83344);
  nand n83343(x83343, x83342, x73994);
  nand n83345(x83345, x68462, x83347);
  nand n83346(x83346, x83345, x73999);
  nand n83348(x83348, x71637, x16709);
  nand n83349(x83349, x71135, x87258);
  nand n83350(x83350, x68462, x83352);
  nand n83351(x83351, x83350, x83349);
  nand n83353(x83353, x71637, x16722);
  nand n83354(x83354, x71135, x87259);
  nand n83355(x83355, x68462, x83357);
  nand n83356(x83356, x83355, x83354);
  nand n83358(x83358, x71637, x16729);
  nand n83359(x83359, x71135, x87260);
  nand n83360(x83360, x68462, x83362);
  nand n83361(x83361, x83360, x83359);
  nand n83363(x83363, x71637, x16732);
  nand n83364(x83364, x71135, x87261);
  nand n83365(x83365, x68462, x83367);
  nand n83366(x83366, x83365, x83364);
  nand n83368(x83368, x71637, x16741);
  nand n83369(x83369, x71135, x87262);
  nand n83370(x83370, x68462, x83372);
  nand n83371(x83371, x83370, x83369);
  nand n83373(x83373, x71637, x16744);
  nand n83374(x83374, x71135, x87263);
  nand n83375(x83375, x68462, x83377);
  nand n83376(x83376, x83375, x83374);
  nand n83378(x83378, x71637, x68469);
  nand n83379(x83379, x71135, x87264);
  nand n83380(x83380, x68462, x83382);
  nand n83381(x83381, x83380, x83379);

  not i0(x0, x71142);
  not i1(x1, x71140);
  not i3(x3, x59);
  not i4(x4, x60);
  not i5(x5, x61);
  not i6(x6, x62);
  not i7(x7, x63);
  not i8(x8, x58);
  not i11(x11, x10);
  not i13(x13, x12);
  not i15(x15, x14);
  not i19(x19, x18);
  not i23(x23, x22);
  not i27(x27, x26);
  not i31(x31, x30);
  not i35(x35, x34);
  not i39(x39, x38);
  not i64(x64, x605);
  not i65(x65, x606);
  not i66(x66, x607);
  not i67(x67, x608);
  not i68(x68, x609);
  not i69(x69, x610);
  not i70(x70, x611);
  not i71(x71, x612);
  not i72(x72, x613);
  not i73(x73, x614);
  not i74(x74, x615);
  not i75(x75, x616);
  not i76(x76, x617);
  not i77(x77, x618);
  not i78(x78, x619);
  not i79(x79, x620);
  not i80(x80, x621);
  not i81(x81, x622);
  not i82(x82, x623);
  not i83(x83, x624);
  not i84(x84, x625);
  not i85(x85, x626);
  not i86(x86, x627);
  not i87(x87, x628);
  not i88(x88, x629);
  not i89(x89, x630);
  not i90(x90, x631);
  not i91(x91, x632);
  not i92(x92, x633);
  not i93(x93, x604);
  not i96(x96, x95);
  not i98(x98, x97);
  not i100(x100, x99);
  not i102(x102, x101);
  not i104(x104, x103);
  not i106(x106, x105);
  not i108(x108, x107);
  not i110(x110, x109);
  not i112(x112, x111);
  not i114(x114, x113);
  not i116(x116, x115);
  not i118(x118, x117);
  not i120(x120, x119);
  not i122(x122, x121);
  not i124(x124, x123);
  not i126(x126, x125);
  not i128(x128, x127);
  not i130(x130, x129);
  not i132(x132, x131);
  not i134(x134, x133);
  not i136(x136, x135);
  not i138(x138, x137);
  not i140(x140, x139);
  not i142(x142, x141);
  not i144(x144, x143);
  not i146(x146, x145);
  not i148(x148, x147);
  not i152(x152, x151);
  not i154(x154, x153);
  not i156(x156, x155);
  not i158(x158, x157);
  not i160(x160, x159);
  not i162(x162, x161);
  not i164(x164, x163);
  not i166(x166, x165);
  not i168(x168, x167);
  not i170(x170, x169);
  not i172(x172, x171);
  not i174(x174, x173);
  not i176(x176, x175);
  not i178(x178, x177);
  not i180(x180, x179);
  not i182(x182, x181);
  not i184(x184, x183);
  not i186(x186, x185);
  not i188(x188, x187);
  not i190(x190, x189);
  not i192(x192, x191);
  not i194(x194, x193);
  not i196(x196, x195);
  not i198(x198, x197);
  not i200(x200, x199);
  not i206(x206, x205);
  not i208(x208, x207);
  not i210(x210, x209);
  not i212(x212, x211);
  not i214(x214, x213);
  not i216(x216, x215);
  not i218(x218, x217);
  not i220(x220, x219);
  not i222(x222, x221);
  not i224(x224, x223);
  not i226(x226, x225);
  not i228(x228, x227);
  not i230(x230, x229);
  not i232(x232, x231);
  not i234(x234, x233);
  not i236(x236, x235);
  not i238(x238, x237);
  not i240(x240, x239);
  not i242(x242, x241);
  not i244(x244, x243);
  not i246(x246, x245);
  not i256(x256, x255);
  not i258(x258, x257);
  not i260(x260, x259);
  not i262(x262, x261);
  not i264(x264, x263);
  not i266(x266, x265);
  not i268(x268, x267);
  not i270(x270, x269);
  not i272(x272, x271);
  not i274(x274, x273);
  not i276(x276, x275);
  not i278(x278, x277);
  not i280(x280, x279);
  not i296(x296, x295);
  not i300(x300, x299);
  not i304(x304, x303);
  not i308(x308, x307);
  not i312(x312, x311);
  not i316(x316, x315);
  not i320(x320, x319);
  not i324(x324, x323);
  not i328(x328, x327);
  not i332(x332, x331);
  not i336(x336, x335);
  not i340(x340, x339);
  not i344(x344, x343);
  not i348(x348, x347);
  not i352(x352, x351);
  not i356(x356, x355);
  not i360(x360, x359);
  not i364(x364, x363);
  not i368(x368, x367);
  not i372(x372, x371);
  not i376(x376, x375);
  not i380(x380, x379);
  not i384(x384, x383);
  not i388(x388, x387);
  not i392(x392, x391);
  not i396(x396, x395);
  not i400(x400, x399);
  not i404(x404, x403);
  not i408(x408, x407);
  not i410(x410, x2);
  not i634(x634, x675);
  not i635(x635, x676);
  not i636(x636, x677);
  not i637(x637, x674);
  not i640(x640, x639);
  not i644(x644, x643);
  not i648(x648, x647);
  not i652(x652, x651);
  not i654(x654, x653);
  not i656(x656, x655);
  not i678(x678, x657);
  not i1000(x1000, x71245);
  not i1001(x1001, x71270);
  not i1003(x1003, x1002);
  not i1005(x1005, x1004);
  not i1007(x1007, x1006);
  not i1009(x1009, x1008);
  not i1011(x1011, x71250);
  not i1012(x1012, x71255);
  not i1014(x1014, x1013);
  not i1016(x1016, x1015);
  not i1018(x1018, x1017);
  not i1020(x1020, x1019);
  not i1022(x1022, x71260);
  not i1024(x1024, x1023);
  not i1026(x1026, x1025);
  not i1028(x1028, x1027);
  not i1031(x1031, x1030);
  not i1033(x1033, x1032);
  not i1035(x1035, x1034);
  not i1038(x1038, x71265);
  not i1040(x1040, x1039);
  not i1042(x1042, x1041);
  not i1046(x1046, x1045);
  not i1048(x1048, x1047);
  not i1050(x1050, x1049);
  not i1052(x1052, x1051);
  not i1059(x1059, x1058);
  not i1062(x1062, x1061);
  not i1068(x1068, x1067);
  not i1075(x1075, x1074);
  not i1077(x1077, x1076);
  not i1079(x1079, x1078);
  not i1081(x1081, x1080);
  not i1083(x1083, x1082);
  not i1085(x1085, x1084);
  not i1087(x1087, x1086);
  not i1089(x1089, x1088);
  not i1091(x1091, x1090);
  not i1093(x1093, x1092);
  not i1095(x1095, x1094);
  not i1097(x1097, x1096);
  not i1101(x1101, x1100);
  not i1103(x1103, x1102);
  not i1106(x1106, x1105);
  not i1110(x1110, x1109);
  not i1116(x1116, x1115);
  not i1125(x1125, x1124);
  not i1127(x1127, x1126);
  not i1129(x1129, x1128);
  not i1131(x1131, x1130);
  not i1133(x1133, x1132);
  not i1135(x1135, x1134);
  not i1137(x1137, x1136);
  not i1139(x1139, x1138);
  not i1141(x1141, x1140);
  not i1145(x1145, x1144);
  not i1148(x1148, x1147);
  not i1152(x1152, x1151);
  not i1159(x1159, x1158);
  not i1161(x1161, x1160);
  not i1162(x1162, x1153);
  not i1163(x1163, x1142);
  not i1164(x1164, x1098);
  not i1168(x1168, x1165);
  not i1169(x1169, x1166);
  not i1170(x1170, x1167);
  not i1172(x1172, x1171);
  not i1175(x1175, x1108);
  not i1177(x1177, x1053);
  not i1179(x1179, x1174);
  not i1180(x1180, x1176);
  not i1181(x1181, x1178);
  not i1183(x1183, x1182);
  not i1186(x1186, x1185);
  not i1188(x1188, x1187);
  not i1190(x1190, x1189);
  not i1193(x1193, x1191);
  not i1194(x1194, x1192);
  not i1196(x1196, x70929);
  not i1198(x1198, x1197);
  not i1200(x1200, x1199);
  not i1201(x1201, x70913);
  not i1203(x1203, x1202);
  not i1205(x1205, x1204);
  not i1207(x1207, x1206);
  not i1209(x1209, x1208);
  not i1210(x1210, x70897);
  not i1212(x1212, x1211);
  not i1214(x1214, x1213);
  not i1216(x1216, x1215);
  not i1218(x1218, x1217);
  not i1220(x1220, x1219);
  not i1222(x1222, x1221);
  not i1224(x1224, x1223);
  not i1226(x1226, x1225);
  not i1228(x1228, x1227);
  not i1234(x1234, x1233);
  not i1240(x1240, x1239);
  not i1246(x1246, x1245);
  not i1252(x1252, x1251);
  not i1258(x1258, x1257);
  not i1264(x1264, x1263);
  not i1270(x1270, x1269);
  not i1276(x1276, x1275);
  not i1280(x1280, x1279);
  not i1282(x1282, x1281);
  not i1284(x1284, x1283);
  not i1290(x1290, x1289);
  not i1296(x1296, x1295);
  not i1302(x1302, x1301);
  not i1308(x1308, x1307);
  not i1314(x1314, x1313);
  not i1320(x1320, x1319);
  not i1326(x1326, x1325);
  not i1332(x1332, x1331);
  not i1338(x1338, x1337);
  not i1344(x1344, x1343);
  not i1350(x1350, x1349);
  not i1356(x1356, x1355);
  not i1362(x1362, x1361);
  not i1368(x1368, x1367);
  not i1374(x1374, x1373);
  not i1378(x1378, x1377);
  not i1380(x1380, x1379);
  not i1382(x1382, x1381);
  not i1388(x1388, x1387);
  not i1394(x1394, x1393);
  not i1400(x1400, x1399);
  not i1406(x1406, x1405);
  not i1412(x1412, x1411);
  not i1418(x1418, x1417);
  not i1424(x1424, x71215);
  not i1437(x1437, x71220);
  not i1444(x1444, x71225);
  not i1448(x1448, x71202);
  not i1461(x1461, x71205);
  not i1468(x1468, x71210);
  not i1472(x1472, x71275);
  not i1485(x1485, x71277);
  not i1492(x1492, x71279);
  not i1684(x1684, x1494);
  not i1686(x1686, x1557);
  not i1688(x1688, x1620);
  not i1690(x1690, x1683);
  not i1693(x1693, x1692);
  not i1695(x1695, x1694);
  not i1697(x1697, x1696);
  not i1699(x1699, x1698);
  not i1701(x1701, x1700);
  not i1703(x1703, x1702);
  not i1705(x1705, x1173);
  not i1707(x1707, x1706);
  not i1709(x1709, x1184);
  not i1711(x1711, x1710);
  not i1714(x1714, x1713);
  not i1717(x1717, x1716);
  not i1724(x1724, x1722);
  not i1725(x1725, x1723);
  not i1727(x1727, x71240);
  not i1729(x1729, x1728);
  not i1731(x1731, x1730);
  not i1732(x1732, x71235);
  not i1734(x1734, x1733);
  not i1736(x1736, x1735);
  not i1738(x1738, x1737);
  not i1740(x1740, x1739);
  not i1741(x1741, x71230);
  not i1751(x1751, x1750);
  not i1754(x1754, x1752);
  not i1757(x1757, x1756);
  not i1759(x1759, x1758);
  not i1761(x1761, x1760);
  not i1764(x1764, x1762);
  not i1767(x1767, x1766);
  not i1769(x1769, x1768);
  not i1771(x1771, x1770);
  not i1774(x1774, x1772);
  not i1777(x1777, x1776);
  not i1779(x1779, x1778);
  not i1781(x1781, x1780);
  not i1784(x1784, x1782);
  not i1787(x1787, x1786);
  not i1789(x1789, x1788);
  not i1791(x1791, x1790);
  not i1794(x1794, x1792);
  not i1797(x1797, x1796);
  not i1799(x1799, x1798);
  not i1801(x1801, x1800);
  not i1804(x1804, x1802);
  not i1807(x1807, x1806);
  not i1809(x1809, x1808);
  not i1811(x1811, x1810);
  not i1814(x1814, x1812);
  not i1817(x1817, x1816);
  not i1819(x1819, x1818);
  not i1821(x1821, x1820);
  not i1824(x1824, x1822);
  not i1827(x1827, x1826);
  not i1829(x1829, x1828);
  not i1893(x1893, x1850);
  not i1896(x1896, x1871);
  not i1897(x1897, x1704);
  not i1899(x1899, x1892);
  not i1901(x1901, x1742);
  not i1902(x1902, x1743);
  not i1903(x1903, x1744);
  not i1904(x1904, x1745);
  not i1905(x1905, x1746);
  not i1906(x1906, x1747);
  not i1907(x1907, x1748);
  not i1908(x1908, x1749);
  not i1910(x1910, x1909);
  not i1936(x1936, x1935);
  not i1962(x1962, x1961);
  not i1988(x1988, x1987);
  not i2014(x2014, x2013);
  not i2040(x2040, x2039);
  not i2066(x2066, x2065);
  not i2092(x2092, x2091);
  not i2244(x2244, x2243);
  not i2247(x2247, x2246);
  not i2250(x2250, x2249);
  not i2253(x2253, x2252);
  not i2256(x2256, x2254);
  not i2267(x2267, x2265);
  not i2278(x2278, x2276);
  not i2279(x2279, x2277);
  not i2281(x2281, x70721);
  not i2283(x2283, x2282);
  not i2285(x2285, x2284);
  not i2286(x2286, x70705);
  not i2288(x2288, x2287);
  not i2290(x2290, x2289);
  not i2292(x2292, x2291);
  not i2294(x2294, x2293);
  not i2295(x2295, x70689);
  not i2297(x2297, x2296);
  not i2299(x2299, x2298);
  not i2301(x2301, x2300);
  not i2303(x2303, x2302);
  not i2305(x2305, x2304);
  not i2307(x2307, x2306);
  not i2309(x2309, x2308);
  not i2311(x2311, x2310);
  not i2313(x2313, x2312);
  not i2443(x2443, x2442);
  not i2573(x2573, x2572);
  not i2703(x2703, x2702);
  not i2833(x2833, x2832);
  not i2963(x2963, x2962);
  not i3093(x3093, x3092);
  not i3223(x3223, x3222);
  not i3353(x3353, x3352);
  not i3357(x3357, x3356);
  not i3359(x3359, x3358);
  not i3485(x3485, x3484);
  not i3615(x3615, x3614);
  not i3745(x3745, x3744);
  not i3875(x3875, x3874);
  not i4005(x4005, x4004);
  not i4135(x4135, x4134);
  not i4265(x4265, x4264);
  not i4395(x4395, x4394);
  not i4403(x4403, x4402);
  not i4405(x4405, x4404);
  not i4527(x4527, x4526);
  not i4657(x4657, x4656);
  not i4787(x4787, x4786);
  not i4917(x4917, x4916);
  not i5047(x5047, x5046);
  not i5177(x5177, x5176);
  not i5307(x5307, x5306);
  not i5437(x5437, x5436);
  not i5441(x5441, x5440);
  not i5443(x5443, x5442);
  not i5447(x5447, x5446);
  not i5449(x5449, x5448);
  not i5571(x5571, x5570);
  not i5701(x5701, x5700);
  not i5831(x5831, x5830);
  not i5961(x5961, x5960);
  not i6091(x6091, x6090);
  not i6221(x6221, x6220);
  not i6351(x6351, x6350);
  not i6481(x6481, x2258);
  not i6494(x6494, x2261);
  not i6501(x6501, x2264);
  not i7156(x7156, x2269);
  not i7169(x7169, x2272);
  not i7176(x7176, x2275);
  not i14555(x14555, x14554);
  not i14557(x14557, x14556);
  not i14560(x14560, x14559);
  not i14567(x14567, x14565);
  not i14568(x14568, x14566);
  not i14571(x14571, x14570);
  not i14573(x14573, x14572);
  not i14575(x14575, x14574);
  not i14577(x14577, x14576);
  not i14579(x14579, x14578);
  not i14581(x14581, x14580);
  not i14591(x14591, x14590);
  not i14594(x14594, x14592);
  not i14597(x14597, x14596);
  not i14599(x14599, x14598);
  not i14601(x14601, x14600);
  not i14604(x14604, x14602);
  not i14607(x14607, x14606);
  not i14609(x14609, x14608);
  not i14611(x14611, x14610);
  not i14614(x14614, x14612);
  not i14617(x14617, x14616);
  not i14619(x14619, x14618);
  not i14621(x14621, x14620);
  not i14624(x14624, x14622);
  not i14627(x14627, x14626);
  not i14629(x14629, x14628);
  not i14631(x14631, x14630);
  not i14634(x14634, x14632);
  not i14637(x14637, x14636);
  not i14639(x14639, x14638);
  not i14641(x14641, x14640);
  not i14644(x14644, x14642);
  not i14647(x14647, x14646);
  not i14649(x14649, x14648);
  not i14651(x14651, x14650);
  not i14654(x14654, x14652);
  not i14657(x14657, x14656);
  not i14659(x14659, x14658);
  not i14661(x14661, x14660);
  not i14664(x14664, x14662);
  not i14667(x14667, x14666);
  not i14669(x14669, x14668);
  not i14733(x14733, x14690);
  not i14735(x14735, x14734);
  not i14737(x14737, x14736);
  not i14739(x14739, x14738);
  not i14741(x14741, x14740);
  not i14743(x14743, x14742);
  not i14746(x14746, x14711);
  not i14748(x14748, x14747);
  not i14751(x14751, x14732);
  not i14752(x14752, x2248);
  not i14754(x14754, x14582);
  not i14755(x14755, x14583);
  not i14756(x14756, x14584);
  not i14757(x14757, x14585);
  not i14758(x14758, x14586);
  not i14759(x14759, x14587);
  not i14760(x14760, x14588);
  not i14761(x14761, x14589);
  not i14763(x14763, x14762);
  not i14789(x14789, x14788);
  not i14815(x14815, x14814);
  not i14841(x14841, x14840);
  not i14867(x14867, x14866);
  not i14893(x14893, x14892);
  not i14919(x14919, x14918);
  not i14945(x14945, x14944);
  not i15096(x15096, x14551);
  not i15152(x15152, x15151);
  not i15217(x15217, x15216);
  not i15219(x15219, x15218);
  not i15222(x15222, x15221);
  not i15224(x15224, x15223);
  not i15227(x15227, x15226);
  not i15229(x15229, x15228);
  not i15231(x15231, x15155);
  not i15232(x15232, x71289);
  not i15236(x15236, x15158);
  not i15237(x15237, x71294);
  not i15240(x15240, x15239);
  not i15242(x15242, x15161);
  not i15243(x15243, x71299);
  not i15246(x15246, x15245);
  not i15248(x15248, x15164);
  not i15249(x15249, x71304);
  not i15252(x15252, x15251);
  not i15254(x15254, x15167);
  not i15255(x15255, x71309);
  not i15258(x15258, x15257);
  not i15260(x15260, x15170);
  not i15261(x15261, x71314);
  not i15264(x15264, x15263);
  not i15266(x15266, x15173);
  not i15267(x15267, x71319);
  not i15270(x15270, x15269);
  not i15272(x15272, x15176);
  not i15273(x15273, x71324);
  not i15276(x15276, x15275);
  not i15278(x15278, x15179);
  not i15279(x15279, x71329);
  not i15282(x15282, x15281);
  not i15284(x15284, x15182);
  not i15285(x15285, x71334);
  not i15288(x15288, x15287);
  not i15290(x15290, x15185);
  not i15291(x15291, x71339);
  not i15294(x15294, x15293);
  not i15296(x15296, x15188);
  not i15297(x15297, x71344);
  not i15300(x15300, x15299);
  not i15302(x15302, x15191);
  not i15303(x15303, x71349);
  not i15306(x15306, x15305);
  not i15308(x15308, x15194);
  not i15309(x15309, x71354);
  not i15312(x15312, x15311);
  not i15314(x15314, x15197);
  not i15315(x15315, x71359);
  not i15318(x15318, x15317);
  not i15320(x15320, x15200);
  not i15321(x15321, x71364);
  not i15324(x15324, x15323);
  not i15326(x15326, x15203);
  not i15327(x15327, x71369);
  not i15330(x15330, x15329);
  not i15332(x15332, x15206);
  not i15333(x15333, x71374);
  not i15336(x15336, x15335);
  not i15338(x15338, x15209);
  not i15339(x15339, x71379);
  not i15342(x15342, x15341);
  not i15344(x15344, x15211);
  not i15345(x15345, x71384);
  not i15348(x15348, x15347);
  not i15350(x15350, x15213);
  not i15351(x15351, x71389);
  not i15354(x15354, x15353);
  not i15356(x15356, x15215);
  not i15357(x15357, x71394);
  not i15360(x15360, x15359);
  not i15362(x15362, x71399);
  not i15365(x15365, x15364);
  not i15367(x15367, x71404);
  not i15370(x15370, x15369);
  not i15372(x15372, x71409);
  not i15375(x15375, x15374);
  not i15377(x15377, x71414);
  not i15380(x15380, x15379);
  not i15382(x15382, x71419);
  not i15385(x15385, x15384);
  not i15387(x15387, x71424);
  not i15390(x15390, x15389);
  not i15392(x15392, x71429);
  not i15395(x15395, x15394);
  not i15397(x15397, x71434);
  not i15400(x15400, x15399);
  not i15402(x15402, x71439);
  not i15405(x15405, x15404);
  not i15407(x15407, x71444);
  not i15410(x15410, x15409);
  not i15411(x15411, x15230);
  not i15412(x15412, x15235);
  not i15413(x15413, x15241);
  not i15414(x15414, x15247);
  not i15415(x15415, x15253);
  not i15416(x15416, x15259);
  not i15417(x15417, x15265);
  not i15418(x15418, x15271);
  not i15419(x15419, x15277);
  not i15420(x15420, x15283);
  not i15421(x15421, x15289);
  not i15422(x15422, x15295);
  not i15423(x15423, x15301);
  not i15424(x15424, x15307);
  not i15425(x15425, x15313);
  not i15426(x15426, x15319);
  not i15427(x15427, x15325);
  not i15428(x15428, x15331);
  not i15429(x15429, x15337);
  not i15430(x15430, x15343);
  not i15431(x15431, x15349);
  not i15432(x15432, x15355);
  not i15433(x15433, x15361);
  not i15434(x15434, x15366);
  not i15435(x15435, x15371);
  not i15436(x15436, x15376);
  not i15437(x15437, x15381);
  not i15438(x15438, x15386);
  not i15439(x15439, x15391);
  not i15440(x15440, x15396);
  not i15446(x15446, x15445);
  not i15450(x15450, x15449);
  not i15454(x15454, x15453);
  not i15458(x15458, x15457);
  not i15462(x15462, x15461);
  not i15466(x15466, x15465);
  not i15470(x15470, x15469);
  not i15474(x15474, x15473);
  not i15478(x15478, x15477);
  not i15482(x15482, x15481);
  not i15486(x15486, x15485);
  not i15490(x15490, x15489);
  not i15494(x15494, x15493);
  not i15498(x15498, x15497);
  not i15502(x15502, x15501);
  not i15506(x15506, x15505);
  not i15510(x15510, x15509);
  not i15514(x15514, x15513);
  not i15518(x15518, x15517);
  not i15522(x15522, x15521);
  not i15526(x15526, x15525);
  not i15530(x15530, x15529);
  not i15534(x15534, x15533);
  not i15538(x15538, x15537);
  not i15542(x15542, x15541);
  not i15546(x15546, x15545);
  not i15550(x15550, x15549);
  not i15554(x15554, x15553);
  not i15558(x15558, x15557);
  not i15559(x15559, x15442);
  not i15561(x15561, x15444);
  not i15564(x15564, x15448);
  not i15567(x15567, x15452);
  not i15570(x15570, x15569);
  not i15572(x15572, x15456);
  not i15575(x15575, x15574);
  not i15577(x15577, x15460);
  not i15580(x15580, x15579);
  not i15582(x15582, x15464);
  not i15585(x15585, x15584);
  not i15587(x15587, x15468);
  not i15590(x15590, x15589);
  not i15592(x15592, x15472);
  not i15595(x15595, x15594);
  not i15597(x15597, x15476);
  not i15600(x15600, x15599);
  not i15602(x15602, x15480);
  not i15605(x15605, x15604);
  not i15607(x15607, x15484);
  not i15610(x15610, x15609);
  not i15612(x15612, x15488);
  not i15615(x15615, x15614);
  not i15617(x15617, x15492);
  not i15620(x15620, x15619);
  not i15622(x15622, x15496);
  not i15625(x15625, x15624);
  not i15627(x15627, x15500);
  not i15630(x15630, x15629);
  not i15632(x15632, x15504);
  not i15635(x15635, x15634);
  not i15637(x15637, x15508);
  not i15640(x15640, x15639);
  not i15642(x15642, x15512);
  not i15645(x15645, x15644);
  not i15647(x15647, x15516);
  not i15650(x15650, x15649);
  not i15652(x15652, x15520);
  not i15655(x15655, x15654);
  not i15657(x15657, x15524);
  not i15660(x15660, x15659);
  not i15662(x15662, x15528);
  not i15665(x15665, x15664);
  not i15667(x15667, x15532);
  not i15670(x15670, x15669);
  not i15672(x15672, x15536);
  not i15675(x15675, x15674);
  not i15677(x15677, x15540);
  not i15680(x15680, x15679);
  not i15682(x15682, x15544);
  not i15685(x15685, x15684);
  not i15687(x15687, x15548);
  not i15690(x15690, x15689);
  not i15692(x15692, x15552);
  not i15695(x15695, x15694);
  not i15697(x15697, x15556);
  not i15700(x15700, x15699);
  not i15701(x15701, x15565);
  not i15703(x15703, x15568);
  not i15706(x15706, x15573);
  not i15709(x15709, x15578);
  not i15712(x15712, x15583);
  not i15715(x15715, x15588);
  not i15718(x15718, x15717);
  not i15720(x15720, x15593);
  not i15723(x15723, x15722);
  not i15725(x15725, x15598);
  not i15728(x15728, x15727);
  not i15730(x15730, x15603);
  not i15733(x15733, x15732);
  not i15735(x15735, x15608);
  not i15738(x15738, x15737);
  not i15740(x15740, x15613);
  not i15743(x15743, x15742);
  not i15745(x15745, x15618);
  not i15748(x15748, x15747);
  not i15750(x15750, x15623);
  not i15753(x15753, x15752);
  not i15755(x15755, x15628);
  not i15758(x15758, x15757);
  not i15760(x15760, x15633);
  not i15763(x15763, x15762);
  not i15765(x15765, x15638);
  not i15768(x15768, x15767);
  not i15770(x15770, x15643);
  not i15773(x15773, x15772);
  not i15775(x15775, x15648);
  not i15778(x15778, x15777);
  not i15780(x15780, x15653);
  not i15783(x15783, x15782);
  not i15785(x15785, x15658);
  not i15788(x15788, x15787);
  not i15790(x15790, x15663);
  not i15793(x15793, x15792);
  not i15795(x15795, x15668);
  not i15798(x15798, x15797);
  not i15800(x15800, x15673);
  not i15803(x15803, x15802);
  not i15805(x15805, x15678);
  not i15808(x15808, x15807);
  not i15810(x15810, x15683);
  not i15813(x15813, x15812);
  not i15815(x15815, x15688);
  not i15818(x15818, x15817);
  not i15820(x15820, x15693);
  not i15823(x15823, x15822);
  not i15825(x15825, x15698);
  not i15828(x15828, x15827);
  not i15829(x15829, x15713);
  not i15831(x15831, x15716);
  not i15834(x15834, x15721);
  not i15837(x15837, x15726);
  not i15840(x15840, x15731);
  not i15843(x15843, x15736);
  not i15846(x15846, x15741);
  not i15849(x15849, x15746);
  not i15852(x15852, x15751);
  not i15855(x15855, x15756);
  not i15858(x15858, x15857);
  not i15860(x15860, x15761);
  not i15863(x15863, x15862);
  not i15865(x15865, x15766);
  not i15868(x15868, x15867);
  not i15870(x15870, x15771);
  not i15873(x15873, x15872);
  not i15875(x15875, x15776);
  not i15878(x15878, x15877);
  not i15880(x15880, x15781);
  not i15883(x15883, x15882);
  not i15885(x15885, x15786);
  not i15888(x15888, x15887);
  not i15890(x15890, x15791);
  not i15893(x15893, x15892);
  not i15895(x15895, x15796);
  not i15898(x15898, x15897);
  not i15900(x15900, x15801);
  not i15903(x15903, x15902);
  not i15905(x15905, x15806);
  not i15908(x15908, x15907);
  not i15910(x15910, x15811);
  not i15913(x15913, x15912);
  not i15915(x15915, x15816);
  not i15918(x15918, x15917);
  not i15920(x15920, x15821);
  not i15923(x15923, x15922);
  not i15925(x15925, x15826);
  not i15928(x15928, x15927);
  not i15929(x15929, x15853);
  not i15931(x15931, x15856);
  not i15934(x15934, x15861);
  not i15937(x15937, x15866);
  not i15940(x15940, x15871);
  not i15943(x15943, x15876);
  not i15946(x15946, x15881);
  not i15949(x15949, x15886);
  not i15952(x15952, x15891);
  not i15955(x15955, x15896);
  not i15958(x15958, x15901);
  not i15961(x15961, x15906);
  not i15964(x15964, x15911);
  not i15967(x15967, x15916);
  not i15970(x15970, x15921);
  not i15973(x15973, x15926);
  not i15980(x15980, x15979);
  not i15982(x15982, x15562);
  not i15989(x15989, x15704);
  not i15993(x15993, x15707);
  not i15997(x15997, x15710);
  not i16004(x16004, x15832);
  not i16008(x16008, x15835);
  not i16012(x16012, x15838);
  not i16016(x16016, x15841);
  not i16020(x16020, x15844);
  not i16024(x16024, x15847);
  not i16028(x16028, x15850);
  not i16035(x16035, x15932);
  not i16039(x16039, x15935);
  not i16043(x16043, x15938);
  not i16047(x16047, x15941);
  not i16051(x16051, x15944);
  not i16055(x16055, x15947);
  not i16059(x16059, x15950);
  not i16063(x16063, x15953);
  not i16067(x16067, x15956);
  not i16071(x16071, x15959);
  not i16075(x16075, x15962);
  not i16079(x16079, x15965);
  not i16083(x16083, x15968);
  not i16087(x16087, x15971);
  not i16091(x16091, x15974);
  not i16096(x16096, x16095);
  not i16098(x16098, x16097);
  not i16100(x16100, x16099);
  not i16102(x16102, x16101);
  not i16104(x16104, x16103);
  not i16106(x16106, x16105);
  not i16108(x16108, x16107);
  not i16110(x16110, x16109);
  not i16112(x16112, x16111);
  not i16114(x16114, x16113);
  not i16116(x16116, x16115);
  not i16118(x16118, x16117);
  not i16120(x16120, x16119);
  not i16122(x16122, x16121);
  not i16124(x16124, x16123);
  not i16126(x16126, x16125);
  not i16128(x16128, x16127);
  not i16130(x16130, x16129);
  not i16132(x16132, x16131);
  not i16134(x16134, x16133);
  not i16136(x16136, x16135);
  not i16138(x16138, x16137);
  not i16140(x16140, x16139);
  not i16142(x16142, x16141);
  not i16144(x16144, x16143);
  not i16146(x16146, x16145);
  not i16148(x16148, x16147);
  not i16152(x16152, x16151);
  not i16154(x16154, x16153);
  not i16156(x16156, x16155);
  not i16158(x16158, x16157);
  not i16160(x16160, x16159);
  not i16162(x16162, x16161);
  not i16164(x16164, x16163);
  not i16166(x16166, x16165);
  not i16168(x16168, x16167);
  not i16170(x16170, x16169);
  not i16172(x16172, x16171);
  not i16174(x16174, x16173);
  not i16176(x16176, x16175);
  not i16178(x16178, x16177);
  not i16180(x16180, x16179);
  not i16182(x16182, x16181);
  not i16184(x16184, x16183);
  not i16186(x16186, x16185);
  not i16188(x16188, x16187);
  not i16190(x16190, x16189);
  not i16192(x16192, x16191);
  not i16194(x16194, x16193);
  not i16196(x16196, x16195);
  not i16198(x16198, x16197);
  not i16200(x16200, x16199);
  not i16206(x16206, x16205);
  not i16208(x16208, x16207);
  not i16210(x16210, x16209);
  not i16212(x16212, x16211);
  not i16214(x16214, x16213);
  not i16216(x16216, x16215);
  not i16218(x16218, x16217);
  not i16220(x16220, x16219);
  not i16222(x16222, x16221);
  not i16224(x16224, x16223);
  not i16226(x16226, x16225);
  not i16228(x16228, x16227);
  not i16230(x16230, x16229);
  not i16232(x16232, x16231);
  not i16234(x16234, x16233);
  not i16236(x16236, x16235);
  not i16238(x16238, x16237);
  not i16240(x16240, x16239);
  not i16242(x16242, x16241);
  not i16244(x16244, x16243);
  not i16246(x16246, x16245);
  not i16256(x16256, x16255);
  not i16258(x16258, x16257);
  not i16260(x16260, x16259);
  not i16262(x16262, x16261);
  not i16264(x16264, x16263);
  not i16266(x16266, x16265);
  not i16268(x16268, x16267);
  not i16270(x16270, x16269);
  not i16272(x16272, x16271);
  not i16274(x16274, x16273);
  not i16276(x16276, x16275);
  not i16278(x16278, x16277);
  not i16280(x16280, x16279);
  not i16296(x16296, x16295);
  not i16300(x16300, x16299);
  not i16304(x16304, x16303);
  not i16308(x16308, x16307);
  not i16312(x16312, x16311);
  not i16316(x16316, x16315);
  not i16320(x16320, x16319);
  not i16324(x16324, x16323);
  not i16328(x16328, x16327);
  not i16332(x16332, x16331);
  not i16336(x16336, x16335);
  not i16340(x16340, x16339);
  not i16344(x16344, x16343);
  not i16348(x16348, x16347);
  not i16352(x16352, x16351);
  not i16356(x16356, x16355);
  not i16360(x16360, x16359);
  not i16364(x16364, x16363);
  not i16368(x16368, x16367);
  not i16372(x16372, x16371);
  not i16376(x16376, x16375);
  not i16380(x16380, x16379);
  not i16384(x16384, x16383);
  not i16388(x16388, x16387);
  not i16392(x16392, x16391);
  not i16396(x16396, x16395);
  not i16400(x16400, x16399);
  not i16404(x16404, x16403);
  not i16408(x16408, x16407);
  not i16410(x16410, x15220);
  not i16508(x16508, x16506);
  not i16509(x16509, x16507);
  not i16512(x16512, x16511);
  not i16514(x16514, x16513);
  not i16516(x16516, x16515);
  not i16518(x16518, x16517);
  not i16520(x16520, x16519);
  not i16522(x16522, x16521);
  not i16524(x16524, x16523);
  not i16526(x16526, x16525);
  not i16528(x16528, x16527);
  not i16530(x16530, x16529);
  not i16532(x16532, x16531);
  not i16534(x16534, x16533);
  not i16536(x16536, x16535);
  not i16538(x16538, x16537);
  not i16540(x16540, x16539);
  not i16542(x16542, x16541);
  not i16544(x16544, x16543);
  not i16546(x16546, x16545);
  not i16548(x16548, x16547);
  not i16550(x16550, x16549);
  not i16552(x16552, x16551);
  not i16554(x16554, x16553);
  not i16556(x16556, x16555);
  not i16558(x16558, x16557);
  not i16560(x16560, x16559);
  not i16562(x16562, x16561);
  not i16564(x16564, x16563);
  not i16566(x16566, x16565);
  not i16568(x16568, x16567);
  not i16570(x16570, x16569);
  not i16572(x16572, x16571);
  not i16574(x16574, x16573);
  not i16576(x16576, x16575);
  not i16578(x16578, x16577);
  not i16580(x16580, x16579);
  not i16582(x16582, x16581);
  not i16584(x16584, x16583);
  not i16586(x16586, x16585);
  not i16588(x16588, x16587);
  not i16590(x16590, x16589);
  not i16592(x16592, x16591);
  not i16594(x16594, x16593);
  not i16596(x16596, x16595);
  not i16598(x16598, x16597);
  not i16600(x16600, x16599);
  not i16602(x16602, x16601);
  not i16604(x16604, x16603);
  not i16606(x16606, x16605);
  not i16608(x16608, x16607);
  not i16610(x16610, x16609);
  not i16612(x16612, x16611);
  not i16658(x16658, x16657);
  not i16659(x16659, x16656);
  not i16661(x16661, x16655);
  not i16662(x16662, x16654);
  not i16664(x16664, x16660);
  not i16665(x16665, x16663);
  not i16667(x16667, x16666);
  not i16679(x16679, x16670);
  not i16680(x16680, x16669);
  not i16682(x16682, x16672);
  not i16683(x16683, x16671);
  not i16685(x16685, x16674);
  not i16686(x16686, x16673);
  not i16688(x16688, x16676);
  not i16689(x16689, x16675);
  not i16691(x16691, x16678);
  not i16692(x16692, x16677);
  not i16694(x16694, x16684);
  not i16695(x16695, x16681);
  not i16697(x16697, x16690);
  not i16698(x16698, x16687);
  not i16700(x16700, x16693);
  not i16702(x16702, x16699);
  not i16703(x16703, x16696);
  not i16705(x16705, x16701);
  not i16706(x16706, x16704);
  not i16709(x16709, x16708);
  not i16713(x16713, x16711);
  not i16714(x16714, x16710);
  not i16716(x16716, x16712);
  not i16718(x16718, x16717);
  not i16719(x16719, x16715);
  not i16722(x16722, x16721);
  not i16725(x16725, x16724);
  not i16726(x16726, x16723);
  not i16729(x16729, x16728);
  not i16732(x16732, x16731);
  not i16735(x16735, x16734);
  not i16736(x16736, x16733);
  not i16738(x16738, x16737);
  not i16741(x16741, x16740);
  not i16744(x16744, x16743);
  not i16745(x16745, x68738);
  not i16747(x16747, x71942);
  not i16843(x16843, x16749);
  not i16844(x16844, x16752);
  not i16845(x16845, x16755);
  not i16846(x16846, x16758);
  not i16847(x16847, x16761);
  not i16848(x16848, x16764);
  not i16849(x16849, x16767);
  not i16850(x16850, x16770);
  not i16851(x16851, x16773);
  not i16852(x16852, x16776);
  not i16853(x16853, x16779);
  not i16854(x16854, x16782);
  not i16855(x16855, x16785);
  not i16856(x16856, x16788);
  not i16857(x16857, x16791);
  not i16858(x16858, x16794);
  not i16859(x16859, x16797);
  not i16860(x16860, x16800);
  not i16861(x16861, x16803);
  not i16862(x16862, x16806);
  not i16863(x16863, x16809);
  not i16864(x16864, x16812);
  not i16865(x16865, x16815);
  not i16866(x16866, x16818);
  not i16867(x16867, x16821);
  not i16868(x16868, x16824);
  not i16869(x16869, x16827);
  not i16870(x16870, x16830);
  not i16871(x16871, x16833);
  not i16872(x16872, x16836);
  not i16873(x16873, x16839);
  not i16874(x16874, x16842);
  not i16876(x16876, x71977);
  not i16973(x16973, x16878);
  not i16974(x16974, x72047);
  not i16977(x16977, x16976);
  not i16979(x16979, x16881);
  not i16980(x16980, x72052);
  not i16983(x16983, x16982);
  not i16985(x16985, x16884);
  not i16986(x16986, x72057);
  not i16989(x16989, x16988);
  not i16991(x16991, x16887);
  not i16992(x16992, x72062);
  not i16995(x16995, x16994);
  not i16997(x16997, x16890);
  not i16998(x16998, x72067);
  not i17001(x17001, x17000);
  not i17003(x17003, x16893);
  not i17004(x17004, x72072);
  not i17007(x17007, x17006);
  not i17009(x17009, x16896);
  not i17010(x17010, x72077);
  not i17013(x17013, x17012);
  not i17015(x17015, x16899);
  not i17016(x17016, x72082);
  not i17019(x17019, x17018);
  not i17021(x17021, x16902);
  not i17022(x17022, x72087);
  not i17025(x17025, x17024);
  not i17027(x17027, x16905);
  not i17028(x17028, x72092);
  not i17031(x17031, x17030);
  not i17033(x17033, x16908);
  not i17034(x17034, x72097);
  not i17037(x17037, x17036);
  not i17039(x17039, x16911);
  not i17040(x17040, x72102);
  not i17043(x17043, x17042);
  not i17045(x17045, x16914);
  not i17046(x17046, x72107);
  not i17049(x17049, x17048);
  not i17051(x17051, x16917);
  not i17052(x17052, x72112);
  not i17055(x17055, x17054);
  not i17057(x17057, x16920);
  not i17058(x17058, x72117);
  not i17061(x17061, x17060);
  not i17063(x17063, x16923);
  not i17064(x17064, x72122);
  not i17067(x17067, x17066);
  not i17069(x17069, x16926);
  not i17070(x17070, x72127);
  not i17073(x17073, x17072);
  not i17075(x17075, x16929);
  not i17076(x17076, x72132);
  not i17079(x17079, x17078);
  not i17081(x17081, x16932);
  not i17082(x17082, x72137);
  not i17085(x17085, x17084);
  not i17087(x17087, x16935);
  not i17088(x17088, x72142);
  not i17091(x17091, x17090);
  not i17093(x17093, x16938);
  not i17094(x17094, x72147);
  not i17097(x17097, x17096);
  not i17099(x17099, x16941);
  not i17100(x17100, x72152);
  not i17103(x17103, x17102);
  not i17105(x17105, x16944);
  not i17106(x17106, x72157);
  not i17109(x17109, x17108);
  not i17111(x17111, x16947);
  not i17112(x17112, x72162);
  not i17115(x17115, x17114);
  not i17117(x17117, x16950);
  not i17118(x17118, x72167);
  not i17121(x17121, x17120);
  not i17123(x17123, x16953);
  not i17124(x17124, x72172);
  not i17127(x17127, x17126);
  not i17129(x17129, x16956);
  not i17130(x17130, x72177);
  not i17133(x17133, x17132);
  not i17135(x17135, x16959);
  not i17136(x17136, x72182);
  not i17139(x17139, x17138);
  not i17141(x17141, x16962);
  not i17142(x17142, x72187);
  not i17145(x17145, x17144);
  not i17147(x17147, x16965);
  not i17148(x17148, x72192);
  not i17151(x17151, x17150);
  not i17153(x17153, x16968);
  not i17154(x17154, x72197);
  not i17157(x17157, x17156);
  not i17159(x17159, x16971);
  not i17160(x17160, x72202);
  not i17163(x17163, x17162);
  not i17164(x17164, x16972);
  not i17165(x17165, x16978);
  not i17166(x17166, x16984);
  not i17167(x17167, x16990);
  not i17168(x17168, x16996);
  not i17169(x17169, x17002);
  not i17170(x17170, x17008);
  not i17171(x17171, x17014);
  not i17172(x17172, x17020);
  not i17173(x17173, x17026);
  not i17174(x17174, x17032);
  not i17175(x17175, x17038);
  not i17176(x17176, x17044);
  not i17177(x17177, x17050);
  not i17178(x17178, x17056);
  not i17179(x17179, x17062);
  not i17180(x17180, x17068);
  not i17181(x17181, x17074);
  not i17182(x17182, x17080);
  not i17183(x17183, x17086);
  not i17184(x17184, x17092);
  not i17185(x17185, x17098);
  not i17186(x17186, x17104);
  not i17187(x17187, x17110);
  not i17188(x17188, x17116);
  not i17189(x17189, x17122);
  not i17190(x17190, x17128);
  not i17191(x17191, x17134);
  not i17192(x17192, x17140);
  not i17193(x17193, x17146);
  not i17199(x17199, x17198);
  not i17203(x17203, x17202);
  not i17207(x17207, x17206);
  not i17211(x17211, x17210);
  not i17215(x17215, x17214);
  not i17219(x17219, x17218);
  not i17223(x17223, x17222);
  not i17227(x17227, x17226);
  not i17231(x17231, x17230);
  not i17235(x17235, x17234);
  not i17239(x17239, x17238);
  not i17243(x17243, x17242);
  not i17247(x17247, x17246);
  not i17251(x17251, x17250);
  not i17255(x17255, x17254);
  not i17259(x17259, x17258);
  not i17263(x17263, x17262);
  not i17267(x17267, x17266);
  not i17271(x17271, x17270);
  not i17275(x17275, x17274);
  not i17279(x17279, x17278);
  not i17283(x17283, x17282);
  not i17287(x17287, x17286);
  not i17291(x17291, x17290);
  not i17295(x17295, x17294);
  not i17299(x17299, x17298);
  not i17303(x17303, x17302);
  not i17307(x17307, x17306);
  not i17311(x17311, x17310);
  not i17315(x17315, x17314);
  not i17317(x17317, x17197);
  not i17320(x17320, x17201);
  not i17323(x17323, x17205);
  not i17326(x17326, x17325);
  not i17328(x17328, x17209);
  not i17331(x17331, x17330);
  not i17333(x17333, x17213);
  not i17336(x17336, x17335);
  not i17338(x17338, x17217);
  not i17341(x17341, x17340);
  not i17343(x17343, x17221);
  not i17346(x17346, x17345);
  not i17348(x17348, x17225);
  not i17351(x17351, x17350);
  not i17353(x17353, x17229);
  not i17356(x17356, x17355);
  not i17358(x17358, x17233);
  not i17361(x17361, x17360);
  not i17363(x17363, x17237);
  not i17366(x17366, x17365);
  not i17368(x17368, x17241);
  not i17371(x17371, x17370);
  not i17373(x17373, x17245);
  not i17376(x17376, x17375);
  not i17378(x17378, x17249);
  not i17381(x17381, x17380);
  not i17383(x17383, x17253);
  not i17386(x17386, x17385);
  not i17388(x17388, x17257);
  not i17391(x17391, x17390);
  not i17393(x17393, x17261);
  not i17396(x17396, x17395);
  not i17398(x17398, x17265);
  not i17401(x17401, x17400);
  not i17403(x17403, x17269);
  not i17406(x17406, x17405);
  not i17408(x17408, x17273);
  not i17411(x17411, x17410);
  not i17413(x17413, x17277);
  not i17416(x17416, x17415);
  not i17418(x17418, x17281);
  not i17421(x17421, x17420);
  not i17423(x17423, x17285);
  not i17426(x17426, x17425);
  not i17428(x17428, x17289);
  not i17431(x17431, x17430);
  not i17433(x17433, x17293);
  not i17436(x17436, x17435);
  not i17438(x17438, x17297);
  not i17441(x17441, x17440);
  not i17443(x17443, x17301);
  not i17446(x17446, x17445);
  not i17448(x17448, x17305);
  not i17451(x17451, x17450);
  not i17453(x17453, x17309);
  not i17456(x17456, x17455);
  not i17458(x17458, x17313);
  not i17461(x17461, x17460);
  not i17463(x17463, x17324);
  not i17466(x17466, x17329);
  not i17469(x17469, x17334);
  not i17472(x17472, x17339);
  not i17475(x17475, x17344);
  not i17478(x17478, x17477);
  not i17480(x17480, x17349);
  not i17483(x17483, x17482);
  not i17485(x17485, x17354);
  not i17488(x17488, x17487);
  not i17490(x17490, x17359);
  not i17493(x17493, x17492);
  not i17495(x17495, x17364);
  not i17498(x17498, x17497);
  not i17500(x17500, x17369);
  not i17503(x17503, x17502);
  not i17505(x17505, x17374);
  not i17508(x17508, x17507);
  not i17510(x17510, x17379);
  not i17513(x17513, x17512);
  not i17515(x17515, x17384);
  not i17518(x17518, x17517);
  not i17520(x17520, x17389);
  not i17523(x17523, x17522);
  not i17525(x17525, x17394);
  not i17528(x17528, x17527);
  not i17530(x17530, x17399);
  not i17533(x17533, x17532);
  not i17535(x17535, x17404);
  not i17538(x17538, x17537);
  not i17540(x17540, x17409);
  not i17543(x17543, x17542);
  not i17545(x17545, x17414);
  not i17548(x17548, x17547);
  not i17550(x17550, x17419);
  not i17553(x17553, x17552);
  not i17555(x17555, x17424);
  not i17558(x17558, x17557);
  not i17560(x17560, x17429);
  not i17563(x17563, x17562);
  not i17565(x17565, x17434);
  not i17568(x17568, x17567);
  not i17570(x17570, x17439);
  not i17573(x17573, x17572);
  not i17575(x17575, x17444);
  not i17578(x17578, x17577);
  not i17580(x17580, x17449);
  not i17583(x17583, x17582);
  not i17585(x17585, x17454);
  not i17588(x17588, x17587);
  not i17590(x17590, x17459);
  not i17593(x17593, x17592);
  not i17595(x17595, x17476);
  not i17598(x17598, x17481);
  not i17601(x17601, x17486);
  not i17604(x17604, x17491);
  not i17607(x17607, x17496);
  not i17610(x17610, x17501);
  not i17613(x17613, x17506);
  not i17616(x17616, x17511);
  not i17619(x17619, x17516);
  not i17622(x17622, x17621);
  not i17624(x17624, x17521);
  not i17627(x17627, x17626);
  not i17629(x17629, x17526);
  not i17632(x17632, x17631);
  not i17634(x17634, x17531);
  not i17637(x17637, x17636);
  not i17639(x17639, x17536);
  not i17642(x17642, x17641);
  not i17644(x17644, x17541);
  not i17647(x17647, x17646);
  not i17649(x17649, x17546);
  not i17652(x17652, x17651);
  not i17654(x17654, x17551);
  not i17657(x17657, x17656);
  not i17659(x17659, x17556);
  not i17662(x17662, x17661);
  not i17664(x17664, x17561);
  not i17667(x17667, x17666);
  not i17669(x17669, x17566);
  not i17672(x17672, x17671);
  not i17674(x17674, x17571);
  not i17677(x17677, x17676);
  not i17679(x17679, x17576);
  not i17682(x17682, x17681);
  not i17684(x17684, x17581);
  not i17687(x17687, x17686);
  not i17689(x17689, x17586);
  not i17692(x17692, x17691);
  not i17694(x17694, x17591);
  not i17697(x17697, x17696);
  not i17699(x17699, x17620);
  not i17702(x17702, x17625);
  not i17705(x17705, x17630);
  not i17708(x17708, x17635);
  not i17711(x17711, x17640);
  not i17714(x17714, x17645);
  not i17717(x17717, x17650);
  not i17720(x17720, x17655);
  not i17723(x17723, x17660);
  not i17726(x17726, x17665);
  not i17729(x17729, x17670);
  not i17732(x17732, x17675);
  not i17735(x17735, x17680);
  not i17738(x17738, x17685);
  not i17741(x17741, x17690);
  not i17744(x17744, x17695);
  not i17748(x17748, x17747);
  not i17750(x17750, x17195);
  not i17753(x17753, x17752);
  not i17755(x17755, x17318);
  not i17758(x17758, x17757);
  not i17760(x17760, x17321);
  not i17763(x17763, x17762);
  not i17765(x17765, x17464);
  not i17768(x17768, x17767);
  not i17770(x17770, x17467);
  not i17773(x17773, x17772);
  not i17775(x17775, x17470);
  not i17778(x17778, x17777);
  not i17780(x17780, x17473);
  not i17783(x17783, x17782);
  not i17785(x17785, x17596);
  not i17788(x17788, x17787);
  not i17790(x17790, x17599);
  not i17793(x17793, x17792);
  not i17795(x17795, x17602);
  not i17798(x17798, x17797);
  not i17800(x17800, x17605);
  not i17803(x17803, x17802);
  not i17805(x17805, x17608);
  not i17808(x17808, x17807);
  not i17810(x17810, x17611);
  not i17813(x17813, x17812);
  not i17815(x17815, x17614);
  not i17818(x17818, x17817);
  not i17820(x17820, x17617);
  not i17823(x17823, x17822);
  not i17825(x17825, x17700);
  not i17828(x17828, x17827);
  not i17830(x17830, x17703);
  not i17833(x17833, x17832);
  not i17835(x17835, x17706);
  not i17838(x17838, x17837);
  not i17840(x17840, x17709);
  not i17843(x17843, x17842);
  not i17845(x17845, x17712);
  not i17848(x17848, x17847);
  not i17850(x17850, x17715);
  not i17853(x17853, x17852);
  not i17855(x17855, x17718);
  not i17858(x17858, x17857);
  not i17860(x17860, x17721);
  not i17863(x17863, x17862);
  not i17865(x17865, x17724);
  not i17868(x17868, x17867);
  not i17870(x17870, x17727);
  not i17873(x17873, x17872);
  not i17875(x17875, x17730);
  not i17878(x17878, x17877);
  not i17880(x17880, x17733);
  not i17883(x17883, x17882);
  not i17885(x17885, x17736);
  not i17888(x17888, x17887);
  not i17890(x17890, x17739);
  not i17893(x17893, x17892);
  not i17895(x17895, x17742);
  not i17898(x17898, x17897);
  not i17900(x17900, x17745);
  not i17903(x17903, x17902);
  not i17906(x17906, x17905);
  not i17908(x17908, x17907);
  not i17910(x17910, x17909);
  not i17912(x17912, x17911);
  not i17914(x17914, x17913);
  not i17916(x17916, x17915);
  not i17918(x17918, x17917);
  not i17920(x17920, x17919);
  not i17923(x17923, x17922);
  not i17925(x17925, x17924);
  not i17927(x17927, x17926);
  not i17929(x17929, x17928);
  not i17931(x17931, x17930);
  not i17933(x17933, x17932);
  not i17935(x17935, x17934);
  not i17937(x17937, x17936);
  not i17939(x17939, x17938);
  not i17941(x17941, x17940);
  not i17943(x17943, x17942);
  not i17945(x17945, x17944);
  not i17947(x17947, x17946);
  not i17949(x17949, x17948);
  not i17951(x17951, x17950);
  not i17953(x17953, x17952);
  not i17955(x17955, x17954);
  not i17958(x17958, x17957);
  not i17960(x17960, x17959);
  not i17962(x17962, x17961);
  not i17964(x17964, x17963);
  not i17966(x17966, x17965);
  not i17968(x17968, x17967);
  not i17970(x17970, x17969);
  not i17972(x17972, x17971);
  not i17974(x17974, x17973);
  not i17976(x17976, x17975);
  not i17978(x17978, x17977);
  not i17980(x17980, x17979);
  not i17982(x17982, x17981);
  not i17984(x17984, x17983);
  not i17986(x17986, x17985);
  not i17988(x17988, x17987);
  not i17990(x17990, x17989);
  not i17992(x17992, x17991);
  not i17994(x17994, x17993);
  not i17996(x17996, x17995);
  not i17998(x17998, x17997);
  not i18000(x18000, x17999);
  not i18002(x18002, x18001);
  not i18004(x18004, x18003);
  not i18006(x18006, x18005);
  not i18008(x18008, x18007);
  not i18011(x18011, x18010);
  not i18013(x18013, x18012);
  not i18015(x18015, x18014);
  not i18017(x18017, x18016);
  not i18019(x18019, x18018);
  not i18021(x18021, x18020);
  not i18023(x18023, x18022);
  not i18025(x18025, x18024);
  not i18027(x18027, x18026);
  not i18029(x18029, x18028);
  not i18031(x18031, x18030);
  not i18033(x18033, x18032);
  not i18035(x18035, x18034);
  not i18037(x18037, x18036);
  not i18039(x18039, x18038);
  not i18041(x18041, x18040);
  not i18043(x18043, x18042);
  not i18045(x18045, x18044);
  not i18047(x18047, x18046);
  not i18049(x18049, x18048);
  not i18051(x18051, x18050);
  not i18053(x18053, x18052);
  not i18055(x18055, x18054);
  not i18057(x18057, x18056);
  not i18059(x18059, x18058);
  not i18061(x18061, x18060);
  not i18063(x18063, x18062);
  not i18065(x18065, x18064);
  not i18067(x18067, x18066);
  not i18069(x18069, x18068);
  not i18071(x18071, x18070);
  not i18073(x18073, x18072);
  not i18075(x18075, x18074);
  not i18077(x18077, x18076);
  not i18079(x18079, x18078);
  not i18082(x18082, x18081);
  not i18084(x18084, x18083);
  not i18086(x18086, x18085);
  not i18088(x18088, x18087);
  not i18090(x18090, x18089);
  not i18092(x18092, x18091);
  not i18094(x18094, x18093);
  not i18096(x18096, x18095);
  not i18098(x18098, x18097);
  not i18100(x18100, x18099);
  not i18102(x18102, x18101);
  not i18104(x18104, x18103);
  not i18106(x18106, x18105);
  not i18108(x18108, x18107);
  not i18110(x18110, x18109);
  not i18112(x18112, x18111);
  not i18114(x18114, x18113);
  not i18116(x18116, x18115);
  not i18118(x18118, x18117);
  not i18120(x18120, x18119);
  not i18122(x18122, x18121);
  not i18124(x18124, x18123);
  not i18126(x18126, x18125);
  not i18128(x18128, x18127);
  not i18130(x18130, x18129);
  not i18132(x18132, x18131);
  not i18134(x18134, x18133);
  not i18136(x18136, x18135);
  not i18138(x18138, x18137);
  not i18140(x18140, x18139);
  not i18142(x18142, x18141);
  not i18144(x18144, x18143);
  not i18146(x18146, x18145);
  not i18148(x18148, x18147);
  not i18150(x18150, x18149);
  not i18152(x18152, x18151);
  not i18154(x18154, x18153);
  not i18156(x18156, x18155);
  not i18158(x18158, x18157);
  not i18160(x18160, x18159);
  not i18162(x18162, x18161);
  not i18164(x18164, x18163);
  not i18166(x18166, x18165);
  not i18168(x18168, x18167);
  not i18171(x18171, x18170);
  not i18173(x18173, x18172);
  not i18175(x18175, x18174);
  not i18177(x18177, x18176);
  not i18179(x18179, x18178);
  not i18181(x18181, x18180);
  not i18183(x18183, x18182);
  not i18185(x18185, x18184);
  not i18187(x18187, x18186);
  not i18189(x18189, x18188);
  not i18191(x18191, x18190);
  not i18193(x18193, x18192);
  not i18195(x18195, x18194);
  not i18197(x18197, x18196);
  not i18199(x18199, x18198);
  not i18201(x18201, x18200);
  not i18203(x18203, x18202);
  not i18205(x18205, x18204);
  not i18207(x18207, x18206);
  not i18209(x18209, x18208);
  not i18211(x18211, x18210);
  not i18213(x18213, x18212);
  not i18215(x18215, x18214);
  not i18217(x18217, x18216);
  not i18219(x18219, x18218);
  not i18221(x18221, x18220);
  not i18223(x18223, x18222);
  not i18225(x18225, x18224);
  not i18227(x18227, x18226);
  not i18229(x18229, x18228);
  not i18231(x18231, x18230);
  not i18233(x18233, x18232);
  not i18235(x18235, x18234);
  not i18237(x18237, x18236);
  not i18239(x18239, x18238);
  not i18241(x18241, x18240);
  not i18243(x18243, x18242);
  not i18245(x18245, x18244);
  not i18247(x18247, x18246);
  not i18249(x18249, x18248);
  not i18251(x18251, x18250);
  not i18253(x18253, x18252);
  not i18255(x18255, x18254);
  not i18257(x18257, x18256);
  not i18259(x18259, x18258);
  not i18261(x18261, x18260);
  not i18263(x18263, x18262);
  not i18265(x18265, x18264);
  not i18267(x18267, x18266);
  not i18269(x18269, x18268);
  not i18271(x18271, x18270);
  not i18273(x18273, x18272);
  not i18275(x18275, x18274);
  not i18278(x18278, x18277);
  not i18280(x18280, x18279);
  not i18282(x18282, x18281);
  not i18284(x18284, x18283);
  not i18286(x18286, x18285);
  not i18288(x18288, x18287);
  not i18290(x18290, x18289);
  not i18292(x18292, x18291);
  not i18294(x18294, x18293);
  not i18296(x18296, x18295);
  not i18298(x18298, x18297);
  not i18300(x18300, x18299);
  not i18302(x18302, x18301);
  not i18304(x18304, x18303);
  not i18306(x18306, x18305);
  not i18308(x18308, x18307);
  not i18310(x18310, x18309);
  not i18312(x18312, x18311);
  not i18314(x18314, x18313);
  not i18316(x18316, x18315);
  not i18318(x18318, x18317);
  not i18320(x18320, x18319);
  not i18322(x18322, x18321);
  not i18324(x18324, x18323);
  not i18326(x18326, x18325);
  not i18328(x18328, x18327);
  not i18330(x18330, x18329);
  not i18332(x18332, x18331);
  not i18334(x18334, x18333);
  not i18336(x18336, x18335);
  not i18338(x18338, x18337);
  not i18340(x18340, x18339);
  not i18342(x18342, x18341);
  not i18344(x18344, x18343);
  not i18346(x18346, x18345);
  not i18348(x18348, x18347);
  not i18350(x18350, x18349);
  not i18352(x18352, x18351);
  not i18354(x18354, x18353);
  not i18356(x18356, x18355);
  not i18358(x18358, x18357);
  not i18360(x18360, x18359);
  not i18362(x18362, x18361);
  not i18364(x18364, x18363);
  not i18366(x18366, x18365);
  not i18368(x18368, x18367);
  not i18370(x18370, x18369);
  not i18372(x18372, x18371);
  not i18374(x18374, x18373);
  not i18376(x18376, x18375);
  not i18378(x18378, x18377);
  not i18380(x18380, x18379);
  not i18382(x18382, x18381);
  not i18384(x18384, x18383);
  not i18386(x18386, x18385);
  not i18388(x18388, x18387);
  not i18390(x18390, x18389);
  not i18392(x18392, x18391);
  not i18394(x18394, x18393);
  not i18396(x18396, x18395);
  not i18398(x18398, x18397);
  not i18400(x18400, x18399);
  not i18403(x18403, x18402);
  not i18405(x18405, x18404);
  not i18407(x18407, x18406);
  not i18409(x18409, x18408);
  not i18411(x18411, x18410);
  not i18413(x18413, x18412);
  not i18415(x18415, x18414);
  not i18417(x18417, x18416);
  not i18419(x18419, x18418);
  not i18421(x18421, x18420);
  not i18423(x18423, x18422);
  not i18425(x18425, x18424);
  not i18427(x18427, x18426);
  not i18429(x18429, x18428);
  not i18431(x18431, x18430);
  not i18433(x18433, x18432);
  not i18435(x18435, x18434);
  not i18437(x18437, x18436);
  not i18439(x18439, x18438);
  not i18441(x18441, x18440);
  not i18443(x18443, x18442);
  not i18445(x18445, x18444);
  not i18447(x18447, x18446);
  not i18449(x18449, x18448);
  not i18451(x18451, x18450);
  not i18453(x18453, x18452);
  not i18455(x18455, x18454);
  not i18457(x18457, x18456);
  not i18459(x18459, x18458);
  not i18461(x18461, x18460);
  not i18463(x18463, x18462);
  not i18465(x18465, x18464);
  not i18467(x18467, x18466);
  not i18469(x18469, x18468);
  not i18471(x18471, x18470);
  not i18473(x18473, x18472);
  not i18475(x18475, x18474);
  not i18477(x18477, x18476);
  not i18479(x18479, x18478);
  not i18481(x18481, x18480);
  not i18483(x18483, x18482);
  not i18485(x18485, x18484);
  not i18487(x18487, x18486);
  not i18489(x18489, x18488);
  not i18491(x18491, x18490);
  not i18493(x18493, x18492);
  not i18495(x18495, x18494);
  not i18497(x18497, x18496);
  not i18499(x18499, x18498);
  not i18501(x18501, x18500);
  not i18503(x18503, x18502);
  not i18505(x18505, x18504);
  not i18507(x18507, x18506);
  not i18509(x18509, x18508);
  not i18511(x18511, x18510);
  not i18513(x18513, x18512);
  not i18515(x18515, x18514);
  not i18517(x18517, x18516);
  not i18519(x18519, x18518);
  not i18521(x18521, x18520);
  not i18523(x18523, x18522);
  not i18525(x18525, x18524);
  not i18527(x18527, x18526);
  not i18529(x18529, x18528);
  not i18531(x18531, x18530);
  not i18533(x18533, x18532);
  not i18535(x18535, x18534);
  not i18537(x18537, x18536);
  not i18539(x18539, x18538);
  not i18541(x18541, x18540);
  not i18543(x18543, x18542);
  not i18546(x18546, x18545);
  not i18548(x18548, x18547);
  not i18550(x18550, x18549);
  not i18552(x18552, x18551);
  not i18554(x18554, x18553);
  not i18556(x18556, x18555);
  not i18558(x18558, x18557);
  not i18560(x18560, x18559);
  not i18562(x18562, x18561);
  not i18564(x18564, x18563);
  not i18566(x18566, x18565);
  not i18568(x18568, x18567);
  not i18570(x18570, x18569);
  not i18572(x18572, x18571);
  not i18574(x18574, x18573);
  not i18576(x18576, x18575);
  not i18578(x18578, x18577);
  not i18580(x18580, x18579);
  not i18582(x18582, x18581);
  not i18584(x18584, x18583);
  not i18586(x18586, x18585);
  not i18588(x18588, x18587);
  not i18590(x18590, x18589);
  not i18592(x18592, x18591);
  not i18594(x18594, x18593);
  not i18596(x18596, x18595);
  not i18598(x18598, x18597);
  not i18600(x18600, x18599);
  not i18602(x18602, x18601);
  not i18604(x18604, x18603);
  not i18606(x18606, x18605);
  not i18608(x18608, x18607);
  not i18610(x18610, x18609);
  not i18612(x18612, x18611);
  not i18614(x18614, x18613);
  not i18616(x18616, x18615);
  not i18618(x18618, x18617);
  not i18620(x18620, x18619);
  not i18622(x18622, x18621);
  not i18624(x18624, x18623);
  not i18626(x18626, x18625);
  not i18628(x18628, x18627);
  not i18630(x18630, x18629);
  not i18632(x18632, x18631);
  not i18634(x18634, x18633);
  not i18636(x18636, x18635);
  not i18638(x18638, x18637);
  not i18640(x18640, x18639);
  not i18642(x18642, x18641);
  not i18644(x18644, x18643);
  not i18646(x18646, x18645);
  not i18648(x18648, x18647);
  not i18650(x18650, x18649);
  not i18652(x18652, x18651);
  not i18654(x18654, x18653);
  not i18656(x18656, x18655);
  not i18658(x18658, x18657);
  not i18660(x18660, x18659);
  not i18662(x18662, x18661);
  not i18664(x18664, x18663);
  not i18666(x18666, x18665);
  not i18668(x18668, x18667);
  not i18670(x18670, x18669);
  not i18672(x18672, x18671);
  not i18674(x18674, x18673);
  not i18676(x18676, x18675);
  not i18678(x18678, x18677);
  not i18680(x18680, x18679);
  not i18682(x18682, x18681);
  not i18684(x18684, x18683);
  not i18686(x18686, x18685);
  not i18688(x18688, x18687);
  not i18690(x18690, x18689);
  not i18692(x18692, x18691);
  not i18694(x18694, x18693);
  not i18696(x18696, x18695);
  not i18698(x18698, x18697);
  not i18700(x18700, x18699);
  not i18702(x18702, x18701);
  not i18704(x18704, x18703);
  not i18707(x18707, x18706);
  not i18709(x18709, x18708);
  not i18711(x18711, x18710);
  not i18713(x18713, x18712);
  not i18715(x18715, x18714);
  not i18717(x18717, x18716);
  not i18719(x18719, x18718);
  not i18721(x18721, x18720);
  not i18723(x18723, x18722);
  not i18725(x18725, x18724);
  not i18727(x18727, x18726);
  not i18729(x18729, x18728);
  not i18731(x18731, x18730);
  not i18733(x18733, x18732);
  not i18735(x18735, x18734);
  not i18737(x18737, x18736);
  not i18739(x18739, x18738);
  not i18741(x18741, x18740);
  not i18743(x18743, x18742);
  not i18745(x18745, x18744);
  not i18747(x18747, x18746);
  not i18749(x18749, x18748);
  not i18751(x18751, x18750);
  not i18753(x18753, x18752);
  not i18755(x18755, x18754);
  not i18757(x18757, x18756);
  not i18759(x18759, x18758);
  not i18761(x18761, x18760);
  not i18763(x18763, x18762);
  not i18765(x18765, x18764);
  not i18767(x18767, x18766);
  not i18769(x18769, x18768);
  not i18771(x18771, x18770);
  not i18773(x18773, x18772);
  not i18775(x18775, x18774);
  not i18777(x18777, x18776);
  not i18779(x18779, x18778);
  not i18781(x18781, x18780);
  not i18783(x18783, x18782);
  not i18785(x18785, x18784);
  not i18787(x18787, x18786);
  not i18789(x18789, x18788);
  not i18791(x18791, x18790);
  not i18793(x18793, x18792);
  not i18795(x18795, x18794);
  not i18797(x18797, x18796);
  not i18799(x18799, x18798);
  not i18801(x18801, x18800);
  not i18803(x18803, x18802);
  not i18805(x18805, x18804);
  not i18807(x18807, x18806);
  not i18809(x18809, x18808);
  not i18811(x18811, x18810);
  not i18813(x18813, x18812);
  not i18815(x18815, x18814);
  not i18817(x18817, x18816);
  not i18819(x18819, x18818);
  not i18821(x18821, x18820);
  not i18823(x18823, x18822);
  not i18825(x18825, x18824);
  not i18827(x18827, x18826);
  not i18829(x18829, x18828);
  not i18831(x18831, x18830);
  not i18833(x18833, x18832);
  not i18835(x18835, x18834);
  not i18837(x18837, x18836);
  not i18839(x18839, x18838);
  not i18841(x18841, x18840);
  not i18843(x18843, x18842);
  not i18845(x18845, x18844);
  not i18847(x18847, x18846);
  not i18849(x18849, x18848);
  not i18851(x18851, x18850);
  not i18853(x18853, x18852);
  not i18855(x18855, x18854);
  not i18857(x18857, x18856);
  not i18859(x18859, x18858);
  not i18861(x18861, x18860);
  not i18863(x18863, x18862);
  not i18865(x18865, x18864);
  not i18867(x18867, x18866);
  not i18869(x18869, x18868);
  not i18871(x18871, x18870);
  not i18873(x18873, x18872);
  not i18875(x18875, x18874);
  not i18877(x18877, x18876);
  not i18879(x18879, x18878);
  not i18881(x18881, x18880);
  not i18883(x18883, x18882);
  not i18886(x18886, x18885);
  not i18888(x18888, x18887);
  not i18890(x18890, x18889);
  not i18892(x18892, x18891);
  not i18894(x18894, x18893);
  not i18896(x18896, x18895);
  not i18898(x18898, x18897);
  not i18900(x18900, x18899);
  not i18902(x18902, x18901);
  not i18904(x18904, x18903);
  not i18906(x18906, x18905);
  not i18908(x18908, x18907);
  not i18910(x18910, x18909);
  not i18912(x18912, x18911);
  not i18914(x18914, x18913);
  not i18916(x18916, x18915);
  not i18918(x18918, x18917);
  not i18920(x18920, x18919);
  not i18922(x18922, x18921);
  not i18924(x18924, x18923);
  not i18926(x18926, x18925);
  not i18928(x18928, x18927);
  not i18930(x18930, x18929);
  not i18932(x18932, x18931);
  not i18934(x18934, x18933);
  not i18936(x18936, x18935);
  not i18938(x18938, x18937);
  not i18940(x18940, x18939);
  not i18942(x18942, x18941);
  not i18944(x18944, x18943);
  not i18946(x18946, x18945);
  not i18948(x18948, x18947);
  not i18955(x18955, x18954);
  not i18963(x18963, x18962);
  not i18971(x18971, x18970);
  not i18982(x18982, x18981);
  not i18990(x18990, x18989);
  not i18998(x18998, x18997);
  not i19006(x19006, x19005);
  not i19010(x19010, x19009);
  not i19015(x19015, x19014);
  not i19023(x19023, x19022);
  not i19027(x19027, x19026);
  not i19035(x19035, x19034);
  not i19043(x19043, x19042);
  not i19047(x19047, x19046);
  not i19052(x19052, x19051);
  not i19056(x19056, x19055);
  not i19061(x19061, x19060);
  not i19069(x19069, x19068);
  not i19073(x19073, x19072);
  not i19078(x19078, x19077);
  not i19082(x19082, x19081);
  not i19087(x19087, x19086);
  not i19095(x19095, x19094);
  not i19099(x19099, x19098);
  not i19104(x19104, x19103);
  not i19108(x19108, x19107);
  not i19116(x19116, x19115);
  not i19124(x19124, x19123);
  not i19128(x19128, x19127);
  not i19133(x19133, x19132);
  not i19137(x19137, x19136);
  not i19142(x19142, x19141);
  not i19146(x19146, x19145);
  not i19151(x19151, x19150);
  not i19159(x19159, x19158);
  not i19163(x19163, x19162);
  not i19168(x19168, x19167);
  not i19172(x19172, x19171);
  not i19177(x19177, x19176);
  not i19181(x19181, x19180);
  not i19186(x19186, x19185);
  not i19194(x19194, x19193);
  not i19198(x19198, x19197);
  not i19203(x19203, x19202);
  not i19207(x19207, x19206);
  not i19212(x19212, x19211);
  not i19216(x19216, x19215);
  not i19224(x19224, x19223);
  not i19232(x19232, x19231);
  not i19236(x19236, x19235);
  not i19241(x19241, x19240);
  not i19245(x19245, x19244);
  not i19250(x19250, x19249);
  not i19254(x19254, x19253);
  not i19259(x19259, x19258);
  not i19267(x19267, x19266);
  not i19275(x19275, x19274);
  not i19279(x19279, x19278);
  not i19284(x19284, x19283);
  not i19288(x19288, x19287);
  not i19293(x19293, x19292);
  not i19297(x19297, x19296);
  not i19302(x19302, x19301);
  not i19306(x19306, x19305);
  not i19311(x19311, x19310);
  not i19319(x19319, x19318);
  not i19323(x19323, x19322);
  not i19328(x19328, x19327);
  not i19332(x19332, x19331);
  not i19337(x19337, x19336);
  not i19341(x19341, x19340);
  not i19346(x19346, x19345);
  not i19350(x19350, x19349);
  not i19358(x19358, x19357);
  not i19366(x19366, x19365);
  not i19370(x19370, x19369);
  not i19375(x19375, x19374);
  not i19379(x19379, x19378);
  not i19384(x19384, x19383);
  not i19388(x19388, x19387);
  not i19393(x19393, x19392);
  not i19397(x19397, x19396);
  not i19402(x19402, x19401);
  not i19406(x19406, x19405);
  not i19411(x19411, x19410);
  not i19419(x19419, x19418);
  not i19423(x19423, x19422);
  not i19428(x19428, x19427);
  not i19432(x19432, x19431);
  not i19437(x19437, x19436);
  not i19441(x19441, x19440);
  not i19446(x19446, x19445);
  not i19450(x19450, x19449);
  not i19455(x19455, x19454);
  not i19459(x19459, x19458);
  not i19464(x19464, x19463);
  not i19472(x19472, x19471);
  not i19476(x19476, x19475);
  not i19481(x19481, x19480);
  not i19485(x19485, x19484);
  not i19490(x19490, x19489);
  not i19494(x19494, x19493);
  not i19499(x19499, x19498);
  not i19503(x19503, x19502);
  not i19508(x19508, x19507);
  not i19512(x19512, x19511);
  not i19520(x19520, x19519);
  not i19528(x19528, x19527);
  not i19532(x19532, x19531);
  not i19537(x19537, x19536);
  not i19541(x19541, x19540);
  not i19546(x19546, x19545);
  not i19550(x19550, x19549);
  not i19555(x19555, x19554);
  not i19559(x19559, x19558);
  not i19564(x19564, x19563);
  not i19568(x19568, x19567);
  not i19573(x19573, x19572);
  not i19577(x19577, x19576);
  not i19582(x19582, x19581);
  not i19590(x19590, x19589);
  not i19594(x19594, x19593);
  not i19599(x19599, x19598);
  not i19603(x19603, x19602);
  not i19608(x19608, x19607);
  not i19612(x19612, x19611);
  not i19617(x19617, x19616);
  not i19621(x19621, x19620);
  not i19626(x19626, x19625);
  not i19630(x19630, x19629);
  not i19635(x19635, x19634);
  not i19639(x19639, x19638);
  not i19644(x19644, x19643);
  not i19652(x19652, x19651);
  not i19656(x19656, x19655);
  not i19661(x19661, x19660);
  not i19665(x19665, x19664);
  not i19670(x19670, x19669);
  not i19674(x19674, x19673);
  not i19679(x19679, x19678);
  not i19683(x19683, x19682);
  not i19688(x19688, x19687);
  not i19692(x19692, x19691);
  not i19697(x19697, x19696);
  not i19701(x19701, x19700);
  not i19709(x19709, x19708);
  not i19717(x19717, x19716);
  not i19721(x19721, x19720);
  not i19726(x19726, x19725);
  not i19730(x19730, x19729);
  not i19735(x19735, x19734);
  not i19739(x19739, x19738);
  not i19744(x19744, x19743);
  not i19748(x19748, x19747);
  not i19753(x19753, x19752);
  not i19757(x19757, x19756);
  not i19762(x19762, x19761);
  not i19766(x19766, x19765);
  not i19771(x19771, x19770);
  not i19779(x19779, x19778);
  not i19787(x19787, x19786);
  not i19791(x19791, x19790);
  not i19796(x19796, x19795);
  not i19800(x19800, x19799);
  not i19805(x19805, x19804);
  not i19809(x19809, x19808);
  not i19814(x19814, x19813);
  not i19818(x19818, x19817);
  not i19823(x19823, x19822);
  not i19827(x19827, x19826);
  not i19832(x19832, x19831);
  not i19836(x19836, x19835);
  not i19841(x19841, x19840);
  not i19845(x19845, x19844);
  not i19850(x19850, x19849);
  not i19858(x19858, x19857);
  not i19862(x19862, x19861);
  not i19867(x19867, x19866);
  not i19871(x19871, x19870);
  not i19876(x19876, x19875);
  not i19880(x19880, x19879);
  not i19885(x19885, x19884);
  not i19889(x19889, x19888);
  not i19894(x19894, x19893);
  not i19898(x19898, x19897);
  not i19903(x19903, x19902);
  not i19907(x19907, x19906);
  not i19912(x19912, x19911);
  not i19916(x19916, x19915);
  not i19924(x19924, x19923);
  not i19932(x19932, x19931);
  not i19936(x19936, x19935);
  not i19941(x19941, x19940);
  not i19945(x19945, x19944);
  not i19950(x19950, x19949);
  not i19954(x19954, x19953);
  not i19959(x19959, x19958);
  not i19963(x19963, x19962);
  not i19968(x19968, x19967);
  not i19972(x19972, x19971);
  not i19977(x19977, x19976);
  not i19981(x19981, x19980);
  not i19986(x19986, x19985);
  not i19990(x19990, x19989);
  not i19995(x19995, x19994);
  not i19999(x19999, x19998);
  not i20004(x20004, x20003);
  not i20012(x20012, x20011);
  not i20016(x20016, x20015);
  not i20021(x20021, x20020);
  not i20025(x20025, x20024);
  not i20030(x20030, x20029);
  not i20034(x20034, x20033);
  not i20039(x20039, x20038);
  not i20043(x20043, x20042);
  not i20048(x20048, x20047);
  not i20052(x20052, x20051);
  not i20057(x20057, x20056);
  not i20061(x20061, x20060);
  not i20066(x20066, x20065);
  not i20070(x20070, x20069);
  not i20075(x20075, x20074);
  not i20079(x20079, x20078);
  not i20084(x20084, x20083);
  not i20092(x20092, x20091);
  not i20096(x20096, x20095);
  not i20101(x20101, x20100);
  not i20105(x20105, x20104);
  not i20110(x20110, x20109);
  not i20114(x20114, x20113);
  not i20119(x20119, x20118);
  not i20123(x20123, x20122);
  not i20128(x20128, x20127);
  not i20132(x20132, x20131);
  not i20137(x20137, x20136);
  not i20141(x20141, x20140);
  not i20146(x20146, x20145);
  not i20150(x20150, x20149);
  not i20155(x20155, x20154);
  not i20159(x20159, x20158);
  not i20167(x20167, x20166);
  not i20171(x20171, x20170);
  not i20176(x20176, x20175);
  not i20180(x20180, x20179);
  not i20185(x20185, x20184);
  not i20189(x20189, x20188);
  not i20194(x20194, x20193);
  not i20198(x20198, x20197);
  not i20203(x20203, x20202);
  not i20207(x20207, x20206);
  not i20212(x20212, x20211);
  not i20216(x20216, x20215);
  not i20221(x20221, x20220);
  not i20225(x20225, x20224);
  not i20230(x20230, x20229);
  not i20234(x20234, x20233);
  not i20239(x20239, x20238);
  not i20243(x20243, x20242);
  not i20248(x20248, x20247);
  not i20252(x20252, x20251);
  not i20257(x20257, x20256);
  not i20261(x20261, x20260);
  not i20266(x20266, x20265);
  not i20270(x20270, x20269);
  not i20275(x20275, x20274);
  not i20279(x20279, x20278);
  not i20284(x20284, x20283);
  not i20288(x20288, x20287);
  not i20293(x20293, x20292);
  not i20297(x20297, x20296);
  not i20302(x20302, x20301);
  not i20306(x20306, x20305);
  not i20311(x20311, x20310);
  not i20315(x20315, x20314);
  not i20320(x20320, x20319);
  not i20324(x20324, x20323);
  not i20329(x20329, x20328);
  not i20333(x20333, x20332);
  not i20338(x20338, x20337);
  not i20342(x20342, x20341);
  not i20347(x20347, x20346);
  not i20351(x20351, x20350);
  not i20355(x20355, x20354);
  not i20359(x20359, x20358);
  not i20363(x20363, x20362);
  not i20367(x20367, x20366);
  not i20371(x20371, x20370);
  not i20375(x20375, x20374);
  not i20379(x20379, x20378);
  not i20383(x20383, x20382);
  not i20387(x20387, x20386);
  not i20391(x20391, x20390);
  not i20395(x20395, x20394);
  not i20399(x20399, x20398);
  not i20403(x20403, x20402);
  not i20407(x20407, x20406);
  not i20411(x20411, x20410);
  not i20415(x20415, x20414);
  not i20419(x20419, x20418);
  not i20423(x20423, x20422);
  not i20427(x20427, x20426);
  not i20428(x20428, x18959);
  not i20429(x20429, x18967);
  not i20431(x20431, x18975);
  not i20435(x20435, x18994);
  not i20436(x20436, x18986);
  not i20443(x20443, x19011);
  not i20444(x20444, x19002);
  not i20451(x20451, x19028);
  not i20452(x20452, x19019);
  not i20455(x20455, x20454);
  not i20464(x20464, x19048);
  not i20465(x20465, x19039);
  not i20468(x20468, x20467);
  not i20470(x20470, x19057);
  not i20477(x20477, x20476);
  not i20481(x20481, x20480);
  not i20484(x20484, x19074);
  not i20485(x20485, x19065);
  not i20488(x20488, x20487);
  not i20490(x20490, x19083);
  not i20497(x20497, x20496);
  not i20501(x20501, x20500);
  not i20504(x20504, x19100);
  not i20505(x20505, x19091);
  not i20508(x20508, x20507);
  not i20510(x20510, x19109);
  not i20517(x20517, x20516);
  not i20521(x20521, x20520);
  not i20524(x20524, x19129);
  not i20525(x20525, x19120);
  not i20528(x20528, x20527);
  not i20530(x20530, x19138);
  not i20534(x20534, x19147);
  not i20538(x20538, x20537);
  not i20542(x20542, x20541);
  not i20545(x20545, x19164);
  not i20546(x20546, x19155);
  not i20549(x20549, x20548);
  not i20551(x20551, x19173);
  not i20555(x20555, x19182);
  not i20559(x20559, x20558);
  not i20563(x20563, x20562);
  not i20566(x20566, x19199);
  not i20567(x20567, x19190);
  not i20570(x20570, x20569);
  not i20572(x20572, x19208);
  not i20577(x20577, x19217);
  not i20583(x20583, x20582);
  not i20587(x20587, x20586);
  not i20590(x20590, x19237);
  not i20591(x20591, x19228);
  not i20594(x20594, x20593);
  not i20596(x20596, x19246);
  not i20601(x20601, x19263);
  not i20602(x20602, x19255);
  not i20608(x20608, x20607);
  not i20612(x20612, x20611);
  not i20618(x20618, x19280);
  not i20619(x20619, x19271);
  not i20622(x20622, x20621);
  not i20624(x20624, x19289);
  not i20629(x20629, x19307);
  not i20630(x20630, x19298);
  not i20636(x20636, x20635);
  not i20640(x20640, x20639);
  not i20646(x20646, x19324);
  not i20647(x20647, x19315);
  not i20650(x20650, x20649);
  not i20652(x20652, x19333);
  not i20657(x20657, x19351);
  not i20658(x20658, x19342);
  not i20661(x20661, x20660);
  not i20665(x20665, x20664);
  not i20670(x20670, x20669);
  not i20674(x20674, x20673);
  not i20680(x20680, x19371);
  not i20681(x20681, x19362);
  not i20684(x20684, x20683);
  not i20686(x20686, x19380);
  not i20691(x20691, x19398);
  not i20692(x20692, x19389);
  not i20695(x20695, x20694);
  not i20697(x20697, x19407);
  not i20700(x20700, x20699);
  not i20705(x20705, x20704);
  not i20709(x20709, x20708);
  not i20714(x20714, x20713);
  not i20720(x20720, x19424);
  not i20721(x20721, x19415);
  not i20724(x20724, x20723);
  not i20726(x20726, x19433);
  not i20731(x20731, x19451);
  not i20732(x20732, x19442);
  not i20735(x20735, x20734);
  not i20737(x20737, x19460);
  not i20740(x20740, x20739);
  not i20745(x20745, x20744);
  not i20749(x20749, x20748);
  not i20754(x20754, x20753);
  not i20760(x20760, x19477);
  not i20761(x20761, x19468);
  not i20764(x20764, x20763);
  not i20766(x20766, x19486);
  not i20771(x20771, x19504);
  not i20772(x20772, x19495);
  not i20775(x20775, x20774);
  not i20777(x20777, x19513);
  not i20780(x20780, x20779);
  not i20785(x20785, x20784);
  not i20789(x20789, x20788);
  not i20794(x20794, x20793);
  not i20800(x20800, x19533);
  not i20801(x20801, x19524);
  not i20804(x20804, x20803);
  not i20806(x20806, x19542);
  not i20811(x20811, x19560);
  not i20812(x20812, x19551);
  not i20815(x20815, x20814);
  not i20817(x20817, x19569);
  not i20820(x20820, x20819);
  not i20822(x20822, x19578);
  not i20826(x20826, x20825);
  not i20830(x20830, x20829);
  not i20835(x20835, x20834);
  not i20839(x20839, x20838);
  not i20842(x20842, x19595);
  not i20843(x20843, x19586);
  not i20846(x20846, x20845);
  not i20848(x20848, x19604);
  not i20853(x20853, x19622);
  not i20854(x20854, x19613);
  not i20857(x20857, x20856);
  not i20859(x20859, x19631);
  not i20862(x20862, x20861);
  not i20864(x20864, x19640);
  not i20868(x20868, x20867);
  not i20872(x20872, x20871);
  not i20877(x20877, x20876);
  not i20881(x20881, x20880);
  not i20884(x20884, x19657);
  not i20885(x20885, x19648);
  not i20888(x20888, x20887);
  not i20890(x20890, x19666);
  not i20895(x20895, x19684);
  not i20896(x20896, x19675);
  not i20899(x20899, x20898);
  not i20901(x20901, x19693);
  not i20904(x20904, x20903);
  not i20907(x20907, x19702);
  not i20913(x20913, x20912);
  not i20917(x20917, x20916);
  not i20922(x20922, x20921);
  not i20926(x20926, x20925);
  not i20929(x20929, x19722);
  not i20930(x20930, x19713);
  not i20933(x20933, x20932);
  not i20935(x20935, x19731);
  not i20940(x20940, x19749);
  not i20941(x20941, x19740);
  not i20944(x20944, x20943);
  not i20946(x20946, x19758);
  not i20949(x20949, x20948);
  not i20952(x20952, x19775);
  not i20953(x20953, x19767);
  not i20959(x20959, x20958);
  not i20963(x20963, x20962);
  not i20968(x20968, x20967);
  not i20972(x20972, x20971);
  not i20978(x20978, x19792);
  not i20979(x20979, x19783);
  not i20982(x20982, x20981);
  not i20984(x20984, x19801);
  not i20987(x20987, x20986);
  not i20990(x20990, x19819);
  not i20991(x20991, x19810);
  not i20994(x20994, x20993);
  not i20996(x20996, x19828);
  not i20999(x20999, x20998);
  not i21002(x21002, x19846);
  not i21003(x21003, x19837);
  not i21009(x21009, x21008);
  not i21013(x21013, x21012);
  not i21018(x21018, x21017);
  not i21022(x21022, x21021);
  not i21028(x21028, x19863);
  not i21029(x21029, x19854);
  not i21032(x21032, x21031);
  not i21034(x21034, x19872);
  not i21037(x21037, x21036);
  not i21040(x21040, x19890);
  not i21041(x21041, x19881);
  not i21044(x21044, x21043);
  not i21046(x21046, x19899);
  not i21049(x21049, x21048);
  not i21052(x21052, x19917);
  not i21053(x21053, x19908);
  not i21056(x21056, x21055);
  not i21060(x21060, x21059);
  not i21065(x21065, x21064);
  not i21069(x21069, x21068);
  not i21074(x21074, x21073);
  not i21078(x21078, x21077);
  not i21084(x21084, x19937);
  not i21085(x21085, x19928);
  not i21088(x21088, x21087);
  not i21090(x21090, x19946);
  not i21093(x21093, x21092);
  not i21096(x21096, x19964);
  not i21097(x21097, x19955);
  not i21100(x21100, x21099);
  not i21102(x21102, x19973);
  not i21105(x21105, x21104);
  not i21108(x21108, x19991);
  not i21109(x21109, x19982);
  not i21112(x21112, x21111);
  not i21114(x21114, x20000);
  not i21117(x21117, x21116);
  not i21122(x21122, x21121);
  not i21126(x21126, x21125);
  not i21131(x21131, x21130);
  not i21135(x21135, x21134);
  not i21140(x21140, x21139);
  not i21144(x21144, x21143);
  not i21147(x21147, x20017);
  not i21148(x21148, x20008);
  not i21151(x21151, x21150);
  not i21153(x21153, x20026);
  not i21156(x21156, x21155);
  not i21159(x21159, x20044);
  not i21160(x21160, x20035);
  not i21163(x21163, x21162);
  not i21165(x21165, x20053);
  not i21168(x21168, x21167);
  not i21171(x21171, x20071);
  not i21172(x21172, x20062);
  not i21175(x21175, x21174);
  not i21177(x21177, x20080);
  not i21180(x21180, x21179);
  not i21185(x21185, x21184);
  not i21189(x21189, x21188);
  not i21194(x21194, x21193);
  not i21198(x21198, x21197);
  not i21203(x21203, x21202);
  not i21207(x21207, x21206);
  not i21210(x21210, x20097);
  not i21211(x21211, x20088);
  not i21214(x21214, x21213);
  not i21216(x21216, x20106);
  not i21219(x21219, x21218);
  not i21222(x21222, x20124);
  not i21223(x21223, x20115);
  not i21226(x21226, x21225);
  not i21228(x21228, x20133);
  not i21231(x21231, x21230);
  not i21234(x21234, x20151);
  not i21235(x21235, x20142);
  not i21238(x21238, x21237);
  not i21240(x21240, x20160);
  not i21243(x21243, x21242);
  not i21248(x21248, x21247);
  not i21252(x21252, x21251);
  not i21256(x21256, x21255);
  not i21261(x21261, x21260);
  not i21265(x21265, x21264);
  not i21270(x21270, x21269);
  not i21274(x21274, x21273);
  not i21277(x21277, x20181);
  not i21278(x21278, x20172);
  not i21281(x21281, x21280);
  not i21283(x21283, x20190);
  not i21286(x21286, x21285);
  not i21289(x21289, x20208);
  not i21290(x21290, x20199);
  not i21293(x21293, x21292);
  not i21295(x21295, x20217);
  not i21298(x21298, x21297);
  not i21301(x21301, x20235);
  not i21302(x21302, x20226);
  not i21305(x21305, x21304);
  not i21307(x21307, x20244);
  not i21310(x21310, x21309);
  not i21312(x21312, x20253);
  not i21316(x21316, x21315);
  not i21320(x21320, x21319);
  not i21324(x21324, x21323);
  not i21329(x21329, x21328);
  not i21333(x21333, x21332);
  not i21338(x21338, x21337);
  not i21342(x21342, x21341);
  not i21345(x21345, x20271);
  not i21346(x21346, x20262);
  not i21349(x21349, x21348);
  not i21351(x21351, x20280);
  not i21354(x21354, x21353);
  not i21356(x21356, x20298);
  not i21357(x21357, x20289);
  not i21360(x21360, x21359);
  not i21362(x21362, x20307);
  not i21365(x21365, x21364);
  not i21367(x21367, x20325);
  not i21368(x21368, x20316);
  not i21371(x21371, x21370);
  not i21373(x21373, x20334);
  not i21376(x21376, x21375);
  not i21377(x21377, x20343);
  not i21381(x21381, x21380);
  not i21385(x21385, x21384);
  not i21389(x21389, x21388);
  not i21393(x21393, x21392);
  not i21397(x21397, x21396);
  not i21401(x21401, x21400);
  not i21405(x21405, x21404);
  not i21409(x21409, x21408);
  not i21413(x21413, x21412);
  not i21417(x21417, x21416);
  not i21421(x21421, x21420);
  not i21425(x21425, x21424);
  not i21429(x21429, x21428);
  not i21430(x21430, x20459);
  not i21434(x21434, x21433);
  not i21435(x21435, x20473);
  not i21436(x21436, x20482);
  not i21440(x21440, x21439);
  not i21441(x21441, x20493);
  not i21442(x21442, x20502);
  not i21446(x21446, x21445);
  not i21450(x21450, x21449);
  not i21451(x21451, x20513);
  not i21452(x21452, x20522);
  not i21456(x21456, x21455);
  not i21460(x21460, x21459);
  not i21461(x21461, x20533);
  not i21462(x21462, x20543);
  not i21466(x21466, x21465);
  not i21470(x21470, x21469);
  not i21471(x21471, x20554);
  not i21472(x21472, x20564);
  not i21476(x21476, x21475);
  not i21480(x21480, x21479);
  not i21482(x21482, x20575);
  not i21485(x21485, x20588);
  not i21489(x21489, x21488);
  not i21493(x21493, x21492);
  not i21495(x21495, x20599);
  not i21498(x21498, x20613);
  not i21502(x21502, x21501);
  not i21506(x21506, x21505);
  not i21510(x21510, x21509);
  not i21512(x21512, x20627);
  not i21515(x21515, x20641);
  not i21519(x21519, x21518);
  not i21523(x21523, x21522);
  not i21527(x21527, x21526);
  not i21529(x21529, x20666);
  not i21530(x21530, x20655);
  not i21533(x21533, x20675);
  not i21537(x21537, x21536);
  not i21541(x21541, x21540);
  not i21545(x21545, x21544);
  not i21547(x21547, x20701);
  not i21548(x21548, x20689);
  not i21551(x21551, x20710);
  not i21553(x21553, x20718);
  not i21556(x21556, x21555);
  not i21560(x21560, x21559);
  not i21564(x21564, x21563);
  not i21566(x21566, x20741);
  not i21567(x21567, x20729);
  not i21570(x21570, x20750);
  not i21572(x21572, x20758);
  not i21575(x21575, x21574);
  not i21579(x21579, x21578);
  not i21583(x21583, x21582);
  not i21587(x21587, x21586);
  not i21590(x21590, x20781);
  not i21591(x21591, x20769);
  not i21594(x21594, x20790);
  not i21596(x21596, x20798);
  not i21599(x21599, x21598);
  not i21603(x21603, x21602);
  not i21607(x21607, x21606);
  not i21611(x21611, x21610);
  not i21617(x21617, x20821);
  not i21618(x21618, x20809);
  not i21621(x21621, x20831);
  not i21623(x21623, x20840);
  not i21626(x21626, x21625);
  not i21630(x21630, x21629);
  not i21634(x21634, x21633);
  not i21638(x21638, x21637);
  not i21644(x21644, x20863);
  not i21645(x21645, x20851);
  not i21648(x21648, x20873);
  not i21650(x21650, x20882);
  not i21653(x21653, x21652);
  not i21657(x21657, x21656);
  not i21661(x21661, x21660);
  not i21665(x21665, x21664);
  not i21671(x21671, x20905);
  not i21672(x21672, x20893);
  not i21675(x21675, x21674);
  not i21679(x21679, x21678);
  not i21681(x21681, x20918);
  not i21683(x21683, x20927);
  not i21686(x21686, x21685);
  not i21690(x21690, x21689);
  not i21694(x21694, x21693);
  not i21698(x21698, x21697);
  not i21704(x21704, x20950);
  not i21705(x21705, x20938);
  not i21708(x21708, x21707);
  not i21712(x21712, x21711);
  not i21714(x21714, x20964);
  not i21716(x21716, x20973);
  not i21719(x21719, x21718);
  not i21723(x21723, x21722);
  not i21727(x21727, x21726);
  not i21732(x21732, x21731);
  not i21736(x21736, x21735);
  not i21742(x21742, x21000);
  not i21743(x21743, x20988);
  not i21746(x21746, x21745);
  not i21750(x21750, x21749);
  not i21752(x21752, x21014);
  not i21754(x21754, x21023);
  not i21757(x21757, x21756);
  not i21761(x21761, x21760);
  not i21765(x21765, x21764);
  not i21770(x21770, x21769);
  not i21774(x21774, x21773);
  not i21780(x21780, x21050);
  not i21781(x21781, x21038);
  not i21784(x21784, x21783);
  not i21786(x21786, x21061);
  not i21789(x21789, x21788);
  not i21791(x21791, x21070);
  not i21793(x21793, x21079);
  not i21796(x21796, x21795);
  not i21800(x21800, x21799);
  not i21804(x21804, x21803);
  not i21809(x21809, x21808);
  not i21813(x21813, x21812);
  not i21819(x21819, x21106);
  not i21820(x21820, x21094);
  not i21823(x21823, x21822);
  not i21825(x21825, x21118);
  not i21828(x21828, x21827);
  not i21830(x21830, x21127);
  not i21832(x21832, x21136);
  not i21835(x21835, x21834);
  not i21837(x21837, x21145);
  not i21840(x21840, x21839);
  not i21844(x21844, x21843);
  not i21849(x21849, x21848);
  not i21853(x21853, x21852);
  not i21859(x21859, x21169);
  not i21860(x21860, x21157);
  not i21863(x21863, x21862);
  not i21865(x21865, x21181);
  not i21868(x21868, x21867);
  not i21870(x21870, x21190);
  not i21872(x21872, x21199);
  not i21875(x21875, x21874);
  not i21877(x21877, x21208);
  not i21880(x21880, x21879);
  not i21884(x21884, x21883);
  not i21889(x21889, x21888);
  not i21893(x21893, x21892);
  not i21899(x21899, x21232);
  not i21900(x21900, x21220);
  not i21903(x21903, x21902);
  not i21905(x21905, x21244);
  not i21908(x21908, x21907);
  not i21911(x21911, x21257);
  not i21914(x21914, x21913);
  not i21916(x21916, x21266);
  not i21919(x21919, x21918);
  not i21922(x21922, x21275);
  not i21925(x21925, x21924);
  not i21929(x21929, x21928);
  not i21934(x21934, x21933);
  not i21938(x21938, x21937);
  not i21943(x21943, x21942);
  not i21947(x21947, x21946);
  not i21950(x21950, x21299);
  not i21951(x21951, x21287);
  not i21954(x21954, x21953);
  not i21956(x21956, x21311);
  not i21959(x21959, x21958);
  not i21961(x21961, x21325);
  not i21964(x21964, x21963);
  not i21966(x21966, x21334);
  not i21969(x21969, x21968);
  not i21971(x21971, x21343);
  not i21974(x21974, x21973);
  not i21978(x21978, x21977);
  not i21982(x21982, x21981);
  not i21986(x21986, x21985);
  not i21990(x21990, x21989);
  not i21994(x21994, x21993);
  not i22004(x22004, x22003);
  not i22008(x22008, x22007);
  not i22015(x22015, x22014);
  not i22022(x22022, x22021);
  not i22026(x22026, x22025);
  not i22034(x22034, x22033);
  not i22038(x22038, x22037);
  not i22046(x22046, x22045);
  not i22050(x22050, x22049);
  not i22058(x22058, x22057);
  not i22062(x22062, x22061);
  not i22070(x22070, x22069);
  not i22074(x22074, x22073);
  not i22079(x22079, x22078);
  not i22083(x22083, x22082);
  not i22087(x22087, x22086);
  not i22092(x22092, x22091);
  not i22096(x22096, x22095);
  not i22100(x22100, x22099);
  not i22105(x22105, x22104);
  not i22109(x22109, x22108);
  not i22113(x22113, x22112);
  not i22118(x22118, x22117);
  not i22122(x22122, x22121);
  not i22126(x22126, x22125);
  not i22131(x22131, x22130);
  not i22135(x22135, x22134);
  not i22139(x22139, x22138);
  not i22143(x22143, x22142);
  not i22148(x22148, x22147);
  not i22152(x22152, x22151);
  not i22157(x22157, x22156);
  not i22161(x22161, x22160);
  not i22165(x22165, x22164);
  not i22170(x22170, x22169);
  not i22174(x22174, x22173);
  not i22179(x22179, x22178);
  not i22183(x22183, x22182);
  not i22187(x22187, x22186);
  not i22192(x22192, x22191);
  not i22196(x22196, x22195);
  not i22201(x22201, x22200);
  not i22205(x22205, x22204);
  not i22209(x22209, x22208);
  not i22214(x22214, x22213);
  not i22218(x22218, x22217);
  not i22223(x22223, x22222);
  not i22227(x22227, x22226);
  not i22231(x22231, x22230);
  not i22236(x22236, x22235);
  not i22240(x22240, x22239);
  not i22242(x22242, x21588);
  not i22246(x22246, x22245);
  not i22250(x22250, x22249);
  not i22254(x22254, x22253);
  not i22259(x22259, x22258);
  not i22263(x22263, x22262);
  not i22266(x22266, x21612);
  not i22269(x22269, x22268);
  not i22273(x22273, x22272);
  not i22278(x22278, x22277);
  not i22282(x22282, x22281);
  not i22287(x22287, x22286);
  not i22291(x22291, x22290);
  not i22294(x22294, x21639);
  not i22297(x22297, x22296);
  not i22301(x22301, x22300);
  not i22306(x22306, x22305);
  not i22310(x22310, x22309);
  not i22315(x22315, x22314);
  not i22319(x22319, x22318);
  not i22322(x22322, x21666);
  not i22325(x22325, x22324);
  not i22329(x22329, x22328);
  not i22334(x22334, x22333);
  not i22338(x22338, x22337);
  not i22341(x22341, x21680);
  not i22344(x22344, x22343);
  not i22348(x22348, x22347);
  not i22351(x22351, x21699);
  not i22354(x22354, x22353);
  not i22358(x22358, x22357);
  not i22363(x22363, x22362);
  not i22367(x22367, x22366);
  not i22370(x22370, x21713);
  not i22373(x22373, x22372);
  not i22375(x22375, x21728);
  not i22378(x22378, x22377);
  not i22381(x22381, x21737);
  not i22384(x22384, x22383);
  not i22388(x22388, x22387);
  not i22393(x22393, x22392);
  not i22397(x22397, x22396);
  not i22400(x22400, x21751);
  not i22403(x22403, x22402);
  not i22405(x22405, x21766);
  not i22408(x22408, x22407);
  not i22411(x22411, x21775);
  not i22414(x22414, x22413);
  not i22418(x22418, x22417);
  not i22423(x22423, x22422);
  not i22427(x22427, x22426);
  not i22430(x22430, x21790);
  not i22433(x22433, x22432);
  not i22435(x22435, x21805);
  not i22438(x22438, x22437);
  not i22441(x22441, x21814);
  not i22444(x22444, x22443);
  not i22448(x22448, x22447);
  not i22453(x22453, x22452);
  not i22457(x22457, x22456);
  not i22460(x22460, x21829);
  not i22463(x22463, x22462);
  not i22465(x22465, x21845);
  not i22468(x22468, x22467);
  not i22471(x22471, x21854);
  not i22474(x22474, x22473);
  not i22478(x22478, x22477);
  not i22483(x22483, x22482);
  not i22487(x22487, x22486);
  not i22490(x22490, x21869);
  not i22493(x22493, x22492);
  not i22495(x22495, x21885);
  not i22498(x22498, x22497);
  not i22501(x22501, x21894);
  not i22504(x22504, x22503);
  not i22508(x22508, x22507);
  not i22513(x22513, x22512);
  not i22517(x22517, x22516);
  not i22520(x22520, x21920);
  not i22521(x22521, x21909);
  not i22524(x22524, x22523);
  not i22526(x22526, x21930);
  not i22529(x22529, x22528);
  not i22531(x22531, x21948);
  not i22532(x22532, x21939);
  not i22535(x22535, x22534);
  not i22539(x22539, x22538);
  not i22543(x22543, x22542);
  not i22547(x22547, x22546);
  not i22560(x22560, x22559);
  not i22565(x22565, x22027);
  not i22568(x22568, x22567);
  not i22573(x22573, x22039);
  not i22576(x22576, x22575);
  not i22581(x22581, x22051);
  not i22584(x22584, x22583);
  not i22589(x22589, x22063);
  not i22592(x22592, x22591);
  not i22597(x22597, x22075);
  not i22600(x22600, x22599);
  not i22604(x22604, x22603);
  not i22608(x22608, x22607);
  not i22611(x22611, x22088);
  not i22614(x22614, x22613);
  not i22618(x22618, x22617);
  not i22622(x22622, x22621);
  not i22625(x22625, x22101);
  not i22628(x22628, x22627);
  not i22632(x22632, x22631);
  not i22636(x22636, x22635);
  not i22639(x22639, x22114);
  not i22642(x22642, x22641);
  not i22646(x22646, x22645);
  not i22650(x22650, x22649);
  not i22653(x22653, x22127);
  not i22656(x22656, x22655);
  not i22660(x22660, x22659);
  not i22664(x22664, x22663);
  not i22669(x22669, x22668);
  not i22671(x22671, x22144);
  not i22674(x22674, x22673);
  not i22679(x22679, x22678);
  not i22683(x22683, x22682);
  not i22686(x22686, x22153);
  not i22689(x22689, x22688);
  not i22691(x22691, x22166);
  not i22694(x22694, x22693);
  not i22699(x22699, x22698);
  not i22703(x22703, x22702);
  not i22706(x22706, x22175);
  not i22709(x22709, x22708);
  not i22711(x22711, x22188);
  not i22714(x22714, x22713);
  not i22719(x22719, x22718);
  not i22723(x22723, x22722);
  not i22726(x22726, x22197);
  not i22729(x22729, x22728);
  not i22731(x22731, x22210);
  not i22734(x22734, x22733);
  not i22739(x22739, x22738);
  not i22743(x22743, x22742);
  not i22746(x22746, x22219);
  not i22749(x22749, x22748);
  not i22751(x22751, x22232);
  not i22754(x22754, x22753);
  not i22759(x22759, x22758);
  not i22763(x22763, x22762);
  not i22766(x22766, x22241);
  not i22769(x22769, x22768);
  not i22771(x22771, x22255);
  not i22774(x22774, x22773);
  not i22779(x22779, x22778);
  not i22783(x22783, x22782);
  not i22786(x22786, x22274);
  not i22787(x22787, x22264);
  not i22790(x22790, x22789);
  not i22792(x22792, x22283);
  not i22795(x22795, x22794);
  not i22800(x22800, x22799);
  not i22804(x22804, x22803);
  not i22807(x22807, x22302);
  not i22808(x22808, x22292);
  not i22811(x22811, x22810);
  not i22813(x22813, x22311);
  not i22816(x22816, x22815);
  not i22821(x22821, x22820);
  not i22825(x22825, x22824);
  not i22828(x22828, x22330);
  not i22829(x22829, x22320);
  not i22832(x22832, x22831);
  not i22834(x22834, x22339);
  not i22837(x22837, x22836);
  not i22842(x22842, x22841);
  not i22846(x22846, x22845);
  not i22849(x22849, x22359);
  not i22850(x22850, x22349);
  not i22853(x22853, x22852);
  not i22855(x22855, x22368);
  not i22858(x22858, x22857);
  not i22863(x22863, x22862);
  not i22867(x22867, x22866);
  not i22870(x22870, x22389);
  not i22871(x22871, x22379);
  not i22874(x22874, x22873);
  not i22876(x22876, x22398);
  not i22879(x22879, x22878);
  not i22884(x22884, x22883);
  not i22888(x22888, x22887);
  not i22891(x22891, x22419);
  not i22892(x22892, x22409);
  not i22895(x22895, x22894);
  not i22897(x22897, x22428);
  not i22900(x22900, x22899);
  not i22905(x22905, x22904);
  not i22909(x22909, x22908);
  not i22912(x22912, x22449);
  not i22913(x22913, x22439);
  not i22916(x22916, x22915);
  not i22918(x22918, x22458);
  not i22921(x22921, x22920);
  not i22926(x22926, x22925);
  not i22930(x22930, x22929);
  not i22933(x22933, x22479);
  not i22934(x22934, x22469);
  not i22937(x22937, x22936);
  not i22939(x22939, x22488);
  not i22942(x22942, x22941);
  not i22947(x22947, x22946);
  not i22951(x22951, x22950);
  not i22954(x22954, x22509);
  not i22955(x22955, x22499);
  not i22958(x22958, x22957);
  not i22960(x22960, x22518);
  not i22963(x22963, x22962);
  not i22967(x22967, x22966);
  not i22971(x22971, x22970);
  not i22978(x22978, x22977);
  not i22982(x22982, x22981);
  not i22986(x22986, x22985);
  not i22990(x22990, x22989);
  not i22995(x22995, x22994);
  not i22999(x22999, x22998);
  not i23004(x23004, x23003);
  not i23008(x23008, x23007);
  not i23013(x23013, x23012);
  not i23017(x23017, x23016);
  not i23022(x23022, x23021);
  not i23026(x23026, x23025);
  not i23031(x23031, x23030);
  not i23032(x23032, x23028);
  not i23034(x23034, x22609);
  not i23037(x23037, x23036);
  not i23041(x23041, x23040);
  not i23046(x23046, x23045);
  not i23047(x23047, x23043);
  not i23049(x23049, x22623);
  not i23052(x23052, x23051);
  not i23056(x23056, x23055);
  not i23061(x23061, x23060);
  not i23062(x23062, x23058);
  not i23064(x23064, x22637);
  not i23067(x23067, x23066);
  not i23071(x23071, x23070);
  not i23076(x23076, x23075);
  not i23077(x23077, x23073);
  not i23079(x23079, x22651);
  not i23082(x23082, x23081);
  not i23086(x23086, x23085);
  not i23091(x23091, x23090);
  not i23092(x23092, x23088);
  not i23094(x23094, x22665);
  not i23097(x23097, x23096);
  not i23101(x23101, x23100);
  not i23106(x23106, x23105);
  not i23107(x23107, x23103);
  not i23109(x23109, x22684);
  not i23110(x23110, x22675);
  not i23113(x23113, x23112);
  not i23117(x23117, x23116);
  not i23122(x23122, x23121);
  not i23123(x23123, x23119);
  not i23125(x23125, x22704);
  not i23126(x23126, x22695);
  not i23129(x23129, x23128);
  not i23133(x23133, x23132);
  not i23138(x23138, x23137);
  not i23139(x23139, x23135);
  not i23141(x23141, x22724);
  not i23142(x23142, x22715);
  not i23145(x23145, x23144);
  not i23149(x23149, x23148);
  not i23154(x23154, x23153);
  not i23155(x23155, x23151);
  not i23157(x23157, x22744);
  not i23158(x23158, x22735);
  not i23161(x23161, x23160);
  not i23165(x23165, x23164);
  not i23170(x23170, x23169);
  not i23171(x23171, x23167);
  not i23173(x23173, x22764);
  not i23174(x23174, x22755);
  not i23177(x23177, x23176);
  not i23181(x23181, x23180);
  not i23186(x23186, x23185);
  not i23187(x23187, x23183);
  not i23189(x23189, x22784);
  not i23190(x23190, x22775);
  not i23193(x23193, x23192);
  not i23197(x23197, x23196);
  not i23202(x23202, x23201);
  not i23203(x23203, x23199);
  not i23205(x23205, x22805);
  not i23206(x23206, x22796);
  not i23209(x23209, x23208);
  not i23213(x23213, x23212);
  not i23218(x23218, x23217);
  not i23219(x23219, x23215);
  not i23221(x23221, x22826);
  not i23222(x23222, x22817);
  not i23225(x23225, x23224);
  not i23229(x23229, x23228);
  not i23234(x23234, x23233);
  not i23235(x23235, x23231);
  not i23237(x23237, x22847);
  not i23238(x23238, x22838);
  not i23241(x23241, x23240);
  not i23245(x23245, x23244);
  not i23250(x23250, x23249);
  not i23251(x23251, x23247);
  not i23253(x23253, x22868);
  not i23254(x23254, x22859);
  not i23257(x23257, x23256);
  not i23261(x23261, x23260);
  not i23266(x23266, x23265);
  not i23267(x23267, x23263);
  not i23269(x23269, x22889);
  not i23270(x23270, x22880);
  not i23273(x23273, x23272);
  not i23277(x23277, x23276);
  not i23282(x23282, x23281);
  not i23283(x23283, x23279);
  not i23285(x23285, x22910);
  not i23286(x23286, x22901);
  not i23289(x23289, x23288);
  not i23293(x23293, x23292);
  not i23298(x23298, x23297);
  not i23299(x23299, x23295);
  not i23301(x23301, x22931);
  not i23302(x23302, x22922);
  not i23305(x23305, x23304);
  not i23309(x23309, x23308);
  not i23314(x23314, x23313);
  not i23315(x23315, x23311);
  not i23317(x23317, x22952);
  not i23318(x23318, x22943);
  not i23321(x23321, x23320);
  not i23325(x23325, x23324);
  not i23329(x23329, x23328);
  not i23339(x23339, x23338);
  not i23343(x23343, x23342);
  not i23344(x23344, x22991);
  not i23348(x23348, x23347);
  not i23349(x23349, x23000);
  not i23353(x23353, x23352);
  not i23354(x23354, x23009);
  not i23358(x23358, x23357);
  not i23359(x23359, x23018);
  not i23363(x23363, x23362);
  not i23365(x23365, x23027);
  not i23368(x23368, x23367);
  not i23372(x23372, x23371);
  not i23375(x23375, x23042);
  not i23378(x23378, x23377);
  not i23382(x23382, x23381);
  not i23385(x23385, x23057);
  not i23388(x23388, x23387);
  not i23392(x23392, x23391);
  not i23395(x23395, x23072);
  not i23398(x23398, x23397);
  not i23402(x23402, x23401);
  not i23405(x23405, x23087);
  not i23408(x23408, x23407);
  not i23412(x23412, x23411);
  not i23415(x23415, x23102);
  not i23418(x23418, x23417);
  not i23422(x23422, x23421);
  not i23425(x23425, x23118);
  not i23428(x23428, x23427);
  not i23432(x23432, x23431);
  not i23435(x23435, x23134);
  not i23438(x23438, x23437);
  not i23442(x23442, x23441);
  not i23445(x23445, x23150);
  not i23448(x23448, x23447);
  not i23452(x23452, x23451);
  not i23455(x23455, x23166);
  not i23458(x23458, x23457);
  not i23462(x23462, x23461);
  not i23465(x23465, x23182);
  not i23468(x23468, x23467);
  not i23472(x23472, x23471);
  not i23475(x23475, x23198);
  not i23478(x23478, x23477);
  not i23482(x23482, x23481);
  not i23485(x23485, x23214);
  not i23488(x23488, x23487);
  not i23492(x23492, x23491);
  not i23495(x23495, x23230);
  not i23498(x23498, x23497);
  not i23502(x23502, x23501);
  not i23505(x23505, x23246);
  not i23508(x23508, x23507);
  not i23512(x23512, x23511);
  not i23515(x23515, x23262);
  not i23518(x23518, x23517);
  not i23522(x23522, x23521);
  not i23525(x23525, x23278);
  not i23528(x23528, x23527);
  not i23532(x23532, x23531);
  not i23535(x23535, x23294);
  not i23538(x23538, x23537);
  not i23542(x23542, x23541);
  not i23545(x23545, x23310);
  not i23548(x23548, x23547);
  not i23552(x23552, x23551);
  not i23556(x23556, x23555);
  not i23564(x23564, x23563);
  not i23568(x23568, x23567);
  not i23572(x23572, x23571);
  not i23576(x23576, x23575);
  not i23581(x23581, x23580);
  not i23585(x23585, x23584);
  not i23590(x23590, x23589);
  not i23594(x23594, x23593);
  not i23599(x23599, x23598);
  not i23603(x23603, x23602);
  not i23608(x23608, x23607);
  not i23612(x23612, x23611);
  not i23617(x23617, x23616);
  not i23621(x23621, x23620);
  not i23626(x23626, x23625);
  not i23630(x23630, x23629);
  not i23633(x23633, x23373);
  not i23636(x23636, x23635);
  not i23640(x23640, x23639);
  not i23643(x23643, x23383);
  not i23646(x23646, x23645);
  not i23650(x23650, x23649);
  not i23653(x23653, x23393);
  not i23656(x23656, x23655);
  not i23660(x23660, x23659);
  not i23663(x23663, x23403);
  not i23666(x23666, x23665);
  not i23670(x23670, x23669);
  not i23673(x23673, x23413);
  not i23676(x23676, x23675);
  not i23680(x23680, x23679);
  not i23683(x23683, x23423);
  not i23686(x23686, x23685);
  not i23690(x23690, x23689);
  not i23693(x23693, x23433);
  not i23696(x23696, x23695);
  not i23700(x23700, x23699);
  not i23703(x23703, x23443);
  not i23706(x23706, x23705);
  not i23710(x23710, x23709);
  not i23713(x23713, x23453);
  not i23716(x23716, x23715);
  not i23720(x23720, x23719);
  not i23723(x23723, x23463);
  not i23726(x23726, x23725);
  not i23730(x23730, x23729);
  not i23733(x23733, x23473);
  not i23736(x23736, x23735);
  not i23740(x23740, x23739);
  not i23743(x23743, x23483);
  not i23746(x23746, x23745);
  not i23750(x23750, x23749);
  not i23753(x23753, x23493);
  not i23756(x23756, x23755);
  not i23760(x23760, x23759);
  not i23763(x23763, x23503);
  not i23766(x23766, x23765);
  not i23770(x23770, x23769);
  not i23773(x23773, x23513);
  not i23776(x23776, x23775);
  not i23780(x23780, x23779);
  not i23783(x23783, x23523);
  not i23786(x23786, x23785);
  not i23790(x23790, x23789);
  not i23793(x23793, x23533);
  not i23796(x23796, x23795);
  not i23800(x23800, x23799);
  not i23803(x23803, x23543);
  not i23806(x23806, x23805);
  not i23810(x23810, x23809);
  not i23812(x23812, x23560);
  not i23818(x23818, x23817);
  not i23822(x23822, x23821);
  not i23824(x23824, x23577);
  not i23827(x23827, x23826);
  not i23829(x23829, x23586);
  not i23832(x23832, x23831);
  not i23834(x23834, x23595);
  not i23837(x23837, x23836);
  not i23839(x23839, x23604);
  not i23842(x23842, x23841);
  not i23844(x23844, x23613);
  not i23847(x23847, x23846);
  not i23849(x23849, x23622);
  not i23852(x23852, x23851);
  not i23854(x23854, x23631);
  not i23857(x23857, x23856);
  not i23859(x23859, x23641);
  not i23862(x23862, x23861);
  not i23864(x23864, x23651);
  not i23867(x23867, x23866);
  not i23869(x23869, x23661);
  not i23872(x23872, x23871);
  not i23874(x23874, x23671);
  not i23877(x23877, x23876);
  not i23879(x23879, x23681);
  not i23882(x23882, x23881);
  not i23884(x23884, x23691);
  not i23887(x23887, x23886);
  not i23889(x23889, x23701);
  not i23892(x23892, x23891);
  not i23894(x23894, x23711);
  not i23897(x23897, x23896);
  not i23899(x23899, x23721);
  not i23902(x23902, x23901);
  not i23904(x23904, x23731);
  not i23907(x23907, x23906);
  not i23909(x23909, x23741);
  not i23912(x23912, x23911);
  not i23914(x23914, x23751);
  not i23917(x23917, x23916);
  not i23919(x23919, x23761);
  not i23922(x23922, x23921);
  not i23924(x23924, x23771);
  not i23927(x23927, x23926);
  not i23929(x23929, x23781);
  not i23932(x23932, x23931);
  not i23934(x23934, x23791);
  not i23937(x23937, x23936);
  not i23939(x23939, x23801);
  not i23942(x23942, x23941);
  not i23943(x23943, x23811);
  not i23944(x23944, x23815);
  not i23945(x23945, x23819);
  not i23946(x23946, x23823);
  not i23947(x23947, x23828);
  not i23948(x23948, x23833);
  not i23949(x23949, x23838);
  not i23950(x23950, x23843);
  not i23951(x23951, x23848);
  not i23952(x23952, x23853);
  not i23953(x23953, x23858);
  not i23954(x23954, x23863);
  not i23955(x23955, x23868);
  not i23956(x23956, x23873);
  not i23957(x23957, x23878);
  not i23958(x23958, x23883);
  not i23959(x23959, x23888);
  not i23960(x23960, x23893);
  not i23961(x23961, x23898);
  not i23962(x23962, x23903);
  not i23963(x23963, x23908);
  not i23964(x23964, x23913);
  not i23965(x23965, x23918);
  not i23966(x23966, x23923);
  not i23967(x23967, x23928);
  not i23973(x23973, x23972);
  not i23977(x23977, x23976);
  not i23981(x23981, x23980);
  not i23985(x23985, x23984);
  not i23989(x23989, x23988);
  not i23993(x23993, x23992);
  not i23997(x23997, x23996);
  not i24001(x24001, x24000);
  not i24005(x24005, x24004);
  not i24009(x24009, x24008);
  not i24013(x24013, x24012);
  not i24017(x24017, x24016);
  not i24021(x24021, x24020);
  not i24025(x24025, x24024);
  not i24029(x24029, x24028);
  not i24033(x24033, x24032);
  not i24037(x24037, x24036);
  not i24041(x24041, x24040);
  not i24045(x24045, x24044);
  not i24049(x24049, x24048);
  not i24053(x24053, x24052);
  not i24057(x24057, x24056);
  not i24061(x24061, x24060);
  not i24065(x24065, x24064);
  not i24066(x24066, x23969);
  not i24068(x24068, x23971);
  not i24071(x24071, x23975);
  not i24074(x24074, x23979);
  not i24077(x24077, x24076);
  not i24079(x24079, x23983);
  not i24082(x24082, x24081);
  not i24084(x24084, x23987);
  not i24087(x24087, x24086);
  not i24089(x24089, x23991);
  not i24092(x24092, x24091);
  not i24094(x24094, x23995);
  not i24097(x24097, x24096);
  not i24099(x24099, x23999);
  not i24102(x24102, x24101);
  not i24104(x24104, x24003);
  not i24107(x24107, x24106);
  not i24109(x24109, x24007);
  not i24112(x24112, x24111);
  not i24114(x24114, x24011);
  not i24117(x24117, x24116);
  not i24119(x24119, x24015);
  not i24122(x24122, x24121);
  not i24124(x24124, x24019);
  not i24127(x24127, x24126);
  not i24129(x24129, x24023);
  not i24132(x24132, x24131);
  not i24134(x24134, x24027);
  not i24137(x24137, x24136);
  not i24139(x24139, x24031);
  not i24142(x24142, x24141);
  not i24144(x24144, x24035);
  not i24147(x24147, x24146);
  not i24149(x24149, x24039);
  not i24152(x24152, x24151);
  not i24154(x24154, x24043);
  not i24157(x24157, x24156);
  not i24159(x24159, x24047);
  not i24162(x24162, x24161);
  not i24164(x24164, x24051);
  not i24167(x24167, x24166);
  not i24169(x24169, x24055);
  not i24172(x24172, x24171);
  not i24174(x24174, x24059);
  not i24177(x24177, x24176);
  not i24179(x24179, x24063);
  not i24182(x24182, x24181);
  not i24183(x24183, x24069);
  not i24184(x24184, x24072);
  not i24186(x24186, x24075);
  not i24189(x24189, x24080);
  not i24192(x24192, x24085);
  not i24195(x24195, x24090);
  not i24198(x24198, x24095);
  not i24201(x24201, x24200);
  not i24203(x24203, x24100);
  not i24206(x24206, x24205);
  not i24208(x24208, x24105);
  not i24211(x24211, x24210);
  not i24213(x24213, x24110);
  not i24216(x24216, x24215);
  not i24218(x24218, x24115);
  not i24221(x24221, x24220);
  not i24223(x24223, x24120);
  not i24226(x24226, x24225);
  not i24228(x24228, x24125);
  not i24231(x24231, x24230);
  not i24233(x24233, x24130);
  not i24236(x24236, x24235);
  not i24238(x24238, x24135);
  not i24241(x24241, x24240);
  not i24243(x24243, x24140);
  not i24246(x24246, x24245);
  not i24248(x24248, x24145);
  not i24251(x24251, x24250);
  not i24253(x24253, x24150);
  not i24256(x24256, x24255);
  not i24258(x24258, x24155);
  not i24261(x24261, x24260);
  not i24263(x24263, x24160);
  not i24266(x24266, x24265);
  not i24268(x24268, x24165);
  not i24271(x24271, x24270);
  not i24273(x24273, x24170);
  not i24276(x24276, x24275);
  not i24278(x24278, x24175);
  not i24281(x24281, x24280);
  not i24283(x24283, x24180);
  not i24286(x24286, x24285);
  not i24287(x24287, x24187);
  not i24288(x24288, x24190);
  not i24289(x24289, x24193);
  not i24290(x24290, x24196);
  not i24292(x24292, x24199);
  not i24295(x24295, x24204);
  not i24298(x24298, x24209);
  not i24301(x24301, x24214);
  not i24304(x24304, x24219);
  not i24307(x24307, x24224);
  not i24310(x24310, x24229);
  not i24313(x24313, x24234);
  not i24316(x24316, x24239);
  not i24319(x24319, x24318);
  not i24321(x24321, x24244);
  not i24324(x24324, x24323);
  not i24326(x24326, x24249);
  not i24329(x24329, x24328);
  not i24331(x24331, x24254);
  not i24334(x24334, x24333);
  not i24336(x24336, x24259);
  not i24339(x24339, x24338);
  not i24341(x24341, x24264);
  not i24344(x24344, x24343);
  not i24346(x24346, x24269);
  not i24349(x24349, x24348);
  not i24351(x24351, x24274);
  not i24354(x24354, x24353);
  not i24356(x24356, x24279);
  not i24359(x24359, x24358);
  not i24361(x24361, x24284);
  not i24364(x24364, x24363);
  not i24365(x24365, x24299);
  not i24366(x24366, x24302);
  not i24367(x24367, x24305);
  not i24368(x24368, x24308);
  not i24369(x24369, x24311);
  not i24370(x24370, x24314);
  not i24372(x24372, x24317);
  not i24375(x24375, x24322);
  not i24378(x24378, x24327);
  not i24381(x24381, x24332);
  not i24384(x24384, x24337);
  not i24387(x24387, x24342);
  not i24390(x24390, x24347);
  not i24393(x24393, x24352);
  not i24396(x24396, x24357);
  not i24399(x24399, x24362);
  not i24403(x24403, x24402);
  not i24407(x24407, x24406);
  not i24411(x24411, x24410);
  not i24415(x24415, x24414);
  not i24419(x24419, x24418);
  not i24423(x24423, x24422);
  not i24427(x24427, x24426);
  not i24431(x24431, x24430);
  not i24433(x24433, x24293);
  not i24436(x24436, x24435);
  not i24438(x24438, x24296);
  not i24441(x24441, x24440);
  not i24445(x24445, x24444);
  not i24449(x24449, x24448);
  not i24453(x24453, x24452);
  not i24457(x24457, x24456);
  not i24461(x24461, x24460);
  not i24465(x24465, x24464);
  not i24467(x24467, x24373);
  not i24470(x24470, x24469);
  not i24472(x24472, x24376);
  not i24475(x24475, x24474);
  not i24477(x24477, x24379);
  not i24480(x24480, x24479);
  not i24482(x24482, x24382);
  not i24485(x24485, x24484);
  not i24487(x24487, x24385);
  not i24490(x24490, x24489);
  not i24492(x24492, x24388);
  not i24495(x24495, x24494);
  not i24497(x24497, x24391);
  not i24500(x24500, x24499);
  not i24502(x24502, x24394);
  not i24505(x24505, x24504);
  not i24507(x24507, x24397);
  not i24510(x24510, x24509);
  not i24512(x24512, x24400);
  not i24515(x24515, x24514);
  not i24517(x24517, x24516);
  not i24519(x24519, x24518);
  not i24521(x24521, x24520);
  not i24523(x24523, x24522);
  not i24525(x24525, x24524);
  not i24527(x24527, x24526);
  not i24529(x24529, x24528);
  not i24531(x24531, x24530);
  not i24533(x24533, x24532);
  not i24535(x24535, x24534);
  not i24537(x24537, x24536);
  not i24539(x24539, x24538);
  not i24541(x24541, x24540);
  not i24543(x24543, x24542);
  not i24545(x24545, x24544);
  not i24547(x24547, x24546);
  not i24549(x24549, x24548);
  not i24551(x24551, x24550);
  not i24553(x24553, x24552);
  not i24555(x24555, x24554);
  not i24557(x24557, x24556);
  not i24559(x24559, x24558);
  not i24561(x24561, x24560);
  not i24563(x24563, x24562);
  not i24565(x24565, x24564);
  not i24567(x24567, x24566);
  not i24569(x24569, x24568);
  not i24571(x24571, x24570);
  not i24573(x24573, x24572);
  not i24575(x24575, x24574);
  not i24578(x24578, x24577);
  not i24580(x24580, x24579);
  not i24582(x24582, x24581);
  not i24584(x24584, x24583);
  not i24586(x24586, x24585);
  not i24588(x24588, x24587);
  not i24590(x24590, x24589);
  not i24592(x24592, x24591);
  not i24594(x24594, x24593);
  not i24596(x24596, x24595);
  not i24598(x24598, x24597);
  not i24600(x24600, x24599);
  not i24602(x24602, x24601);
  not i24604(x24604, x24603);
  not i24606(x24606, x24605);
  not i24608(x24608, x24607);
  not i24610(x24610, x24609);
  not i24612(x24612, x24611);
  not i24614(x24614, x24613);
  not i24616(x24616, x24615);
  not i24618(x24618, x24617);
  not i24620(x24620, x24619);
  not i24622(x24622, x24621);
  not i24624(x24624, x24623);
  not i24626(x24626, x24625);
  not i24628(x24628, x24627);
  not i24630(x24630, x24629);
  not i24632(x24632, x24631);
  not i24637(x24637, x24636);
  not i24639(x24639, x24638);
  not i24641(x24641, x24640);
  not i24643(x24643, x24642);
  not i24645(x24645, x24644);
  not i24647(x24647, x24646);
  not i24649(x24649, x24648);
  not i24651(x24651, x24650);
  not i24653(x24653, x24652);
  not i24655(x24655, x24654);
  not i24657(x24657, x24656);
  not i24659(x24659, x24658);
  not i24661(x24661, x24660);
  not i24663(x24663, x24662);
  not i24665(x24665, x24664);
  not i24667(x24667, x24666);
  not i24669(x24669, x24668);
  not i24671(x24671, x24670);
  not i24673(x24673, x24672);
  not i24675(x24675, x24674);
  not i24677(x24677, x24676);
  not i24679(x24679, x24678);
  not i24681(x24681, x24680);
  not i24683(x24683, x24682);
  not i24693(x24693, x24692);
  not i24695(x24695, x24694);
  not i24697(x24697, x24696);
  not i24699(x24699, x24698);
  not i24701(x24701, x24700);
  not i24703(x24703, x24702);
  not i24705(x24705, x24704);
  not i24707(x24707, x24706);
  not i24709(x24709, x24708);
  not i24711(x24711, x24710);
  not i24713(x24713, x24712);
  not i24715(x24715, x24714);
  not i24717(x24717, x24716);
  not i24719(x24719, x24718);
  not i24721(x24721, x24720);
  not i24739(x24739, x24738);
  not i24743(x24743, x24742);
  not i24747(x24747, x24746);
  not i24751(x24751, x24750);
  not i24755(x24755, x24754);
  not i24759(x24759, x24758);
  not i24763(x24763, x24762);
  not i24767(x24767, x24766);
  not i24771(x24771, x24770);
  not i24775(x24775, x24774);
  not i24779(x24779, x24778);
  not i24783(x24783, x24782);
  not i24787(x24787, x24786);
  not i24791(x24791, x24790);
  not i24795(x24795, x24794);
  not i24799(x24799, x24798);
  not i24803(x24803, x24802);
  not i24807(x24807, x24806);
  not i24811(x24811, x24810);
  not i24815(x24815, x24814);
  not i24819(x24819, x24818);
  not i24823(x24823, x24822);
  not i24827(x24827, x24826);
  not i24831(x24831, x24830);
  not i24835(x24835, x24834);
  not i24839(x24839, x24838);
  not i24843(x24843, x24842);
  not i24847(x24847, x24846);
  not i24851(x24851, x24850);
  not i24855(x24855, x24854);
  not i24859(x24859, x24858);
  not i24860(x24860, x17904);
  not i24862(x24862, x24861);
  not i24864(x24864, x24863);
  not i24866(x24866, x24865);
  not i24868(x24868, x24867);
  not i24870(x24870, x24869);
  not i24872(x24872, x24871);
  not i24874(x24874, x24873);
  not i24876(x24876, x24875);
  not i24878(x24878, x24877);
  not i24880(x24880, x24879);
  not i24882(x24882, x24881);
  not i24884(x24884, x24883);
  not i24886(x24886, x24885);
  not i24888(x24888, x24887);
  not i24890(x24890, x24889);
  not i24892(x24892, x24891);
  not i24926(x24926, x24925);
  not i24928(x24928, x24927);
  not i24930(x24930, x24929);
  not i24932(x24932, x24931);
  not i24934(x24934, x24933);
  not i24936(x24936, x24935);
  not i24938(x24938, x24937);
  not i24940(x24940, x24939);
  not i24942(x24942, x24941);
  not i24944(x24944, x24943);
  not i24946(x24946, x24945);
  not i24948(x24948, x24947);
  not i24950(x24950, x24949);
  not i24952(x24952, x24951);
  not i24954(x24954, x24953);
  not i24956(x24956, x24955);
  not i24958(x24958, x24957);
  not i24960(x24960, x24959);
  not i24962(x24962, x24961);
  not i24964(x24964, x24963);
  not i24966(x24966, x24965);
  not i24968(x24968, x24967);
  not i24970(x24970, x24969);
  not i24972(x24972, x24971);
  not i24974(x24974, x24973);
  not i24976(x24976, x24975);
  not i24978(x24978, x24977);
  not i24980(x24980, x24979);
  not i24982(x24982, x24981);
  not i24984(x24984, x24983);
  not i24986(x24986, x24985);
  not i24988(x24988, x24987);
  not i25749(x25749, x71982);
  not i25772(x25772, x71987);
  not i25782(x25782, x71992);
  not i25790(x25790, x71997);
  not i25796(x25796, x72002);
  not i27944(x27944, x27881);
  not i27945(x27945, x27883);
  not i27946(x27946, x27885);
  not i27947(x27947, x27887);
  not i27948(x27948, x27889);
  not i27949(x27949, x27891);
  not i27950(x27950, x27893);
  not i27951(x27951, x27895);
  not i27952(x27952, x27897);
  not i27953(x27953, x27899);
  not i27954(x27954, x27901);
  not i27955(x27955, x27903);
  not i27956(x27956, x27905);
  not i27957(x27957, x27907);
  not i27958(x27958, x27909);
  not i27959(x27959, x27911);
  not i27960(x27960, x27913);
  not i27961(x27961, x27915);
  not i27962(x27962, x27917);
  not i27963(x27963, x27919);
  not i27964(x27964, x27921);
  not i27965(x27965, x27923);
  not i27966(x27966, x27925);
  not i27967(x27967, x27927);
  not i27968(x27968, x27929);
  not i27969(x27969, x27931);
  not i27970(x27970, x27933);
  not i27971(x27971, x27935);
  not i27972(x27972, x27937);
  not i27973(x27973, x27939);
  not i27974(x27974, x27941);
  not i27975(x27975, x27943);
  not i28073(x28073, x27978);
  not i28074(x28074, x72537);
  not i28077(x28077, x28076);
  not i28079(x28079, x27981);
  not i28080(x28080, x72542);
  not i28083(x28083, x28082);
  not i28085(x28085, x27984);
  not i28086(x28086, x72547);
  not i28089(x28089, x28088);
  not i28091(x28091, x27987);
  not i28092(x28092, x72552);
  not i28095(x28095, x28094);
  not i28097(x28097, x27990);
  not i28098(x28098, x72557);
  not i28101(x28101, x28100);
  not i28103(x28103, x27993);
  not i28104(x28104, x72562);
  not i28107(x28107, x28106);
  not i28109(x28109, x27996);
  not i28110(x28110, x72567);
  not i28113(x28113, x28112);
  not i28115(x28115, x27999);
  not i28116(x28116, x72572);
  not i28119(x28119, x28118);
  not i28121(x28121, x28002);
  not i28122(x28122, x72577);
  not i28125(x28125, x28124);
  not i28127(x28127, x28005);
  not i28128(x28128, x72582);
  not i28131(x28131, x28130);
  not i28133(x28133, x28008);
  not i28134(x28134, x72587);
  not i28137(x28137, x28136);
  not i28139(x28139, x28011);
  not i28140(x28140, x72592);
  not i28143(x28143, x28142);
  not i28145(x28145, x28014);
  not i28146(x28146, x72597);
  not i28149(x28149, x28148);
  not i28151(x28151, x28017);
  not i28152(x28152, x72602);
  not i28155(x28155, x28154);
  not i28157(x28157, x28020);
  not i28158(x28158, x72607);
  not i28161(x28161, x28160);
  not i28163(x28163, x28023);
  not i28164(x28164, x72612);
  not i28167(x28167, x28166);
  not i28169(x28169, x28026);
  not i28170(x28170, x72617);
  not i28173(x28173, x28172);
  not i28175(x28175, x28029);
  not i28176(x28176, x72622);
  not i28179(x28179, x28178);
  not i28181(x28181, x28032);
  not i28182(x28182, x72627);
  not i28185(x28185, x28184);
  not i28187(x28187, x28035);
  not i28188(x28188, x72632);
  not i28191(x28191, x28190);
  not i28193(x28193, x28038);
  not i28194(x28194, x72637);
  not i28197(x28197, x28196);
  not i28199(x28199, x28041);
  not i28200(x28200, x72642);
  not i28203(x28203, x28202);
  not i28205(x28205, x28044);
  not i28206(x28206, x72647);
  not i28209(x28209, x28208);
  not i28211(x28211, x28047);
  not i28212(x28212, x72652);
  not i28215(x28215, x28214);
  not i28217(x28217, x28050);
  not i28218(x28218, x72657);
  not i28221(x28221, x28220);
  not i28223(x28223, x28053);
  not i28224(x28224, x72662);
  not i28227(x28227, x28226);
  not i28229(x28229, x28056);
  not i28230(x28230, x72667);
  not i28233(x28233, x28232);
  not i28235(x28235, x28059);
  not i28236(x28236, x72672);
  not i28239(x28239, x28238);
  not i28241(x28241, x28062);
  not i28242(x28242, x72677);
  not i28245(x28245, x28244);
  not i28247(x28247, x28065);
  not i28248(x28248, x72682);
  not i28251(x28251, x28250);
  not i28253(x28253, x28068);
  not i28254(x28254, x72687);
  not i28257(x28257, x28256);
  not i28259(x28259, x28071);
  not i28260(x28260, x72692);
  not i28263(x28263, x28262);
  not i28264(x28264, x28072);
  not i28265(x28265, x28078);
  not i28266(x28266, x28084);
  not i28267(x28267, x28090);
  not i28268(x28268, x28096);
  not i28269(x28269, x28102);
  not i28270(x28270, x28108);
  not i28271(x28271, x28114);
  not i28272(x28272, x28120);
  not i28273(x28273, x28126);
  not i28274(x28274, x28132);
  not i28275(x28275, x28138);
  not i28276(x28276, x28144);
  not i28277(x28277, x28150);
  not i28278(x28278, x28156);
  not i28279(x28279, x28162);
  not i28280(x28280, x28168);
  not i28281(x28281, x28174);
  not i28282(x28282, x28180);
  not i28283(x28283, x28186);
  not i28284(x28284, x28192);
  not i28285(x28285, x28198);
  not i28286(x28286, x28204);
  not i28287(x28287, x28210);
  not i28288(x28288, x28216);
  not i28289(x28289, x28222);
  not i28290(x28290, x28228);
  not i28291(x28291, x28234);
  not i28292(x28292, x28240);
  not i28293(x28293, x28246);
  not i28299(x28299, x28298);
  not i28303(x28303, x28302);
  not i28307(x28307, x28306);
  not i28311(x28311, x28310);
  not i28315(x28315, x28314);
  not i28319(x28319, x28318);
  not i28323(x28323, x28322);
  not i28327(x28327, x28326);
  not i28331(x28331, x28330);
  not i28335(x28335, x28334);
  not i28339(x28339, x28338);
  not i28343(x28343, x28342);
  not i28347(x28347, x28346);
  not i28351(x28351, x28350);
  not i28355(x28355, x28354);
  not i28359(x28359, x28358);
  not i28363(x28363, x28362);
  not i28367(x28367, x28366);
  not i28371(x28371, x28370);
  not i28375(x28375, x28374);
  not i28379(x28379, x28378);
  not i28383(x28383, x28382);
  not i28387(x28387, x28386);
  not i28391(x28391, x28390);
  not i28395(x28395, x28394);
  not i28399(x28399, x28398);
  not i28403(x28403, x28402);
  not i28407(x28407, x28406);
  not i28411(x28411, x28410);
  not i28415(x28415, x28414);
  not i28417(x28417, x28297);
  not i28420(x28420, x28301);
  not i28423(x28423, x28305);
  not i28426(x28426, x28425);
  not i28428(x28428, x28309);
  not i28431(x28431, x28430);
  not i28433(x28433, x28313);
  not i28436(x28436, x28435);
  not i28438(x28438, x28317);
  not i28441(x28441, x28440);
  not i28443(x28443, x28321);
  not i28446(x28446, x28445);
  not i28448(x28448, x28325);
  not i28451(x28451, x28450);
  not i28453(x28453, x28329);
  not i28456(x28456, x28455);
  not i28458(x28458, x28333);
  not i28461(x28461, x28460);
  not i28463(x28463, x28337);
  not i28466(x28466, x28465);
  not i28468(x28468, x28341);
  not i28471(x28471, x28470);
  not i28473(x28473, x28345);
  not i28476(x28476, x28475);
  not i28478(x28478, x28349);
  not i28481(x28481, x28480);
  not i28483(x28483, x28353);
  not i28486(x28486, x28485);
  not i28488(x28488, x28357);
  not i28491(x28491, x28490);
  not i28493(x28493, x28361);
  not i28496(x28496, x28495);
  not i28498(x28498, x28365);
  not i28501(x28501, x28500);
  not i28503(x28503, x28369);
  not i28506(x28506, x28505);
  not i28508(x28508, x28373);
  not i28511(x28511, x28510);
  not i28513(x28513, x28377);
  not i28516(x28516, x28515);
  not i28518(x28518, x28381);
  not i28521(x28521, x28520);
  not i28523(x28523, x28385);
  not i28526(x28526, x28525);
  not i28528(x28528, x28389);
  not i28531(x28531, x28530);
  not i28533(x28533, x28393);
  not i28536(x28536, x28535);
  not i28538(x28538, x28397);
  not i28541(x28541, x28540);
  not i28543(x28543, x28401);
  not i28546(x28546, x28545);
  not i28548(x28548, x28405);
  not i28551(x28551, x28550);
  not i28553(x28553, x28409);
  not i28556(x28556, x28555);
  not i28558(x28558, x28413);
  not i28561(x28561, x28560);
  not i28563(x28563, x28424);
  not i28566(x28566, x28429);
  not i28569(x28569, x28434);
  not i28572(x28572, x28439);
  not i28575(x28575, x28444);
  not i28578(x28578, x28577);
  not i28580(x28580, x28449);
  not i28583(x28583, x28582);
  not i28585(x28585, x28454);
  not i28588(x28588, x28587);
  not i28590(x28590, x28459);
  not i28593(x28593, x28592);
  not i28595(x28595, x28464);
  not i28598(x28598, x28597);
  not i28600(x28600, x28469);
  not i28603(x28603, x28602);
  not i28605(x28605, x28474);
  not i28608(x28608, x28607);
  not i28610(x28610, x28479);
  not i28613(x28613, x28612);
  not i28615(x28615, x28484);
  not i28618(x28618, x28617);
  not i28620(x28620, x28489);
  not i28623(x28623, x28622);
  not i28625(x28625, x28494);
  not i28628(x28628, x28627);
  not i28630(x28630, x28499);
  not i28633(x28633, x28632);
  not i28635(x28635, x28504);
  not i28638(x28638, x28637);
  not i28640(x28640, x28509);
  not i28643(x28643, x28642);
  not i28645(x28645, x28514);
  not i28648(x28648, x28647);
  not i28650(x28650, x28519);
  not i28653(x28653, x28652);
  not i28655(x28655, x28524);
  not i28658(x28658, x28657);
  not i28660(x28660, x28529);
  not i28663(x28663, x28662);
  not i28665(x28665, x28534);
  not i28668(x28668, x28667);
  not i28670(x28670, x28539);
  not i28673(x28673, x28672);
  not i28675(x28675, x28544);
  not i28678(x28678, x28677);
  not i28680(x28680, x28549);
  not i28683(x28683, x28682);
  not i28685(x28685, x28554);
  not i28688(x28688, x28687);
  not i28690(x28690, x28559);
  not i28693(x28693, x28692);
  not i28695(x28695, x28576);
  not i28698(x28698, x28581);
  not i28701(x28701, x28586);
  not i28704(x28704, x28591);
  not i28707(x28707, x28596);
  not i28710(x28710, x28601);
  not i28713(x28713, x28606);
  not i28716(x28716, x28611);
  not i28719(x28719, x28616);
  not i28722(x28722, x28721);
  not i28724(x28724, x28621);
  not i28727(x28727, x28726);
  not i28729(x28729, x28626);
  not i28732(x28732, x28731);
  not i28734(x28734, x28631);
  not i28737(x28737, x28736);
  not i28739(x28739, x28636);
  not i28742(x28742, x28741);
  not i28744(x28744, x28641);
  not i28747(x28747, x28746);
  not i28749(x28749, x28646);
  not i28752(x28752, x28751);
  not i28754(x28754, x28651);
  not i28757(x28757, x28756);
  not i28759(x28759, x28656);
  not i28762(x28762, x28761);
  not i28764(x28764, x28661);
  not i28767(x28767, x28766);
  not i28769(x28769, x28666);
  not i28772(x28772, x28771);
  not i28774(x28774, x28671);
  not i28777(x28777, x28776);
  not i28779(x28779, x28676);
  not i28782(x28782, x28781);
  not i28784(x28784, x28681);
  not i28787(x28787, x28786);
  not i28789(x28789, x28686);
  not i28792(x28792, x28791);
  not i28794(x28794, x28691);
  not i28797(x28797, x28796);
  not i28799(x28799, x28720);
  not i28802(x28802, x28725);
  not i28805(x28805, x28730);
  not i28808(x28808, x28735);
  not i28811(x28811, x28740);
  not i28814(x28814, x28745);
  not i28817(x28817, x28750);
  not i28820(x28820, x28755);
  not i28823(x28823, x28760);
  not i28826(x28826, x28765);
  not i28829(x28829, x28770);
  not i28832(x28832, x28775);
  not i28835(x28835, x28780);
  not i28838(x28838, x28785);
  not i28841(x28841, x28790);
  not i28844(x28844, x28795);
  not i28848(x28848, x28847);
  not i28850(x28850, x28295);
  not i28853(x28853, x28852);
  not i28855(x28855, x28418);
  not i28858(x28858, x28857);
  not i28860(x28860, x28421);
  not i28863(x28863, x28862);
  not i28865(x28865, x28564);
  not i28868(x28868, x28867);
  not i28870(x28870, x28567);
  not i28873(x28873, x28872);
  not i28875(x28875, x28570);
  not i28878(x28878, x28877);
  not i28880(x28880, x28573);
  not i28883(x28883, x28882);
  not i28885(x28885, x28696);
  not i28888(x28888, x28887);
  not i28890(x28890, x28699);
  not i28893(x28893, x28892);
  not i28895(x28895, x28702);
  not i28898(x28898, x28897);
  not i28900(x28900, x28705);
  not i28903(x28903, x28902);
  not i28905(x28905, x28708);
  not i28908(x28908, x28907);
  not i28910(x28910, x28711);
  not i28913(x28913, x28912);
  not i28915(x28915, x28714);
  not i28918(x28918, x28917);
  not i28920(x28920, x28717);
  not i28923(x28923, x28922);
  not i28925(x28925, x28800);
  not i28928(x28928, x28927);
  not i28930(x28930, x28803);
  not i28933(x28933, x28932);
  not i28935(x28935, x28806);
  not i28938(x28938, x28937);
  not i28940(x28940, x28809);
  not i28943(x28943, x28942);
  not i28945(x28945, x28812);
  not i28948(x28948, x28947);
  not i28950(x28950, x28815);
  not i28953(x28953, x28952);
  not i28955(x28955, x28818);
  not i28958(x28958, x28957);
  not i28960(x28960, x28821);
  not i28963(x28963, x28962);
  not i28965(x28965, x28824);
  not i28968(x28968, x28967);
  not i28970(x28970, x28827);
  not i28973(x28973, x28972);
  not i28975(x28975, x28830);
  not i28978(x28978, x28977);
  not i28980(x28980, x28833);
  not i28983(x28983, x28982);
  not i28985(x28985, x28836);
  not i28988(x28988, x28987);
  not i28990(x28990, x28839);
  not i28993(x28993, x28992);
  not i28995(x28995, x28842);
  not i28998(x28998, x28997);
  not i29000(x29000, x28845);
  not i29003(x29003, x29002);
  not i29006(x29006, x29005);
  not i29008(x29008, x29007);
  not i29010(x29010, x29009);
  not i29012(x29012, x29011);
  not i29014(x29014, x29013);
  not i29016(x29016, x29015);
  not i29018(x29018, x29017);
  not i29020(x29020, x29019);
  not i29023(x29023, x29022);
  not i29025(x29025, x29024);
  not i29027(x29027, x29026);
  not i29029(x29029, x29028);
  not i29031(x29031, x29030);
  not i29033(x29033, x29032);
  not i29035(x29035, x29034);
  not i29037(x29037, x29036);
  not i29039(x29039, x29038);
  not i29041(x29041, x29040);
  not i29043(x29043, x29042);
  not i29045(x29045, x29044);
  not i29047(x29047, x29046);
  not i29049(x29049, x29048);
  not i29051(x29051, x29050);
  not i29053(x29053, x29052);
  not i29055(x29055, x29054);
  not i29058(x29058, x29057);
  not i29060(x29060, x29059);
  not i29062(x29062, x29061);
  not i29064(x29064, x29063);
  not i29066(x29066, x29065);
  not i29068(x29068, x29067);
  not i29070(x29070, x29069);
  not i29072(x29072, x29071);
  not i29074(x29074, x29073);
  not i29076(x29076, x29075);
  not i29078(x29078, x29077);
  not i29080(x29080, x29079);
  not i29082(x29082, x29081);
  not i29084(x29084, x29083);
  not i29086(x29086, x29085);
  not i29088(x29088, x29087);
  not i29090(x29090, x29089);
  not i29092(x29092, x29091);
  not i29094(x29094, x29093);
  not i29096(x29096, x29095);
  not i29098(x29098, x29097);
  not i29100(x29100, x29099);
  not i29102(x29102, x29101);
  not i29104(x29104, x29103);
  not i29106(x29106, x29105);
  not i29108(x29108, x29107);
  not i29111(x29111, x29110);
  not i29113(x29113, x29112);
  not i29115(x29115, x29114);
  not i29117(x29117, x29116);
  not i29119(x29119, x29118);
  not i29121(x29121, x29120);
  not i29123(x29123, x29122);
  not i29125(x29125, x29124);
  not i29127(x29127, x29126);
  not i29129(x29129, x29128);
  not i29131(x29131, x29130);
  not i29133(x29133, x29132);
  not i29135(x29135, x29134);
  not i29137(x29137, x29136);
  not i29139(x29139, x29138);
  not i29141(x29141, x29140);
  not i29143(x29143, x29142);
  not i29145(x29145, x29144);
  not i29147(x29147, x29146);
  not i29149(x29149, x29148);
  not i29151(x29151, x29150);
  not i29153(x29153, x29152);
  not i29155(x29155, x29154);
  not i29157(x29157, x29156);
  not i29159(x29159, x29158);
  not i29161(x29161, x29160);
  not i29163(x29163, x29162);
  not i29165(x29165, x29164);
  not i29167(x29167, x29166);
  not i29169(x29169, x29168);
  not i29171(x29171, x29170);
  not i29173(x29173, x29172);
  not i29175(x29175, x29174);
  not i29177(x29177, x29176);
  not i29179(x29179, x29178);
  not i29182(x29182, x29181);
  not i29184(x29184, x29183);
  not i29186(x29186, x29185);
  not i29188(x29188, x29187);
  not i29190(x29190, x29189);
  not i29192(x29192, x29191);
  not i29194(x29194, x29193);
  not i29196(x29196, x29195);
  not i29198(x29198, x29197);
  not i29200(x29200, x29199);
  not i29202(x29202, x29201);
  not i29204(x29204, x29203);
  not i29206(x29206, x29205);
  not i29208(x29208, x29207);
  not i29210(x29210, x29209);
  not i29212(x29212, x29211);
  not i29214(x29214, x29213);
  not i29216(x29216, x29215);
  not i29218(x29218, x29217);
  not i29220(x29220, x29219);
  not i29222(x29222, x29221);
  not i29224(x29224, x29223);
  not i29226(x29226, x29225);
  not i29228(x29228, x29227);
  not i29230(x29230, x29229);
  not i29232(x29232, x29231);
  not i29234(x29234, x29233);
  not i29236(x29236, x29235);
  not i29238(x29238, x29237);
  not i29240(x29240, x29239);
  not i29242(x29242, x29241);
  not i29244(x29244, x29243);
  not i29246(x29246, x29245);
  not i29248(x29248, x29247);
  not i29250(x29250, x29249);
  not i29252(x29252, x29251);
  not i29254(x29254, x29253);
  not i29256(x29256, x29255);
  not i29258(x29258, x29257);
  not i29260(x29260, x29259);
  not i29262(x29262, x29261);
  not i29264(x29264, x29263);
  not i29266(x29266, x29265);
  not i29268(x29268, x29267);
  not i29271(x29271, x29270);
  not i29273(x29273, x29272);
  not i29275(x29275, x29274);
  not i29277(x29277, x29276);
  not i29279(x29279, x29278);
  not i29281(x29281, x29280);
  not i29283(x29283, x29282);
  not i29285(x29285, x29284);
  not i29287(x29287, x29286);
  not i29289(x29289, x29288);
  not i29291(x29291, x29290);
  not i29293(x29293, x29292);
  not i29295(x29295, x29294);
  not i29297(x29297, x29296);
  not i29299(x29299, x29298);
  not i29301(x29301, x29300);
  not i29303(x29303, x29302);
  not i29305(x29305, x29304);
  not i29307(x29307, x29306);
  not i29309(x29309, x29308);
  not i29311(x29311, x29310);
  not i29313(x29313, x29312);
  not i29315(x29315, x29314);
  not i29317(x29317, x29316);
  not i29319(x29319, x29318);
  not i29321(x29321, x29320);
  not i29323(x29323, x29322);
  not i29325(x29325, x29324);
  not i29327(x29327, x29326);
  not i29329(x29329, x29328);
  not i29331(x29331, x29330);
  not i29333(x29333, x29332);
  not i29335(x29335, x29334);
  not i29337(x29337, x29336);
  not i29339(x29339, x29338);
  not i29341(x29341, x29340);
  not i29343(x29343, x29342);
  not i29345(x29345, x29344);
  not i29347(x29347, x29346);
  not i29349(x29349, x29348);
  not i29351(x29351, x29350);
  not i29353(x29353, x29352);
  not i29355(x29355, x29354);
  not i29357(x29357, x29356);
  not i29359(x29359, x29358);
  not i29361(x29361, x29360);
  not i29363(x29363, x29362);
  not i29365(x29365, x29364);
  not i29367(x29367, x29366);
  not i29369(x29369, x29368);
  not i29371(x29371, x29370);
  not i29373(x29373, x29372);
  not i29375(x29375, x29374);
  not i29378(x29378, x29377);
  not i29380(x29380, x29379);
  not i29382(x29382, x29381);
  not i29384(x29384, x29383);
  not i29386(x29386, x29385);
  not i29388(x29388, x29387);
  not i29390(x29390, x29389);
  not i29392(x29392, x29391);
  not i29394(x29394, x29393);
  not i29396(x29396, x29395);
  not i29398(x29398, x29397);
  not i29400(x29400, x29399);
  not i29402(x29402, x29401);
  not i29404(x29404, x29403);
  not i29406(x29406, x29405);
  not i29408(x29408, x29407);
  not i29410(x29410, x29409);
  not i29412(x29412, x29411);
  not i29414(x29414, x29413);
  not i29416(x29416, x29415);
  not i29418(x29418, x29417);
  not i29420(x29420, x29419);
  not i29422(x29422, x29421);
  not i29424(x29424, x29423);
  not i29426(x29426, x29425);
  not i29428(x29428, x29427);
  not i29430(x29430, x29429);
  not i29432(x29432, x29431);
  not i29434(x29434, x29433);
  not i29436(x29436, x29435);
  not i29438(x29438, x29437);
  not i29440(x29440, x29439);
  not i29442(x29442, x29441);
  not i29444(x29444, x29443);
  not i29446(x29446, x29445);
  not i29448(x29448, x29447);
  not i29450(x29450, x29449);
  not i29452(x29452, x29451);
  not i29454(x29454, x29453);
  not i29456(x29456, x29455);
  not i29458(x29458, x29457);
  not i29460(x29460, x29459);
  not i29462(x29462, x29461);
  not i29464(x29464, x29463);
  not i29466(x29466, x29465);
  not i29468(x29468, x29467);
  not i29470(x29470, x29469);
  not i29472(x29472, x29471);
  not i29474(x29474, x29473);
  not i29476(x29476, x29475);
  not i29478(x29478, x29477);
  not i29480(x29480, x29479);
  not i29482(x29482, x29481);
  not i29484(x29484, x29483);
  not i29486(x29486, x29485);
  not i29488(x29488, x29487);
  not i29490(x29490, x29489);
  not i29492(x29492, x29491);
  not i29494(x29494, x29493);
  not i29496(x29496, x29495);
  not i29498(x29498, x29497);
  not i29500(x29500, x29499);
  not i29503(x29503, x29502);
  not i29505(x29505, x29504);
  not i29507(x29507, x29506);
  not i29509(x29509, x29508);
  not i29511(x29511, x29510);
  not i29513(x29513, x29512);
  not i29515(x29515, x29514);
  not i29517(x29517, x29516);
  not i29519(x29519, x29518);
  not i29521(x29521, x29520);
  not i29523(x29523, x29522);
  not i29525(x29525, x29524);
  not i29527(x29527, x29526);
  not i29529(x29529, x29528);
  not i29531(x29531, x29530);
  not i29533(x29533, x29532);
  not i29535(x29535, x29534);
  not i29537(x29537, x29536);
  not i29539(x29539, x29538);
  not i29541(x29541, x29540);
  not i29543(x29543, x29542);
  not i29545(x29545, x29544);
  not i29547(x29547, x29546);
  not i29549(x29549, x29548);
  not i29551(x29551, x29550);
  not i29553(x29553, x29552);
  not i29555(x29555, x29554);
  not i29557(x29557, x29556);
  not i29559(x29559, x29558);
  not i29561(x29561, x29560);
  not i29563(x29563, x29562);
  not i29565(x29565, x29564);
  not i29567(x29567, x29566);
  not i29569(x29569, x29568);
  not i29571(x29571, x29570);
  not i29573(x29573, x29572);
  not i29575(x29575, x29574);
  not i29577(x29577, x29576);
  not i29579(x29579, x29578);
  not i29581(x29581, x29580);
  not i29583(x29583, x29582);
  not i29585(x29585, x29584);
  not i29587(x29587, x29586);
  not i29589(x29589, x29588);
  not i29591(x29591, x29590);
  not i29593(x29593, x29592);
  not i29595(x29595, x29594);
  not i29597(x29597, x29596);
  not i29599(x29599, x29598);
  not i29601(x29601, x29600);
  not i29603(x29603, x29602);
  not i29605(x29605, x29604);
  not i29607(x29607, x29606);
  not i29609(x29609, x29608);
  not i29611(x29611, x29610);
  not i29613(x29613, x29612);
  not i29615(x29615, x29614);
  not i29617(x29617, x29616);
  not i29619(x29619, x29618);
  not i29621(x29621, x29620);
  not i29623(x29623, x29622);
  not i29625(x29625, x29624);
  not i29627(x29627, x29626);
  not i29629(x29629, x29628);
  not i29631(x29631, x29630);
  not i29633(x29633, x29632);
  not i29635(x29635, x29634);
  not i29637(x29637, x29636);
  not i29639(x29639, x29638);
  not i29641(x29641, x29640);
  not i29643(x29643, x29642);
  not i29646(x29646, x29645);
  not i29648(x29648, x29647);
  not i29650(x29650, x29649);
  not i29652(x29652, x29651);
  not i29654(x29654, x29653);
  not i29656(x29656, x29655);
  not i29658(x29658, x29657);
  not i29660(x29660, x29659);
  not i29662(x29662, x29661);
  not i29664(x29664, x29663);
  not i29666(x29666, x29665);
  not i29668(x29668, x29667);
  not i29670(x29670, x29669);
  not i29672(x29672, x29671);
  not i29674(x29674, x29673);
  not i29676(x29676, x29675);
  not i29678(x29678, x29677);
  not i29680(x29680, x29679);
  not i29682(x29682, x29681);
  not i29684(x29684, x29683);
  not i29686(x29686, x29685);
  not i29688(x29688, x29687);
  not i29690(x29690, x29689);
  not i29692(x29692, x29691);
  not i29694(x29694, x29693);
  not i29696(x29696, x29695);
  not i29698(x29698, x29697);
  not i29700(x29700, x29699);
  not i29702(x29702, x29701);
  not i29704(x29704, x29703);
  not i29706(x29706, x29705);
  not i29708(x29708, x29707);
  not i29710(x29710, x29709);
  not i29712(x29712, x29711);
  not i29714(x29714, x29713);
  not i29716(x29716, x29715);
  not i29718(x29718, x29717);
  not i29720(x29720, x29719);
  not i29722(x29722, x29721);
  not i29724(x29724, x29723);
  not i29726(x29726, x29725);
  not i29728(x29728, x29727);
  not i29730(x29730, x29729);
  not i29732(x29732, x29731);
  not i29734(x29734, x29733);
  not i29736(x29736, x29735);
  not i29738(x29738, x29737);
  not i29740(x29740, x29739);
  not i29742(x29742, x29741);
  not i29744(x29744, x29743);
  not i29746(x29746, x29745);
  not i29748(x29748, x29747);
  not i29750(x29750, x29749);
  not i29752(x29752, x29751);
  not i29754(x29754, x29753);
  not i29756(x29756, x29755);
  not i29758(x29758, x29757);
  not i29760(x29760, x29759);
  not i29762(x29762, x29761);
  not i29764(x29764, x29763);
  not i29766(x29766, x29765);
  not i29768(x29768, x29767);
  not i29770(x29770, x29769);
  not i29772(x29772, x29771);
  not i29774(x29774, x29773);
  not i29776(x29776, x29775);
  not i29778(x29778, x29777);
  not i29780(x29780, x29779);
  not i29782(x29782, x29781);
  not i29784(x29784, x29783);
  not i29786(x29786, x29785);
  not i29788(x29788, x29787);
  not i29790(x29790, x29789);
  not i29792(x29792, x29791);
  not i29794(x29794, x29793);
  not i29796(x29796, x29795);
  not i29798(x29798, x29797);
  not i29800(x29800, x29799);
  not i29802(x29802, x29801);
  not i29804(x29804, x29803);
  not i29807(x29807, x29806);
  not i29809(x29809, x29808);
  not i29811(x29811, x29810);
  not i29813(x29813, x29812);
  not i29815(x29815, x29814);
  not i29817(x29817, x29816);
  not i29819(x29819, x29818);
  not i29821(x29821, x29820);
  not i29823(x29823, x29822);
  not i29825(x29825, x29824);
  not i29827(x29827, x29826);
  not i29829(x29829, x29828);
  not i29831(x29831, x29830);
  not i29833(x29833, x29832);
  not i29835(x29835, x29834);
  not i29837(x29837, x29836);
  not i29839(x29839, x29838);
  not i29841(x29841, x29840);
  not i29843(x29843, x29842);
  not i29845(x29845, x29844);
  not i29847(x29847, x29846);
  not i29849(x29849, x29848);
  not i29851(x29851, x29850);
  not i29853(x29853, x29852);
  not i29855(x29855, x29854);
  not i29857(x29857, x29856);
  not i29859(x29859, x29858);
  not i29861(x29861, x29860);
  not i29863(x29863, x29862);
  not i29865(x29865, x29864);
  not i29867(x29867, x29866);
  not i29869(x29869, x29868);
  not i29871(x29871, x29870);
  not i29873(x29873, x29872);
  not i29875(x29875, x29874);
  not i29877(x29877, x29876);
  not i29879(x29879, x29878);
  not i29881(x29881, x29880);
  not i29883(x29883, x29882);
  not i29885(x29885, x29884);
  not i29887(x29887, x29886);
  not i29889(x29889, x29888);
  not i29891(x29891, x29890);
  not i29893(x29893, x29892);
  not i29895(x29895, x29894);
  not i29897(x29897, x29896);
  not i29899(x29899, x29898);
  not i29901(x29901, x29900);
  not i29903(x29903, x29902);
  not i29905(x29905, x29904);
  not i29907(x29907, x29906);
  not i29909(x29909, x29908);
  not i29911(x29911, x29910);
  not i29913(x29913, x29912);
  not i29915(x29915, x29914);
  not i29917(x29917, x29916);
  not i29919(x29919, x29918);
  not i29921(x29921, x29920);
  not i29923(x29923, x29922);
  not i29925(x29925, x29924);
  not i29927(x29927, x29926);
  not i29929(x29929, x29928);
  not i29931(x29931, x29930);
  not i29933(x29933, x29932);
  not i29935(x29935, x29934);
  not i29937(x29937, x29936);
  not i29939(x29939, x29938);
  not i29941(x29941, x29940);
  not i29943(x29943, x29942);
  not i29945(x29945, x29944);
  not i29947(x29947, x29946);
  not i29949(x29949, x29948);
  not i29951(x29951, x29950);
  not i29953(x29953, x29952);
  not i29955(x29955, x29954);
  not i29957(x29957, x29956);
  not i29959(x29959, x29958);
  not i29961(x29961, x29960);
  not i29963(x29963, x29962);
  not i29965(x29965, x29964);
  not i29967(x29967, x29966);
  not i29969(x29969, x29968);
  not i29971(x29971, x29970);
  not i29973(x29973, x29972);
  not i29975(x29975, x29974);
  not i29977(x29977, x29976);
  not i29979(x29979, x29978);
  not i29981(x29981, x29980);
  not i29983(x29983, x29982);
  not i29986(x29986, x29985);
  not i29988(x29988, x29987);
  not i29990(x29990, x29989);
  not i29992(x29992, x29991);
  not i29994(x29994, x29993);
  not i29996(x29996, x29995);
  not i29998(x29998, x29997);
  not i30000(x30000, x29999);
  not i30002(x30002, x30001);
  not i30004(x30004, x30003);
  not i30006(x30006, x30005);
  not i30008(x30008, x30007);
  not i30010(x30010, x30009);
  not i30012(x30012, x30011);
  not i30014(x30014, x30013);
  not i30016(x30016, x30015);
  not i30018(x30018, x30017);
  not i30020(x30020, x30019);
  not i30022(x30022, x30021);
  not i30024(x30024, x30023);
  not i30026(x30026, x30025);
  not i30028(x30028, x30027);
  not i30030(x30030, x30029);
  not i30032(x30032, x30031);
  not i30034(x30034, x30033);
  not i30036(x30036, x30035);
  not i30038(x30038, x30037);
  not i30040(x30040, x30039);
  not i30042(x30042, x30041);
  not i30044(x30044, x30043);
  not i30046(x30046, x30045);
  not i30048(x30048, x30047);
  not i30055(x30055, x30054);
  not i30063(x30063, x30062);
  not i30071(x30071, x30070);
  not i30082(x30082, x30081);
  not i30090(x30090, x30089);
  not i30098(x30098, x30097);
  not i30106(x30106, x30105);
  not i30110(x30110, x30109);
  not i30115(x30115, x30114);
  not i30123(x30123, x30122);
  not i30127(x30127, x30126);
  not i30135(x30135, x30134);
  not i30143(x30143, x30142);
  not i30147(x30147, x30146);
  not i30152(x30152, x30151);
  not i30156(x30156, x30155);
  not i30161(x30161, x30160);
  not i30169(x30169, x30168);
  not i30173(x30173, x30172);
  not i30178(x30178, x30177);
  not i30182(x30182, x30181);
  not i30187(x30187, x30186);
  not i30195(x30195, x30194);
  not i30199(x30199, x30198);
  not i30204(x30204, x30203);
  not i30208(x30208, x30207);
  not i30216(x30216, x30215);
  not i30224(x30224, x30223);
  not i30228(x30228, x30227);
  not i30233(x30233, x30232);
  not i30237(x30237, x30236);
  not i30242(x30242, x30241);
  not i30246(x30246, x30245);
  not i30251(x30251, x30250);
  not i30259(x30259, x30258);
  not i30263(x30263, x30262);
  not i30268(x30268, x30267);
  not i30272(x30272, x30271);
  not i30277(x30277, x30276);
  not i30281(x30281, x30280);
  not i30286(x30286, x30285);
  not i30294(x30294, x30293);
  not i30298(x30298, x30297);
  not i30303(x30303, x30302);
  not i30307(x30307, x30306);
  not i30312(x30312, x30311);
  not i30316(x30316, x30315);
  not i30324(x30324, x30323);
  not i30332(x30332, x30331);
  not i30336(x30336, x30335);
  not i30341(x30341, x30340);
  not i30345(x30345, x30344);
  not i30350(x30350, x30349);
  not i30354(x30354, x30353);
  not i30359(x30359, x30358);
  not i30367(x30367, x30366);
  not i30375(x30375, x30374);
  not i30379(x30379, x30378);
  not i30384(x30384, x30383);
  not i30388(x30388, x30387);
  not i30393(x30393, x30392);
  not i30397(x30397, x30396);
  not i30402(x30402, x30401);
  not i30406(x30406, x30405);
  not i30411(x30411, x30410);
  not i30419(x30419, x30418);
  not i30423(x30423, x30422);
  not i30428(x30428, x30427);
  not i30432(x30432, x30431);
  not i30437(x30437, x30436);
  not i30441(x30441, x30440);
  not i30446(x30446, x30445);
  not i30450(x30450, x30449);
  not i30458(x30458, x30457);
  not i30466(x30466, x30465);
  not i30470(x30470, x30469);
  not i30475(x30475, x30474);
  not i30479(x30479, x30478);
  not i30484(x30484, x30483);
  not i30488(x30488, x30487);
  not i30493(x30493, x30492);
  not i30497(x30497, x30496);
  not i30502(x30502, x30501);
  not i30506(x30506, x30505);
  not i30511(x30511, x30510);
  not i30519(x30519, x30518);
  not i30523(x30523, x30522);
  not i30528(x30528, x30527);
  not i30532(x30532, x30531);
  not i30537(x30537, x30536);
  not i30541(x30541, x30540);
  not i30546(x30546, x30545);
  not i30550(x30550, x30549);
  not i30555(x30555, x30554);
  not i30559(x30559, x30558);
  not i30564(x30564, x30563);
  not i30572(x30572, x30571);
  not i30576(x30576, x30575);
  not i30581(x30581, x30580);
  not i30585(x30585, x30584);
  not i30590(x30590, x30589);
  not i30594(x30594, x30593);
  not i30599(x30599, x30598);
  not i30603(x30603, x30602);
  not i30608(x30608, x30607);
  not i30612(x30612, x30611);
  not i30620(x30620, x30619);
  not i30628(x30628, x30627);
  not i30632(x30632, x30631);
  not i30637(x30637, x30636);
  not i30641(x30641, x30640);
  not i30646(x30646, x30645);
  not i30650(x30650, x30649);
  not i30655(x30655, x30654);
  not i30659(x30659, x30658);
  not i30664(x30664, x30663);
  not i30668(x30668, x30667);
  not i30673(x30673, x30672);
  not i30677(x30677, x30676);
  not i30682(x30682, x30681);
  not i30690(x30690, x30689);
  not i30694(x30694, x30693);
  not i30699(x30699, x30698);
  not i30703(x30703, x30702);
  not i30708(x30708, x30707);
  not i30712(x30712, x30711);
  not i30717(x30717, x30716);
  not i30721(x30721, x30720);
  not i30726(x30726, x30725);
  not i30730(x30730, x30729);
  not i30735(x30735, x30734);
  not i30739(x30739, x30738);
  not i30744(x30744, x30743);
  not i30752(x30752, x30751);
  not i30756(x30756, x30755);
  not i30761(x30761, x30760);
  not i30765(x30765, x30764);
  not i30770(x30770, x30769);
  not i30774(x30774, x30773);
  not i30779(x30779, x30778);
  not i30783(x30783, x30782);
  not i30788(x30788, x30787);
  not i30792(x30792, x30791);
  not i30797(x30797, x30796);
  not i30801(x30801, x30800);
  not i30809(x30809, x30808);
  not i30817(x30817, x30816);
  not i30821(x30821, x30820);
  not i30826(x30826, x30825);
  not i30830(x30830, x30829);
  not i30835(x30835, x30834);
  not i30839(x30839, x30838);
  not i30844(x30844, x30843);
  not i30848(x30848, x30847);
  not i30853(x30853, x30852);
  not i30857(x30857, x30856);
  not i30862(x30862, x30861);
  not i30866(x30866, x30865);
  not i30871(x30871, x30870);
  not i30879(x30879, x30878);
  not i30887(x30887, x30886);
  not i30891(x30891, x30890);
  not i30896(x30896, x30895);
  not i30900(x30900, x30899);
  not i30905(x30905, x30904);
  not i30909(x30909, x30908);
  not i30914(x30914, x30913);
  not i30918(x30918, x30917);
  not i30923(x30923, x30922);
  not i30927(x30927, x30926);
  not i30932(x30932, x30931);
  not i30936(x30936, x30935);
  not i30941(x30941, x30940);
  not i30945(x30945, x30944);
  not i30950(x30950, x30949);
  not i30958(x30958, x30957);
  not i30962(x30962, x30961);
  not i30967(x30967, x30966);
  not i30971(x30971, x30970);
  not i30976(x30976, x30975);
  not i30980(x30980, x30979);
  not i30985(x30985, x30984);
  not i30989(x30989, x30988);
  not i30994(x30994, x30993);
  not i30998(x30998, x30997);
  not i31003(x31003, x31002);
  not i31007(x31007, x31006);
  not i31012(x31012, x31011);
  not i31016(x31016, x31015);
  not i31024(x31024, x31023);
  not i31032(x31032, x31031);
  not i31036(x31036, x31035);
  not i31041(x31041, x31040);
  not i31045(x31045, x31044);
  not i31050(x31050, x31049);
  not i31054(x31054, x31053);
  not i31059(x31059, x31058);
  not i31063(x31063, x31062);
  not i31068(x31068, x31067);
  not i31072(x31072, x31071);
  not i31077(x31077, x31076);
  not i31081(x31081, x31080);
  not i31086(x31086, x31085);
  not i31090(x31090, x31089);
  not i31095(x31095, x31094);
  not i31099(x31099, x31098);
  not i31104(x31104, x31103);
  not i31112(x31112, x31111);
  not i31116(x31116, x31115);
  not i31121(x31121, x31120);
  not i31125(x31125, x31124);
  not i31130(x31130, x31129);
  not i31134(x31134, x31133);
  not i31139(x31139, x31138);
  not i31143(x31143, x31142);
  not i31148(x31148, x31147);
  not i31152(x31152, x31151);
  not i31157(x31157, x31156);
  not i31161(x31161, x31160);
  not i31166(x31166, x31165);
  not i31170(x31170, x31169);
  not i31175(x31175, x31174);
  not i31179(x31179, x31178);
  not i31184(x31184, x31183);
  not i31192(x31192, x31191);
  not i31196(x31196, x31195);
  not i31201(x31201, x31200);
  not i31205(x31205, x31204);
  not i31210(x31210, x31209);
  not i31214(x31214, x31213);
  not i31219(x31219, x31218);
  not i31223(x31223, x31222);
  not i31228(x31228, x31227);
  not i31232(x31232, x31231);
  not i31237(x31237, x31236);
  not i31241(x31241, x31240);
  not i31246(x31246, x31245);
  not i31250(x31250, x31249);
  not i31255(x31255, x31254);
  not i31259(x31259, x31258);
  not i31267(x31267, x31266);
  not i31271(x31271, x31270);
  not i31276(x31276, x31275);
  not i31280(x31280, x31279);
  not i31285(x31285, x31284);
  not i31289(x31289, x31288);
  not i31294(x31294, x31293);
  not i31298(x31298, x31297);
  not i31303(x31303, x31302);
  not i31307(x31307, x31306);
  not i31312(x31312, x31311);
  not i31316(x31316, x31315);
  not i31321(x31321, x31320);
  not i31325(x31325, x31324);
  not i31330(x31330, x31329);
  not i31334(x31334, x31333);
  not i31339(x31339, x31338);
  not i31343(x31343, x31342);
  not i31348(x31348, x31347);
  not i31352(x31352, x31351);
  not i31357(x31357, x31356);
  not i31361(x31361, x31360);
  not i31366(x31366, x31365);
  not i31370(x31370, x31369);
  not i31375(x31375, x31374);
  not i31379(x31379, x31378);
  not i31384(x31384, x31383);
  not i31388(x31388, x31387);
  not i31393(x31393, x31392);
  not i31397(x31397, x31396);
  not i31402(x31402, x31401);
  not i31406(x31406, x31405);
  not i31411(x31411, x31410);
  not i31415(x31415, x31414);
  not i31420(x31420, x31419);
  not i31424(x31424, x31423);
  not i31429(x31429, x31428);
  not i31433(x31433, x31432);
  not i31438(x31438, x31437);
  not i31442(x31442, x31441);
  not i31447(x31447, x31446);
  not i31451(x31451, x31450);
  not i31455(x31455, x31454);
  not i31459(x31459, x31458);
  not i31463(x31463, x31462);
  not i31467(x31467, x31466);
  not i31471(x31471, x31470);
  not i31475(x31475, x31474);
  not i31479(x31479, x31478);
  not i31483(x31483, x31482);
  not i31487(x31487, x31486);
  not i31491(x31491, x31490);
  not i31495(x31495, x31494);
  not i31499(x31499, x31498);
  not i31503(x31503, x31502);
  not i31507(x31507, x31506);
  not i31511(x31511, x31510);
  not i31515(x31515, x31514);
  not i31519(x31519, x31518);
  not i31523(x31523, x31522);
  not i31527(x31527, x31526);
  not i31528(x31528, x30059);
  not i31529(x31529, x30067);
  not i31531(x31531, x30075);
  not i31535(x31535, x30094);
  not i31536(x31536, x30086);
  not i31543(x31543, x30111);
  not i31544(x31544, x30102);
  not i31551(x31551, x30128);
  not i31552(x31552, x30119);
  not i31555(x31555, x31554);
  not i31564(x31564, x30148);
  not i31565(x31565, x30139);
  not i31568(x31568, x31567);
  not i31570(x31570, x30157);
  not i31577(x31577, x31576);
  not i31581(x31581, x31580);
  not i31584(x31584, x30174);
  not i31585(x31585, x30165);
  not i31588(x31588, x31587);
  not i31590(x31590, x30183);
  not i31597(x31597, x31596);
  not i31601(x31601, x31600);
  not i31604(x31604, x30200);
  not i31605(x31605, x30191);
  not i31608(x31608, x31607);
  not i31610(x31610, x30209);
  not i31617(x31617, x31616);
  not i31621(x31621, x31620);
  not i31624(x31624, x30229);
  not i31625(x31625, x30220);
  not i31628(x31628, x31627);
  not i31630(x31630, x30238);
  not i31634(x31634, x30247);
  not i31638(x31638, x31637);
  not i31642(x31642, x31641);
  not i31645(x31645, x30264);
  not i31646(x31646, x30255);
  not i31649(x31649, x31648);
  not i31651(x31651, x30273);
  not i31655(x31655, x30282);
  not i31659(x31659, x31658);
  not i31663(x31663, x31662);
  not i31666(x31666, x30299);
  not i31667(x31667, x30290);
  not i31670(x31670, x31669);
  not i31672(x31672, x30308);
  not i31677(x31677, x30317);
  not i31683(x31683, x31682);
  not i31687(x31687, x31686);
  not i31690(x31690, x30337);
  not i31691(x31691, x30328);
  not i31694(x31694, x31693);
  not i31696(x31696, x30346);
  not i31701(x31701, x30363);
  not i31702(x31702, x30355);
  not i31708(x31708, x31707);
  not i31712(x31712, x31711);
  not i31718(x31718, x30380);
  not i31719(x31719, x30371);
  not i31722(x31722, x31721);
  not i31724(x31724, x30389);
  not i31729(x31729, x30407);
  not i31730(x31730, x30398);
  not i31736(x31736, x31735);
  not i31740(x31740, x31739);
  not i31746(x31746, x30424);
  not i31747(x31747, x30415);
  not i31750(x31750, x31749);
  not i31752(x31752, x30433);
  not i31757(x31757, x30451);
  not i31758(x31758, x30442);
  not i31761(x31761, x31760);
  not i31765(x31765, x31764);
  not i31770(x31770, x31769);
  not i31774(x31774, x31773);
  not i31780(x31780, x30471);
  not i31781(x31781, x30462);
  not i31784(x31784, x31783);
  not i31786(x31786, x30480);
  not i31791(x31791, x30498);
  not i31792(x31792, x30489);
  not i31795(x31795, x31794);
  not i31797(x31797, x30507);
  not i31800(x31800, x31799);
  not i31805(x31805, x31804);
  not i31809(x31809, x31808);
  not i31814(x31814, x31813);
  not i31820(x31820, x30524);
  not i31821(x31821, x30515);
  not i31824(x31824, x31823);
  not i31826(x31826, x30533);
  not i31831(x31831, x30551);
  not i31832(x31832, x30542);
  not i31835(x31835, x31834);
  not i31837(x31837, x30560);
  not i31840(x31840, x31839);
  not i31845(x31845, x31844);
  not i31849(x31849, x31848);
  not i31854(x31854, x31853);
  not i31860(x31860, x30577);
  not i31861(x31861, x30568);
  not i31864(x31864, x31863);
  not i31866(x31866, x30586);
  not i31871(x31871, x30604);
  not i31872(x31872, x30595);
  not i31875(x31875, x31874);
  not i31877(x31877, x30613);
  not i31880(x31880, x31879);
  not i31885(x31885, x31884);
  not i31889(x31889, x31888);
  not i31894(x31894, x31893);
  not i31900(x31900, x30633);
  not i31901(x31901, x30624);
  not i31904(x31904, x31903);
  not i31906(x31906, x30642);
  not i31911(x31911, x30660);
  not i31912(x31912, x30651);
  not i31915(x31915, x31914);
  not i31917(x31917, x30669);
  not i31920(x31920, x31919);
  not i31922(x31922, x30678);
  not i31926(x31926, x31925);
  not i31930(x31930, x31929);
  not i31935(x31935, x31934);
  not i31939(x31939, x31938);
  not i31942(x31942, x30695);
  not i31943(x31943, x30686);
  not i31946(x31946, x31945);
  not i31948(x31948, x30704);
  not i31953(x31953, x30722);
  not i31954(x31954, x30713);
  not i31957(x31957, x31956);
  not i31959(x31959, x30731);
  not i31962(x31962, x31961);
  not i31964(x31964, x30740);
  not i31968(x31968, x31967);
  not i31972(x31972, x31971);
  not i31977(x31977, x31976);
  not i31981(x31981, x31980);
  not i31984(x31984, x30757);
  not i31985(x31985, x30748);
  not i31988(x31988, x31987);
  not i31990(x31990, x30766);
  not i31995(x31995, x30784);
  not i31996(x31996, x30775);
  not i31999(x31999, x31998);
  not i32001(x32001, x30793);
  not i32004(x32004, x32003);
  not i32007(x32007, x30802);
  not i32013(x32013, x32012);
  not i32017(x32017, x32016);
  not i32022(x32022, x32021);
  not i32026(x32026, x32025);
  not i32029(x32029, x30822);
  not i32030(x32030, x30813);
  not i32033(x32033, x32032);
  not i32035(x32035, x30831);
  not i32040(x32040, x30849);
  not i32041(x32041, x30840);
  not i32044(x32044, x32043);
  not i32046(x32046, x30858);
  not i32049(x32049, x32048);
  not i32052(x32052, x30875);
  not i32053(x32053, x30867);
  not i32059(x32059, x32058);
  not i32063(x32063, x32062);
  not i32068(x32068, x32067);
  not i32072(x32072, x32071);
  not i32078(x32078, x30892);
  not i32079(x32079, x30883);
  not i32082(x32082, x32081);
  not i32084(x32084, x30901);
  not i32087(x32087, x32086);
  not i32090(x32090, x30919);
  not i32091(x32091, x30910);
  not i32094(x32094, x32093);
  not i32096(x32096, x30928);
  not i32099(x32099, x32098);
  not i32102(x32102, x30946);
  not i32103(x32103, x30937);
  not i32109(x32109, x32108);
  not i32113(x32113, x32112);
  not i32118(x32118, x32117);
  not i32122(x32122, x32121);
  not i32128(x32128, x30963);
  not i32129(x32129, x30954);
  not i32132(x32132, x32131);
  not i32134(x32134, x30972);
  not i32137(x32137, x32136);
  not i32140(x32140, x30990);
  not i32141(x32141, x30981);
  not i32144(x32144, x32143);
  not i32146(x32146, x30999);
  not i32149(x32149, x32148);
  not i32152(x32152, x31017);
  not i32153(x32153, x31008);
  not i32156(x32156, x32155);
  not i32160(x32160, x32159);
  not i32165(x32165, x32164);
  not i32169(x32169, x32168);
  not i32174(x32174, x32173);
  not i32178(x32178, x32177);
  not i32184(x32184, x31037);
  not i32185(x32185, x31028);
  not i32188(x32188, x32187);
  not i32190(x32190, x31046);
  not i32193(x32193, x32192);
  not i32196(x32196, x31064);
  not i32197(x32197, x31055);
  not i32200(x32200, x32199);
  not i32202(x32202, x31073);
  not i32205(x32205, x32204);
  not i32208(x32208, x31091);
  not i32209(x32209, x31082);
  not i32212(x32212, x32211);
  not i32214(x32214, x31100);
  not i32217(x32217, x32216);
  not i32222(x32222, x32221);
  not i32226(x32226, x32225);
  not i32231(x32231, x32230);
  not i32235(x32235, x32234);
  not i32240(x32240, x32239);
  not i32244(x32244, x32243);
  not i32247(x32247, x31117);
  not i32248(x32248, x31108);
  not i32251(x32251, x32250);
  not i32253(x32253, x31126);
  not i32256(x32256, x32255);
  not i32259(x32259, x31144);
  not i32260(x32260, x31135);
  not i32263(x32263, x32262);
  not i32265(x32265, x31153);
  not i32268(x32268, x32267);
  not i32271(x32271, x31171);
  not i32272(x32272, x31162);
  not i32275(x32275, x32274);
  not i32277(x32277, x31180);
  not i32280(x32280, x32279);
  not i32285(x32285, x32284);
  not i32289(x32289, x32288);
  not i32294(x32294, x32293);
  not i32298(x32298, x32297);
  not i32303(x32303, x32302);
  not i32307(x32307, x32306);
  not i32310(x32310, x31197);
  not i32311(x32311, x31188);
  not i32314(x32314, x32313);
  not i32316(x32316, x31206);
  not i32319(x32319, x32318);
  not i32322(x32322, x31224);
  not i32323(x32323, x31215);
  not i32326(x32326, x32325);
  not i32328(x32328, x31233);
  not i32331(x32331, x32330);
  not i32334(x32334, x31251);
  not i32335(x32335, x31242);
  not i32338(x32338, x32337);
  not i32340(x32340, x31260);
  not i32343(x32343, x32342);
  not i32348(x32348, x32347);
  not i32352(x32352, x32351);
  not i32356(x32356, x32355);
  not i32361(x32361, x32360);
  not i32365(x32365, x32364);
  not i32370(x32370, x32369);
  not i32374(x32374, x32373);
  not i32377(x32377, x31281);
  not i32378(x32378, x31272);
  not i32381(x32381, x32380);
  not i32383(x32383, x31290);
  not i32386(x32386, x32385);
  not i32389(x32389, x31308);
  not i32390(x32390, x31299);
  not i32393(x32393, x32392);
  not i32395(x32395, x31317);
  not i32398(x32398, x32397);
  not i32401(x32401, x31335);
  not i32402(x32402, x31326);
  not i32405(x32405, x32404);
  not i32407(x32407, x31344);
  not i32410(x32410, x32409);
  not i32412(x32412, x31353);
  not i32416(x32416, x32415);
  not i32420(x32420, x32419);
  not i32424(x32424, x32423);
  not i32429(x32429, x32428);
  not i32433(x32433, x32432);
  not i32438(x32438, x32437);
  not i32442(x32442, x32441);
  not i32445(x32445, x31371);
  not i32446(x32446, x31362);
  not i32449(x32449, x32448);
  not i32451(x32451, x31380);
  not i32454(x32454, x32453);
  not i32456(x32456, x31398);
  not i32457(x32457, x31389);
  not i32460(x32460, x32459);
  not i32462(x32462, x31407);
  not i32465(x32465, x32464);
  not i32467(x32467, x31425);
  not i32468(x32468, x31416);
  not i32471(x32471, x32470);
  not i32473(x32473, x31434);
  not i32476(x32476, x32475);
  not i32477(x32477, x31443);
  not i32481(x32481, x32480);
  not i32485(x32485, x32484);
  not i32489(x32489, x32488);
  not i32493(x32493, x32492);
  not i32497(x32497, x32496);
  not i32501(x32501, x32500);
  not i32505(x32505, x32504);
  not i32509(x32509, x32508);
  not i32513(x32513, x32512);
  not i32517(x32517, x32516);
  not i32521(x32521, x32520);
  not i32525(x32525, x32524);
  not i32529(x32529, x32528);
  not i32530(x32530, x31559);
  not i32534(x32534, x32533);
  not i32535(x32535, x31573);
  not i32536(x32536, x31582);
  not i32540(x32540, x32539);
  not i32541(x32541, x31593);
  not i32542(x32542, x31602);
  not i32546(x32546, x32545);
  not i32550(x32550, x32549);
  not i32551(x32551, x31613);
  not i32552(x32552, x31622);
  not i32556(x32556, x32555);
  not i32560(x32560, x32559);
  not i32561(x32561, x31633);
  not i32562(x32562, x31643);
  not i32566(x32566, x32565);
  not i32570(x32570, x32569);
  not i32571(x32571, x31654);
  not i32572(x32572, x31664);
  not i32576(x32576, x32575);
  not i32580(x32580, x32579);
  not i32582(x32582, x31675);
  not i32585(x32585, x31688);
  not i32589(x32589, x32588);
  not i32593(x32593, x32592);
  not i32595(x32595, x31699);
  not i32598(x32598, x31713);
  not i32602(x32602, x32601);
  not i32606(x32606, x32605);
  not i32610(x32610, x32609);
  not i32612(x32612, x31727);
  not i32615(x32615, x31741);
  not i32619(x32619, x32618);
  not i32623(x32623, x32622);
  not i32627(x32627, x32626);
  not i32629(x32629, x31766);
  not i32630(x32630, x31755);
  not i32633(x32633, x31775);
  not i32637(x32637, x32636);
  not i32641(x32641, x32640);
  not i32645(x32645, x32644);
  not i32647(x32647, x31801);
  not i32648(x32648, x31789);
  not i32651(x32651, x31810);
  not i32653(x32653, x31818);
  not i32656(x32656, x32655);
  not i32660(x32660, x32659);
  not i32664(x32664, x32663);
  not i32666(x32666, x31841);
  not i32667(x32667, x31829);
  not i32670(x32670, x31850);
  not i32672(x32672, x31858);
  not i32675(x32675, x32674);
  not i32679(x32679, x32678);
  not i32683(x32683, x32682);
  not i32687(x32687, x32686);
  not i32690(x32690, x31881);
  not i32691(x32691, x31869);
  not i32694(x32694, x31890);
  not i32696(x32696, x31898);
  not i32699(x32699, x32698);
  not i32703(x32703, x32702);
  not i32707(x32707, x32706);
  not i32711(x32711, x32710);
  not i32717(x32717, x31921);
  not i32718(x32718, x31909);
  not i32721(x32721, x31931);
  not i32723(x32723, x31940);
  not i32726(x32726, x32725);
  not i32730(x32730, x32729);
  not i32734(x32734, x32733);
  not i32738(x32738, x32737);
  not i32744(x32744, x31963);
  not i32745(x32745, x31951);
  not i32748(x32748, x31973);
  not i32750(x32750, x31982);
  not i32753(x32753, x32752);
  not i32757(x32757, x32756);
  not i32761(x32761, x32760);
  not i32765(x32765, x32764);
  not i32771(x32771, x32005);
  not i32772(x32772, x31993);
  not i32775(x32775, x32774);
  not i32779(x32779, x32778);
  not i32781(x32781, x32018);
  not i32783(x32783, x32027);
  not i32786(x32786, x32785);
  not i32790(x32790, x32789);
  not i32794(x32794, x32793);
  not i32798(x32798, x32797);
  not i32804(x32804, x32050);
  not i32805(x32805, x32038);
  not i32808(x32808, x32807);
  not i32812(x32812, x32811);
  not i32814(x32814, x32064);
  not i32816(x32816, x32073);
  not i32819(x32819, x32818);
  not i32823(x32823, x32822);
  not i32827(x32827, x32826);
  not i32832(x32832, x32831);
  not i32836(x32836, x32835);
  not i32842(x32842, x32100);
  not i32843(x32843, x32088);
  not i32846(x32846, x32845);
  not i32850(x32850, x32849);
  not i32852(x32852, x32114);
  not i32854(x32854, x32123);
  not i32857(x32857, x32856);
  not i32861(x32861, x32860);
  not i32865(x32865, x32864);
  not i32870(x32870, x32869);
  not i32874(x32874, x32873);
  not i32880(x32880, x32150);
  not i32881(x32881, x32138);
  not i32884(x32884, x32883);
  not i32886(x32886, x32161);
  not i32889(x32889, x32888);
  not i32891(x32891, x32170);
  not i32893(x32893, x32179);
  not i32896(x32896, x32895);
  not i32900(x32900, x32899);
  not i32904(x32904, x32903);
  not i32909(x32909, x32908);
  not i32913(x32913, x32912);
  not i32919(x32919, x32206);
  not i32920(x32920, x32194);
  not i32923(x32923, x32922);
  not i32925(x32925, x32218);
  not i32928(x32928, x32927);
  not i32930(x32930, x32227);
  not i32932(x32932, x32236);
  not i32935(x32935, x32934);
  not i32937(x32937, x32245);
  not i32940(x32940, x32939);
  not i32944(x32944, x32943);
  not i32949(x32949, x32948);
  not i32953(x32953, x32952);
  not i32959(x32959, x32269);
  not i32960(x32960, x32257);
  not i32963(x32963, x32962);
  not i32965(x32965, x32281);
  not i32968(x32968, x32967);
  not i32970(x32970, x32290);
  not i32972(x32972, x32299);
  not i32975(x32975, x32974);
  not i32977(x32977, x32308);
  not i32980(x32980, x32979);
  not i32984(x32984, x32983);
  not i32989(x32989, x32988);
  not i32993(x32993, x32992);
  not i32999(x32999, x32332);
  not i33000(x33000, x32320);
  not i33003(x33003, x33002);
  not i33005(x33005, x32344);
  not i33008(x33008, x33007);
  not i33011(x33011, x32357);
  not i33014(x33014, x33013);
  not i33016(x33016, x32366);
  not i33019(x33019, x33018);
  not i33022(x33022, x32375);
  not i33025(x33025, x33024);
  not i33029(x33029, x33028);
  not i33034(x33034, x33033);
  not i33038(x33038, x33037);
  not i33043(x33043, x33042);
  not i33047(x33047, x33046);
  not i33050(x33050, x32399);
  not i33051(x33051, x32387);
  not i33054(x33054, x33053);
  not i33056(x33056, x32411);
  not i33059(x33059, x33058);
  not i33061(x33061, x32425);
  not i33064(x33064, x33063);
  not i33066(x33066, x32434);
  not i33069(x33069, x33068);
  not i33071(x33071, x32443);
  not i33074(x33074, x33073);
  not i33078(x33078, x33077);
  not i33082(x33082, x33081);
  not i33086(x33086, x33085);
  not i33090(x33090, x33089);
  not i33094(x33094, x33093);
  not i33104(x33104, x33103);
  not i33108(x33108, x33107);
  not i33115(x33115, x33114);
  not i33122(x33122, x33121);
  not i33126(x33126, x33125);
  not i33134(x33134, x33133);
  not i33138(x33138, x33137);
  not i33146(x33146, x33145);
  not i33150(x33150, x33149);
  not i33158(x33158, x33157);
  not i33162(x33162, x33161);
  not i33170(x33170, x33169);
  not i33174(x33174, x33173);
  not i33179(x33179, x33178);
  not i33183(x33183, x33182);
  not i33187(x33187, x33186);
  not i33192(x33192, x33191);
  not i33196(x33196, x33195);
  not i33200(x33200, x33199);
  not i33205(x33205, x33204);
  not i33209(x33209, x33208);
  not i33213(x33213, x33212);
  not i33218(x33218, x33217);
  not i33222(x33222, x33221);
  not i33226(x33226, x33225);
  not i33231(x33231, x33230);
  not i33235(x33235, x33234);
  not i33239(x33239, x33238);
  not i33243(x33243, x33242);
  not i33248(x33248, x33247);
  not i33252(x33252, x33251);
  not i33257(x33257, x33256);
  not i33261(x33261, x33260);
  not i33265(x33265, x33264);
  not i33270(x33270, x33269);
  not i33274(x33274, x33273);
  not i33279(x33279, x33278);
  not i33283(x33283, x33282);
  not i33287(x33287, x33286);
  not i33292(x33292, x33291);
  not i33296(x33296, x33295);
  not i33301(x33301, x33300);
  not i33305(x33305, x33304);
  not i33309(x33309, x33308);
  not i33314(x33314, x33313);
  not i33318(x33318, x33317);
  not i33323(x33323, x33322);
  not i33327(x33327, x33326);
  not i33331(x33331, x33330);
  not i33336(x33336, x33335);
  not i33340(x33340, x33339);
  not i33342(x33342, x32688);
  not i33346(x33346, x33345);
  not i33350(x33350, x33349);
  not i33354(x33354, x33353);
  not i33359(x33359, x33358);
  not i33363(x33363, x33362);
  not i33366(x33366, x32712);
  not i33369(x33369, x33368);
  not i33373(x33373, x33372);
  not i33378(x33378, x33377);
  not i33382(x33382, x33381);
  not i33387(x33387, x33386);
  not i33391(x33391, x33390);
  not i33394(x33394, x32739);
  not i33397(x33397, x33396);
  not i33401(x33401, x33400);
  not i33406(x33406, x33405);
  not i33410(x33410, x33409);
  not i33415(x33415, x33414);
  not i33419(x33419, x33418);
  not i33422(x33422, x32766);
  not i33425(x33425, x33424);
  not i33429(x33429, x33428);
  not i33434(x33434, x33433);
  not i33438(x33438, x33437);
  not i33441(x33441, x32780);
  not i33444(x33444, x33443);
  not i33448(x33448, x33447);
  not i33451(x33451, x32799);
  not i33454(x33454, x33453);
  not i33458(x33458, x33457);
  not i33463(x33463, x33462);
  not i33467(x33467, x33466);
  not i33470(x33470, x32813);
  not i33473(x33473, x33472);
  not i33475(x33475, x32828);
  not i33478(x33478, x33477);
  not i33481(x33481, x32837);
  not i33484(x33484, x33483);
  not i33488(x33488, x33487);
  not i33493(x33493, x33492);
  not i33497(x33497, x33496);
  not i33500(x33500, x32851);
  not i33503(x33503, x33502);
  not i33505(x33505, x32866);
  not i33508(x33508, x33507);
  not i33511(x33511, x32875);
  not i33514(x33514, x33513);
  not i33518(x33518, x33517);
  not i33523(x33523, x33522);
  not i33527(x33527, x33526);
  not i33530(x33530, x32890);
  not i33533(x33533, x33532);
  not i33535(x33535, x32905);
  not i33538(x33538, x33537);
  not i33541(x33541, x32914);
  not i33544(x33544, x33543);
  not i33548(x33548, x33547);
  not i33553(x33553, x33552);
  not i33557(x33557, x33556);
  not i33560(x33560, x32929);
  not i33563(x33563, x33562);
  not i33565(x33565, x32945);
  not i33568(x33568, x33567);
  not i33571(x33571, x32954);
  not i33574(x33574, x33573);
  not i33578(x33578, x33577);
  not i33583(x33583, x33582);
  not i33587(x33587, x33586);
  not i33590(x33590, x32969);
  not i33593(x33593, x33592);
  not i33595(x33595, x32985);
  not i33598(x33598, x33597);
  not i33601(x33601, x32994);
  not i33604(x33604, x33603);
  not i33608(x33608, x33607);
  not i33613(x33613, x33612);
  not i33617(x33617, x33616);
  not i33620(x33620, x33020);
  not i33621(x33621, x33009);
  not i33624(x33624, x33623);
  not i33626(x33626, x33030);
  not i33629(x33629, x33628);
  not i33631(x33631, x33048);
  not i33632(x33632, x33039);
  not i33635(x33635, x33634);
  not i33639(x33639, x33638);
  not i33643(x33643, x33642);
  not i33647(x33647, x33646);
  not i33660(x33660, x33659);
  not i33665(x33665, x33127);
  not i33668(x33668, x33667);
  not i33673(x33673, x33139);
  not i33676(x33676, x33675);
  not i33681(x33681, x33151);
  not i33684(x33684, x33683);
  not i33689(x33689, x33163);
  not i33692(x33692, x33691);
  not i33697(x33697, x33175);
  not i33700(x33700, x33699);
  not i33704(x33704, x33703);
  not i33708(x33708, x33707);
  not i33711(x33711, x33188);
  not i33714(x33714, x33713);
  not i33718(x33718, x33717);
  not i33722(x33722, x33721);
  not i33725(x33725, x33201);
  not i33728(x33728, x33727);
  not i33732(x33732, x33731);
  not i33736(x33736, x33735);
  not i33739(x33739, x33214);
  not i33742(x33742, x33741);
  not i33746(x33746, x33745);
  not i33750(x33750, x33749);
  not i33753(x33753, x33227);
  not i33756(x33756, x33755);
  not i33760(x33760, x33759);
  not i33764(x33764, x33763);
  not i33769(x33769, x33768);
  not i33771(x33771, x33244);
  not i33774(x33774, x33773);
  not i33779(x33779, x33778);
  not i33783(x33783, x33782);
  not i33786(x33786, x33253);
  not i33789(x33789, x33788);
  not i33791(x33791, x33266);
  not i33794(x33794, x33793);
  not i33799(x33799, x33798);
  not i33803(x33803, x33802);
  not i33806(x33806, x33275);
  not i33809(x33809, x33808);
  not i33811(x33811, x33288);
  not i33814(x33814, x33813);
  not i33819(x33819, x33818);
  not i33823(x33823, x33822);
  not i33826(x33826, x33297);
  not i33829(x33829, x33828);
  not i33831(x33831, x33310);
  not i33834(x33834, x33833);
  not i33839(x33839, x33838);
  not i33843(x33843, x33842);
  not i33846(x33846, x33319);
  not i33849(x33849, x33848);
  not i33851(x33851, x33332);
  not i33854(x33854, x33853);
  not i33859(x33859, x33858);
  not i33863(x33863, x33862);
  not i33866(x33866, x33341);
  not i33869(x33869, x33868);
  not i33871(x33871, x33355);
  not i33874(x33874, x33873);
  not i33879(x33879, x33878);
  not i33883(x33883, x33882);
  not i33886(x33886, x33374);
  not i33887(x33887, x33364);
  not i33890(x33890, x33889);
  not i33892(x33892, x33383);
  not i33895(x33895, x33894);
  not i33900(x33900, x33899);
  not i33904(x33904, x33903);
  not i33907(x33907, x33402);
  not i33908(x33908, x33392);
  not i33911(x33911, x33910);
  not i33913(x33913, x33411);
  not i33916(x33916, x33915);
  not i33921(x33921, x33920);
  not i33925(x33925, x33924);
  not i33928(x33928, x33430);
  not i33929(x33929, x33420);
  not i33932(x33932, x33931);
  not i33934(x33934, x33439);
  not i33937(x33937, x33936);
  not i33942(x33942, x33941);
  not i33946(x33946, x33945);
  not i33949(x33949, x33459);
  not i33950(x33950, x33449);
  not i33953(x33953, x33952);
  not i33955(x33955, x33468);
  not i33958(x33958, x33957);
  not i33963(x33963, x33962);
  not i33967(x33967, x33966);
  not i33970(x33970, x33489);
  not i33971(x33971, x33479);
  not i33974(x33974, x33973);
  not i33976(x33976, x33498);
  not i33979(x33979, x33978);
  not i33984(x33984, x33983);
  not i33988(x33988, x33987);
  not i33991(x33991, x33519);
  not i33992(x33992, x33509);
  not i33995(x33995, x33994);
  not i33997(x33997, x33528);
  not i34000(x34000, x33999);
  not i34005(x34005, x34004);
  not i34009(x34009, x34008);
  not i34012(x34012, x33549);
  not i34013(x34013, x33539);
  not i34016(x34016, x34015);
  not i34018(x34018, x33558);
  not i34021(x34021, x34020);
  not i34026(x34026, x34025);
  not i34030(x34030, x34029);
  not i34033(x34033, x33579);
  not i34034(x34034, x33569);
  not i34037(x34037, x34036);
  not i34039(x34039, x33588);
  not i34042(x34042, x34041);
  not i34047(x34047, x34046);
  not i34051(x34051, x34050);
  not i34054(x34054, x33609);
  not i34055(x34055, x33599);
  not i34058(x34058, x34057);
  not i34060(x34060, x33618);
  not i34063(x34063, x34062);
  not i34067(x34067, x34066);
  not i34071(x34071, x34070);
  not i34078(x34078, x34077);
  not i34082(x34082, x34081);
  not i34086(x34086, x34085);
  not i34090(x34090, x34089);
  not i34095(x34095, x34094);
  not i34099(x34099, x34098);
  not i34104(x34104, x34103);
  not i34108(x34108, x34107);
  not i34113(x34113, x34112);
  not i34117(x34117, x34116);
  not i34122(x34122, x34121);
  not i34126(x34126, x34125);
  not i34131(x34131, x34130);
  not i34132(x34132, x34128);
  not i34134(x34134, x33709);
  not i34137(x34137, x34136);
  not i34141(x34141, x34140);
  not i34146(x34146, x34145);
  not i34147(x34147, x34143);
  not i34149(x34149, x33723);
  not i34152(x34152, x34151);
  not i34156(x34156, x34155);
  not i34161(x34161, x34160);
  not i34162(x34162, x34158);
  not i34164(x34164, x33737);
  not i34167(x34167, x34166);
  not i34171(x34171, x34170);
  not i34176(x34176, x34175);
  not i34177(x34177, x34173);
  not i34179(x34179, x33751);
  not i34182(x34182, x34181);
  not i34186(x34186, x34185);
  not i34191(x34191, x34190);
  not i34192(x34192, x34188);
  not i34194(x34194, x33765);
  not i34197(x34197, x34196);
  not i34201(x34201, x34200);
  not i34206(x34206, x34205);
  not i34207(x34207, x34203);
  not i34209(x34209, x33784);
  not i34210(x34210, x33775);
  not i34213(x34213, x34212);
  not i34217(x34217, x34216);
  not i34222(x34222, x34221);
  not i34223(x34223, x34219);
  not i34225(x34225, x33804);
  not i34226(x34226, x33795);
  not i34229(x34229, x34228);
  not i34233(x34233, x34232);
  not i34238(x34238, x34237);
  not i34239(x34239, x34235);
  not i34241(x34241, x33824);
  not i34242(x34242, x33815);
  not i34245(x34245, x34244);
  not i34249(x34249, x34248);
  not i34254(x34254, x34253);
  not i34255(x34255, x34251);
  not i34257(x34257, x33844);
  not i34258(x34258, x33835);
  not i34261(x34261, x34260);
  not i34265(x34265, x34264);
  not i34270(x34270, x34269);
  not i34271(x34271, x34267);
  not i34273(x34273, x33864);
  not i34274(x34274, x33855);
  not i34277(x34277, x34276);
  not i34281(x34281, x34280);
  not i34286(x34286, x34285);
  not i34287(x34287, x34283);
  not i34289(x34289, x33884);
  not i34290(x34290, x33875);
  not i34293(x34293, x34292);
  not i34297(x34297, x34296);
  not i34302(x34302, x34301);
  not i34303(x34303, x34299);
  not i34305(x34305, x33905);
  not i34306(x34306, x33896);
  not i34309(x34309, x34308);
  not i34313(x34313, x34312);
  not i34318(x34318, x34317);
  not i34319(x34319, x34315);
  not i34321(x34321, x33926);
  not i34322(x34322, x33917);
  not i34325(x34325, x34324);
  not i34329(x34329, x34328);
  not i34334(x34334, x34333);
  not i34335(x34335, x34331);
  not i34337(x34337, x33947);
  not i34338(x34338, x33938);
  not i34341(x34341, x34340);
  not i34345(x34345, x34344);
  not i34350(x34350, x34349);
  not i34351(x34351, x34347);
  not i34353(x34353, x33968);
  not i34354(x34354, x33959);
  not i34357(x34357, x34356);
  not i34361(x34361, x34360);
  not i34366(x34366, x34365);
  not i34367(x34367, x34363);
  not i34369(x34369, x33989);
  not i34370(x34370, x33980);
  not i34373(x34373, x34372);
  not i34377(x34377, x34376);
  not i34382(x34382, x34381);
  not i34383(x34383, x34379);
  not i34385(x34385, x34010);
  not i34386(x34386, x34001);
  not i34389(x34389, x34388);
  not i34393(x34393, x34392);
  not i34398(x34398, x34397);
  not i34399(x34399, x34395);
  not i34401(x34401, x34031);
  not i34402(x34402, x34022);
  not i34405(x34405, x34404);
  not i34409(x34409, x34408);
  not i34414(x34414, x34413);
  not i34415(x34415, x34411);
  not i34417(x34417, x34052);
  not i34418(x34418, x34043);
  not i34421(x34421, x34420);
  not i34425(x34425, x34424);
  not i34429(x34429, x34428);
  not i34439(x34439, x34438);
  not i34443(x34443, x34442);
  not i34444(x34444, x34091);
  not i34448(x34448, x34447);
  not i34449(x34449, x34100);
  not i34453(x34453, x34452);
  not i34454(x34454, x34109);
  not i34458(x34458, x34457);
  not i34459(x34459, x34118);
  not i34463(x34463, x34462);
  not i34465(x34465, x34127);
  not i34468(x34468, x34467);
  not i34472(x34472, x34471);
  not i34475(x34475, x34142);
  not i34478(x34478, x34477);
  not i34482(x34482, x34481);
  not i34485(x34485, x34157);
  not i34488(x34488, x34487);
  not i34492(x34492, x34491);
  not i34495(x34495, x34172);
  not i34498(x34498, x34497);
  not i34502(x34502, x34501);
  not i34505(x34505, x34187);
  not i34508(x34508, x34507);
  not i34512(x34512, x34511);
  not i34515(x34515, x34202);
  not i34518(x34518, x34517);
  not i34522(x34522, x34521);
  not i34525(x34525, x34218);
  not i34528(x34528, x34527);
  not i34532(x34532, x34531);
  not i34535(x34535, x34234);
  not i34538(x34538, x34537);
  not i34542(x34542, x34541);
  not i34545(x34545, x34250);
  not i34548(x34548, x34547);
  not i34552(x34552, x34551);
  not i34555(x34555, x34266);
  not i34558(x34558, x34557);
  not i34562(x34562, x34561);
  not i34565(x34565, x34282);
  not i34568(x34568, x34567);
  not i34572(x34572, x34571);
  not i34575(x34575, x34298);
  not i34578(x34578, x34577);
  not i34582(x34582, x34581);
  not i34585(x34585, x34314);
  not i34588(x34588, x34587);
  not i34592(x34592, x34591);
  not i34595(x34595, x34330);
  not i34598(x34598, x34597);
  not i34602(x34602, x34601);
  not i34605(x34605, x34346);
  not i34608(x34608, x34607);
  not i34612(x34612, x34611);
  not i34615(x34615, x34362);
  not i34618(x34618, x34617);
  not i34622(x34622, x34621);
  not i34625(x34625, x34378);
  not i34628(x34628, x34627);
  not i34632(x34632, x34631);
  not i34635(x34635, x34394);
  not i34638(x34638, x34637);
  not i34642(x34642, x34641);
  not i34645(x34645, x34410);
  not i34648(x34648, x34647);
  not i34652(x34652, x34651);
  not i34656(x34656, x34655);
  not i34664(x34664, x34663);
  not i34668(x34668, x34667);
  not i34672(x34672, x34671);
  not i34676(x34676, x34675);
  not i34681(x34681, x34680);
  not i34685(x34685, x34684);
  not i34690(x34690, x34689);
  not i34694(x34694, x34693);
  not i34699(x34699, x34698);
  not i34703(x34703, x34702);
  not i34708(x34708, x34707);
  not i34712(x34712, x34711);
  not i34717(x34717, x34716);
  not i34721(x34721, x34720);
  not i34726(x34726, x34725);
  not i34730(x34730, x34729);
  not i34733(x34733, x34473);
  not i34736(x34736, x34735);
  not i34740(x34740, x34739);
  not i34743(x34743, x34483);
  not i34746(x34746, x34745);
  not i34750(x34750, x34749);
  not i34753(x34753, x34493);
  not i34756(x34756, x34755);
  not i34760(x34760, x34759);
  not i34763(x34763, x34503);
  not i34766(x34766, x34765);
  not i34770(x34770, x34769);
  not i34773(x34773, x34513);
  not i34776(x34776, x34775);
  not i34780(x34780, x34779);
  not i34783(x34783, x34523);
  not i34786(x34786, x34785);
  not i34790(x34790, x34789);
  not i34793(x34793, x34533);
  not i34796(x34796, x34795);
  not i34800(x34800, x34799);
  not i34803(x34803, x34543);
  not i34806(x34806, x34805);
  not i34810(x34810, x34809);
  not i34813(x34813, x34553);
  not i34816(x34816, x34815);
  not i34820(x34820, x34819);
  not i34823(x34823, x34563);
  not i34826(x34826, x34825);
  not i34830(x34830, x34829);
  not i34833(x34833, x34573);
  not i34836(x34836, x34835);
  not i34840(x34840, x34839);
  not i34843(x34843, x34583);
  not i34846(x34846, x34845);
  not i34850(x34850, x34849);
  not i34853(x34853, x34593);
  not i34856(x34856, x34855);
  not i34860(x34860, x34859);
  not i34863(x34863, x34603);
  not i34866(x34866, x34865);
  not i34870(x34870, x34869);
  not i34873(x34873, x34613);
  not i34876(x34876, x34875);
  not i34880(x34880, x34879);
  not i34883(x34883, x34623);
  not i34886(x34886, x34885);
  not i34890(x34890, x34889);
  not i34893(x34893, x34633);
  not i34896(x34896, x34895);
  not i34900(x34900, x34899);
  not i34903(x34903, x34643);
  not i34906(x34906, x34905);
  not i34910(x34910, x34909);
  not i34912(x34912, x34660);
  not i34918(x34918, x34917);
  not i34922(x34922, x34921);
  not i34924(x34924, x34677);
  not i34927(x34927, x34926);
  not i34929(x34929, x34686);
  not i34932(x34932, x34931);
  not i34934(x34934, x34695);
  not i34937(x34937, x34936);
  not i34939(x34939, x34704);
  not i34942(x34942, x34941);
  not i34944(x34944, x34713);
  not i34947(x34947, x34946);
  not i34949(x34949, x34722);
  not i34952(x34952, x34951);
  not i34954(x34954, x34731);
  not i34957(x34957, x34956);
  not i34959(x34959, x34741);
  not i34962(x34962, x34961);
  not i34964(x34964, x34751);
  not i34967(x34967, x34966);
  not i34969(x34969, x34761);
  not i34972(x34972, x34971);
  not i34974(x34974, x34771);
  not i34977(x34977, x34976);
  not i34979(x34979, x34781);
  not i34982(x34982, x34981);
  not i34984(x34984, x34791);
  not i34987(x34987, x34986);
  not i34989(x34989, x34801);
  not i34992(x34992, x34991);
  not i34994(x34994, x34811);
  not i34997(x34997, x34996);
  not i34999(x34999, x34821);
  not i35002(x35002, x35001);
  not i35004(x35004, x34831);
  not i35007(x35007, x35006);
  not i35009(x35009, x34841);
  not i35012(x35012, x35011);
  not i35014(x35014, x34851);
  not i35017(x35017, x35016);
  not i35019(x35019, x34861);
  not i35022(x35022, x35021);
  not i35024(x35024, x34871);
  not i35027(x35027, x35026);
  not i35029(x35029, x34881);
  not i35032(x35032, x35031);
  not i35034(x35034, x34891);
  not i35037(x35037, x35036);
  not i35039(x35039, x34901);
  not i35042(x35042, x35041);
  not i35043(x35043, x34911);
  not i35044(x35044, x34915);
  not i35045(x35045, x34919);
  not i35046(x35046, x34923);
  not i35047(x35047, x34928);
  not i35048(x35048, x34933);
  not i35049(x35049, x34938);
  not i35050(x35050, x34943);
  not i35051(x35051, x34948);
  not i35052(x35052, x34953);
  not i35053(x35053, x34958);
  not i35054(x35054, x34963);
  not i35055(x35055, x34968);
  not i35056(x35056, x34973);
  not i35057(x35057, x34978);
  not i35058(x35058, x34983);
  not i35059(x35059, x34988);
  not i35060(x35060, x34993);
  not i35061(x35061, x34998);
  not i35062(x35062, x35003);
  not i35063(x35063, x35008);
  not i35064(x35064, x35013);
  not i35065(x35065, x35018);
  not i35066(x35066, x35023);
  not i35067(x35067, x35028);
  not i35073(x35073, x35072);
  not i35077(x35077, x35076);
  not i35081(x35081, x35080);
  not i35085(x35085, x35084);
  not i35089(x35089, x35088);
  not i35093(x35093, x35092);
  not i35097(x35097, x35096);
  not i35101(x35101, x35100);
  not i35105(x35105, x35104);
  not i35109(x35109, x35108);
  not i35113(x35113, x35112);
  not i35117(x35117, x35116);
  not i35121(x35121, x35120);
  not i35125(x35125, x35124);
  not i35129(x35129, x35128);
  not i35133(x35133, x35132);
  not i35137(x35137, x35136);
  not i35141(x35141, x35140);
  not i35145(x35145, x35144);
  not i35149(x35149, x35148);
  not i35153(x35153, x35152);
  not i35157(x35157, x35156);
  not i35161(x35161, x35160);
  not i35165(x35165, x35164);
  not i35166(x35166, x35069);
  not i35168(x35168, x35071);
  not i35171(x35171, x35075);
  not i35174(x35174, x35079);
  not i35177(x35177, x35176);
  not i35179(x35179, x35083);
  not i35182(x35182, x35181);
  not i35184(x35184, x35087);
  not i35187(x35187, x35186);
  not i35189(x35189, x35091);
  not i35192(x35192, x35191);
  not i35194(x35194, x35095);
  not i35197(x35197, x35196);
  not i35199(x35199, x35099);
  not i35202(x35202, x35201);
  not i35204(x35204, x35103);
  not i35207(x35207, x35206);
  not i35209(x35209, x35107);
  not i35212(x35212, x35211);
  not i35214(x35214, x35111);
  not i35217(x35217, x35216);
  not i35219(x35219, x35115);
  not i35222(x35222, x35221);
  not i35224(x35224, x35119);
  not i35227(x35227, x35226);
  not i35229(x35229, x35123);
  not i35232(x35232, x35231);
  not i35234(x35234, x35127);
  not i35237(x35237, x35236);
  not i35239(x35239, x35131);
  not i35242(x35242, x35241);
  not i35244(x35244, x35135);
  not i35247(x35247, x35246);
  not i35249(x35249, x35139);
  not i35252(x35252, x35251);
  not i35254(x35254, x35143);
  not i35257(x35257, x35256);
  not i35259(x35259, x35147);
  not i35262(x35262, x35261);
  not i35264(x35264, x35151);
  not i35267(x35267, x35266);
  not i35269(x35269, x35155);
  not i35272(x35272, x35271);
  not i35274(x35274, x35159);
  not i35277(x35277, x35276);
  not i35279(x35279, x35163);
  not i35282(x35282, x35281);
  not i35283(x35283, x35169);
  not i35284(x35284, x35172);
  not i35286(x35286, x35175);
  not i35289(x35289, x35180);
  not i35292(x35292, x35185);
  not i35295(x35295, x35190);
  not i35298(x35298, x35195);
  not i35301(x35301, x35300);
  not i35303(x35303, x35200);
  not i35306(x35306, x35305);
  not i35308(x35308, x35205);
  not i35311(x35311, x35310);
  not i35313(x35313, x35210);
  not i35316(x35316, x35315);
  not i35318(x35318, x35215);
  not i35321(x35321, x35320);
  not i35323(x35323, x35220);
  not i35326(x35326, x35325);
  not i35328(x35328, x35225);
  not i35331(x35331, x35330);
  not i35333(x35333, x35230);
  not i35336(x35336, x35335);
  not i35338(x35338, x35235);
  not i35341(x35341, x35340);
  not i35343(x35343, x35240);
  not i35346(x35346, x35345);
  not i35348(x35348, x35245);
  not i35351(x35351, x35350);
  not i35353(x35353, x35250);
  not i35356(x35356, x35355);
  not i35358(x35358, x35255);
  not i35361(x35361, x35360);
  not i35363(x35363, x35260);
  not i35366(x35366, x35365);
  not i35368(x35368, x35265);
  not i35371(x35371, x35370);
  not i35373(x35373, x35270);
  not i35376(x35376, x35375);
  not i35378(x35378, x35275);
  not i35381(x35381, x35380);
  not i35383(x35383, x35280);
  not i35386(x35386, x35385);
  not i35387(x35387, x35287);
  not i35388(x35388, x35290);
  not i35389(x35389, x35293);
  not i35390(x35390, x35296);
  not i35392(x35392, x35299);
  not i35395(x35395, x35304);
  not i35398(x35398, x35309);
  not i35401(x35401, x35314);
  not i35404(x35404, x35319);
  not i35407(x35407, x35324);
  not i35410(x35410, x35329);
  not i35413(x35413, x35334);
  not i35416(x35416, x35339);
  not i35419(x35419, x35418);
  not i35421(x35421, x35344);
  not i35424(x35424, x35423);
  not i35426(x35426, x35349);
  not i35429(x35429, x35428);
  not i35431(x35431, x35354);
  not i35434(x35434, x35433);
  not i35436(x35436, x35359);
  not i35439(x35439, x35438);
  not i35441(x35441, x35364);
  not i35444(x35444, x35443);
  not i35446(x35446, x35369);
  not i35449(x35449, x35448);
  not i35451(x35451, x35374);
  not i35454(x35454, x35453);
  not i35456(x35456, x35379);
  not i35459(x35459, x35458);
  not i35461(x35461, x35384);
  not i35464(x35464, x35463);
  not i35465(x35465, x35399);
  not i35466(x35466, x35402);
  not i35467(x35467, x35405);
  not i35468(x35468, x35408);
  not i35469(x35469, x35411);
  not i35470(x35470, x35414);
  not i35472(x35472, x35417);
  not i35475(x35475, x35422);
  not i35478(x35478, x35427);
  not i35481(x35481, x35432);
  not i35484(x35484, x35437);
  not i35487(x35487, x35442);
  not i35490(x35490, x35447);
  not i35493(x35493, x35452);
  not i35496(x35496, x35457);
  not i35499(x35499, x35462);
  not i35503(x35503, x35502);
  not i35507(x35507, x35506);
  not i35511(x35511, x35510);
  not i35515(x35515, x35514);
  not i35519(x35519, x35518);
  not i35523(x35523, x35522);
  not i35527(x35527, x35526);
  not i35531(x35531, x35530);
  not i35533(x35533, x35393);
  not i35536(x35536, x35535);
  not i35538(x35538, x35396);
  not i35541(x35541, x35540);
  not i35545(x35545, x35544);
  not i35549(x35549, x35548);
  not i35553(x35553, x35552);
  not i35557(x35557, x35556);
  not i35561(x35561, x35560);
  not i35565(x35565, x35564);
  not i35567(x35567, x35473);
  not i35570(x35570, x35569);
  not i35572(x35572, x35476);
  not i35575(x35575, x35574);
  not i35577(x35577, x35479);
  not i35580(x35580, x35579);
  not i35582(x35582, x35482);
  not i35585(x35585, x35584);
  not i35587(x35587, x35485);
  not i35590(x35590, x35589);
  not i35592(x35592, x35488);
  not i35595(x35595, x35594);
  not i35597(x35597, x35491);
  not i35600(x35600, x35599);
  not i35602(x35602, x35494);
  not i35605(x35605, x35604);
  not i35607(x35607, x35497);
  not i35610(x35610, x35609);
  not i35612(x35612, x35500);
  not i35615(x35615, x35614);
  not i35617(x35617, x35616);
  not i35619(x35619, x35618);
  not i35621(x35621, x35620);
  not i35623(x35623, x35622);
  not i35625(x35625, x35624);
  not i35627(x35627, x35626);
  not i35629(x35629, x35628);
  not i35631(x35631, x35630);
  not i35633(x35633, x35632);
  not i35635(x35635, x35634);
  not i35637(x35637, x35636);
  not i35639(x35639, x35638);
  not i35641(x35641, x35640);
  not i35643(x35643, x35642);
  not i35645(x35645, x35644);
  not i35647(x35647, x35646);
  not i35649(x35649, x35648);
  not i35651(x35651, x35650);
  not i35653(x35653, x35652);
  not i35655(x35655, x35654);
  not i35657(x35657, x35656);
  not i35659(x35659, x35658);
  not i35661(x35661, x35660);
  not i35663(x35663, x35662);
  not i35665(x35665, x35664);
  not i35667(x35667, x35666);
  not i35669(x35669, x35668);
  not i35671(x35671, x35670);
  not i35673(x35673, x35672);
  not i35675(x35675, x35674);
  not i35678(x35678, x35677);
  not i35680(x35680, x35679);
  not i35682(x35682, x35681);
  not i35684(x35684, x35683);
  not i35686(x35686, x35685);
  not i35688(x35688, x35687);
  not i35690(x35690, x35689);
  not i35692(x35692, x35691);
  not i35694(x35694, x35693);
  not i35696(x35696, x35695);
  not i35698(x35698, x35697);
  not i35700(x35700, x35699);
  not i35702(x35702, x35701);
  not i35704(x35704, x35703);
  not i35706(x35706, x35705);
  not i35708(x35708, x35707);
  not i35710(x35710, x35709);
  not i35712(x35712, x35711);
  not i35714(x35714, x35713);
  not i35716(x35716, x35715);
  not i35718(x35718, x35717);
  not i35720(x35720, x35719);
  not i35722(x35722, x35721);
  not i35724(x35724, x35723);
  not i35726(x35726, x35725);
  not i35728(x35728, x35727);
  not i35730(x35730, x35729);
  not i35732(x35732, x35731);
  not i35737(x35737, x35736);
  not i35739(x35739, x35738);
  not i35741(x35741, x35740);
  not i35743(x35743, x35742);
  not i35745(x35745, x35744);
  not i35747(x35747, x35746);
  not i35749(x35749, x35748);
  not i35751(x35751, x35750);
  not i35753(x35753, x35752);
  not i35755(x35755, x35754);
  not i35757(x35757, x35756);
  not i35759(x35759, x35758);
  not i35761(x35761, x35760);
  not i35763(x35763, x35762);
  not i35765(x35765, x35764);
  not i35767(x35767, x35766);
  not i35769(x35769, x35768);
  not i35771(x35771, x35770);
  not i35773(x35773, x35772);
  not i35775(x35775, x35774);
  not i35777(x35777, x35776);
  not i35779(x35779, x35778);
  not i35781(x35781, x35780);
  not i35783(x35783, x35782);
  not i35793(x35793, x35792);
  not i35795(x35795, x35794);
  not i35797(x35797, x35796);
  not i35799(x35799, x35798);
  not i35801(x35801, x35800);
  not i35803(x35803, x35802);
  not i35805(x35805, x35804);
  not i35807(x35807, x35806);
  not i35809(x35809, x35808);
  not i35811(x35811, x35810);
  not i35813(x35813, x35812);
  not i35815(x35815, x35814);
  not i35817(x35817, x35816);
  not i35819(x35819, x35818);
  not i35821(x35821, x35820);
  not i35839(x35839, x35838);
  not i35843(x35843, x35842);
  not i35847(x35847, x35846);
  not i35851(x35851, x35850);
  not i35855(x35855, x35854);
  not i35859(x35859, x35858);
  not i35863(x35863, x35862);
  not i35867(x35867, x35866);
  not i35871(x35871, x35870);
  not i35875(x35875, x35874);
  not i35879(x35879, x35878);
  not i35883(x35883, x35882);
  not i35887(x35887, x35886);
  not i35891(x35891, x35890);
  not i35895(x35895, x35894);
  not i35899(x35899, x35898);
  not i35903(x35903, x35902);
  not i35907(x35907, x35906);
  not i35911(x35911, x35910);
  not i35915(x35915, x35914);
  not i35919(x35919, x35918);
  not i35923(x35923, x35922);
  not i35927(x35927, x35926);
  not i35931(x35931, x35930);
  not i35935(x35935, x35934);
  not i35939(x35939, x35938);
  not i35943(x35943, x35942);
  not i35947(x35947, x35946);
  not i35951(x35951, x35950);
  not i35955(x35955, x35954);
  not i35959(x35959, x35958);
  not i35960(x35960, x29004);
  not i35962(x35962, x35961);
  not i35964(x35964, x35963);
  not i35966(x35966, x35965);
  not i35968(x35968, x35967);
  not i35970(x35970, x35969);
  not i35972(x35972, x35971);
  not i35974(x35974, x35973);
  not i35976(x35976, x35975);
  not i35978(x35978, x35977);
  not i35980(x35980, x35979);
  not i35982(x35982, x35981);
  not i35984(x35984, x35983);
  not i35986(x35986, x35985);
  not i35988(x35988, x35987);
  not i35990(x35990, x35989);
  not i35992(x35992, x35991);
  not i36026(x36026, x36025);
  not i36028(x36028, x36027);
  not i36030(x36030, x36029);
  not i36032(x36032, x36031);
  not i36034(x36034, x36033);
  not i36036(x36036, x36035);
  not i36038(x36038, x36037);
  not i36040(x36040, x36039);
  not i36042(x36042, x36041);
  not i36044(x36044, x36043);
  not i36046(x36046, x36045);
  not i36048(x36048, x36047);
  not i36050(x36050, x36049);
  not i36052(x36052, x36051);
  not i36054(x36054, x36053);
  not i36056(x36056, x36055);
  not i36058(x36058, x36057);
  not i36060(x36060, x36059);
  not i36062(x36062, x36061);
  not i36064(x36064, x36063);
  not i36066(x36066, x36065);
  not i36068(x36068, x36067);
  not i36070(x36070, x36069);
  not i36072(x36072, x36071);
  not i36074(x36074, x36073);
  not i36076(x36076, x36075);
  not i36078(x36078, x36077);
  not i36080(x36080, x36079);
  not i36082(x36082, x36081);
  not i36084(x36084, x36083);
  not i36086(x36086, x36085);
  not i36088(x36088, x36087);
  not i38911(x38911, x38848);
  not i38912(x38912, x38850);
  not i38913(x38913, x38852);
  not i38914(x38914, x38854);
  not i38915(x38915, x38856);
  not i38916(x38916, x38858);
  not i38917(x38917, x38860);
  not i38918(x38918, x38862);
  not i38919(x38919, x38864);
  not i38920(x38920, x38866);
  not i38921(x38921, x38868);
  not i38922(x38922, x38870);
  not i38923(x38923, x38872);
  not i38924(x38924, x38874);
  not i38925(x38925, x38876);
  not i38926(x38926, x38878);
  not i38927(x38927, x38880);
  not i38928(x38928, x38882);
  not i38929(x38929, x38884);
  not i38930(x38930, x38886);
  not i38931(x38931, x38888);
  not i38932(x38932, x38890);
  not i38933(x38933, x38892);
  not i38934(x38934, x38894);
  not i38935(x38935, x38896);
  not i38936(x38936, x38898);
  not i38937(x38937, x38900);
  not i38938(x38938, x38902);
  not i38939(x38939, x38904);
  not i38940(x38940, x38906);
  not i38941(x38941, x38908);
  not i38942(x38942, x38910);
  not i39040(x39040, x38945);
  not i39041(x39041, x73027);
  not i39044(x39044, x39043);
  not i39046(x39046, x38948);
  not i39047(x39047, x73032);
  not i39050(x39050, x39049);
  not i39052(x39052, x38951);
  not i39053(x39053, x73037);
  not i39056(x39056, x39055);
  not i39058(x39058, x38954);
  not i39059(x39059, x73042);
  not i39062(x39062, x39061);
  not i39064(x39064, x38957);
  not i39065(x39065, x73047);
  not i39068(x39068, x39067);
  not i39070(x39070, x38960);
  not i39071(x39071, x73052);
  not i39074(x39074, x39073);
  not i39076(x39076, x38963);
  not i39077(x39077, x73057);
  not i39080(x39080, x39079);
  not i39082(x39082, x38966);
  not i39083(x39083, x73062);
  not i39086(x39086, x39085);
  not i39088(x39088, x38969);
  not i39089(x39089, x73067);
  not i39092(x39092, x39091);
  not i39094(x39094, x38972);
  not i39095(x39095, x73072);
  not i39098(x39098, x39097);
  not i39100(x39100, x38975);
  not i39101(x39101, x73077);
  not i39104(x39104, x39103);
  not i39106(x39106, x38978);
  not i39107(x39107, x73082);
  not i39110(x39110, x39109);
  not i39112(x39112, x38981);
  not i39113(x39113, x73087);
  not i39116(x39116, x39115);
  not i39118(x39118, x38984);
  not i39119(x39119, x73092);
  not i39122(x39122, x39121);
  not i39124(x39124, x38987);
  not i39125(x39125, x73097);
  not i39128(x39128, x39127);
  not i39130(x39130, x38990);
  not i39131(x39131, x73102);
  not i39134(x39134, x39133);
  not i39136(x39136, x38993);
  not i39137(x39137, x73107);
  not i39140(x39140, x39139);
  not i39142(x39142, x38996);
  not i39143(x39143, x73112);
  not i39146(x39146, x39145);
  not i39148(x39148, x38999);
  not i39149(x39149, x73117);
  not i39152(x39152, x39151);
  not i39154(x39154, x39002);
  not i39155(x39155, x73122);
  not i39158(x39158, x39157);
  not i39160(x39160, x39005);
  not i39161(x39161, x73127);
  not i39164(x39164, x39163);
  not i39166(x39166, x39008);
  not i39167(x39167, x73132);
  not i39170(x39170, x39169);
  not i39172(x39172, x39011);
  not i39173(x39173, x73137);
  not i39176(x39176, x39175);
  not i39178(x39178, x39014);
  not i39179(x39179, x73142);
  not i39182(x39182, x39181);
  not i39184(x39184, x39017);
  not i39185(x39185, x73147);
  not i39188(x39188, x39187);
  not i39190(x39190, x39020);
  not i39191(x39191, x73152);
  not i39194(x39194, x39193);
  not i39196(x39196, x39023);
  not i39197(x39197, x73157);
  not i39200(x39200, x39199);
  not i39202(x39202, x39026);
  not i39203(x39203, x73162);
  not i39206(x39206, x39205);
  not i39208(x39208, x39029);
  not i39209(x39209, x73167);
  not i39212(x39212, x39211);
  not i39214(x39214, x39032);
  not i39215(x39215, x73172);
  not i39218(x39218, x39217);
  not i39220(x39220, x39035);
  not i39221(x39221, x73177);
  not i39224(x39224, x39223);
  not i39226(x39226, x39038);
  not i39227(x39227, x73182);
  not i39230(x39230, x39229);
  not i39231(x39231, x39039);
  not i39232(x39232, x39045);
  not i39233(x39233, x39051);
  not i39234(x39234, x39057);
  not i39235(x39235, x39063);
  not i39236(x39236, x39069);
  not i39237(x39237, x39075);
  not i39238(x39238, x39081);
  not i39239(x39239, x39087);
  not i39240(x39240, x39093);
  not i39241(x39241, x39099);
  not i39242(x39242, x39105);
  not i39243(x39243, x39111);
  not i39244(x39244, x39117);
  not i39245(x39245, x39123);
  not i39246(x39246, x39129);
  not i39247(x39247, x39135);
  not i39248(x39248, x39141);
  not i39249(x39249, x39147);
  not i39250(x39250, x39153);
  not i39251(x39251, x39159);
  not i39252(x39252, x39165);
  not i39253(x39253, x39171);
  not i39254(x39254, x39177);
  not i39255(x39255, x39183);
  not i39256(x39256, x39189);
  not i39257(x39257, x39195);
  not i39258(x39258, x39201);
  not i39259(x39259, x39207);
  not i39260(x39260, x39213);
  not i39266(x39266, x39265);
  not i39270(x39270, x39269);
  not i39274(x39274, x39273);
  not i39278(x39278, x39277);
  not i39282(x39282, x39281);
  not i39286(x39286, x39285);
  not i39290(x39290, x39289);
  not i39294(x39294, x39293);
  not i39298(x39298, x39297);
  not i39302(x39302, x39301);
  not i39306(x39306, x39305);
  not i39310(x39310, x39309);
  not i39314(x39314, x39313);
  not i39318(x39318, x39317);
  not i39322(x39322, x39321);
  not i39326(x39326, x39325);
  not i39330(x39330, x39329);
  not i39334(x39334, x39333);
  not i39338(x39338, x39337);
  not i39342(x39342, x39341);
  not i39346(x39346, x39345);
  not i39350(x39350, x39349);
  not i39354(x39354, x39353);
  not i39358(x39358, x39357);
  not i39362(x39362, x39361);
  not i39366(x39366, x39365);
  not i39370(x39370, x39369);
  not i39374(x39374, x39373);
  not i39378(x39378, x39377);
  not i39382(x39382, x39381);
  not i39384(x39384, x39264);
  not i39387(x39387, x39268);
  not i39390(x39390, x39272);
  not i39393(x39393, x39392);
  not i39395(x39395, x39276);
  not i39398(x39398, x39397);
  not i39400(x39400, x39280);
  not i39403(x39403, x39402);
  not i39405(x39405, x39284);
  not i39408(x39408, x39407);
  not i39410(x39410, x39288);
  not i39413(x39413, x39412);
  not i39415(x39415, x39292);
  not i39418(x39418, x39417);
  not i39420(x39420, x39296);
  not i39423(x39423, x39422);
  not i39425(x39425, x39300);
  not i39428(x39428, x39427);
  not i39430(x39430, x39304);
  not i39433(x39433, x39432);
  not i39435(x39435, x39308);
  not i39438(x39438, x39437);
  not i39440(x39440, x39312);
  not i39443(x39443, x39442);
  not i39445(x39445, x39316);
  not i39448(x39448, x39447);
  not i39450(x39450, x39320);
  not i39453(x39453, x39452);
  not i39455(x39455, x39324);
  not i39458(x39458, x39457);
  not i39460(x39460, x39328);
  not i39463(x39463, x39462);
  not i39465(x39465, x39332);
  not i39468(x39468, x39467);
  not i39470(x39470, x39336);
  not i39473(x39473, x39472);
  not i39475(x39475, x39340);
  not i39478(x39478, x39477);
  not i39480(x39480, x39344);
  not i39483(x39483, x39482);
  not i39485(x39485, x39348);
  not i39488(x39488, x39487);
  not i39490(x39490, x39352);
  not i39493(x39493, x39492);
  not i39495(x39495, x39356);
  not i39498(x39498, x39497);
  not i39500(x39500, x39360);
  not i39503(x39503, x39502);
  not i39505(x39505, x39364);
  not i39508(x39508, x39507);
  not i39510(x39510, x39368);
  not i39513(x39513, x39512);
  not i39515(x39515, x39372);
  not i39518(x39518, x39517);
  not i39520(x39520, x39376);
  not i39523(x39523, x39522);
  not i39525(x39525, x39380);
  not i39528(x39528, x39527);
  not i39530(x39530, x39391);
  not i39533(x39533, x39396);
  not i39536(x39536, x39401);
  not i39539(x39539, x39406);
  not i39542(x39542, x39411);
  not i39545(x39545, x39544);
  not i39547(x39547, x39416);
  not i39550(x39550, x39549);
  not i39552(x39552, x39421);
  not i39555(x39555, x39554);
  not i39557(x39557, x39426);
  not i39560(x39560, x39559);
  not i39562(x39562, x39431);
  not i39565(x39565, x39564);
  not i39567(x39567, x39436);
  not i39570(x39570, x39569);
  not i39572(x39572, x39441);
  not i39575(x39575, x39574);
  not i39577(x39577, x39446);
  not i39580(x39580, x39579);
  not i39582(x39582, x39451);
  not i39585(x39585, x39584);
  not i39587(x39587, x39456);
  not i39590(x39590, x39589);
  not i39592(x39592, x39461);
  not i39595(x39595, x39594);
  not i39597(x39597, x39466);
  not i39600(x39600, x39599);
  not i39602(x39602, x39471);
  not i39605(x39605, x39604);
  not i39607(x39607, x39476);
  not i39610(x39610, x39609);
  not i39612(x39612, x39481);
  not i39615(x39615, x39614);
  not i39617(x39617, x39486);
  not i39620(x39620, x39619);
  not i39622(x39622, x39491);
  not i39625(x39625, x39624);
  not i39627(x39627, x39496);
  not i39630(x39630, x39629);
  not i39632(x39632, x39501);
  not i39635(x39635, x39634);
  not i39637(x39637, x39506);
  not i39640(x39640, x39639);
  not i39642(x39642, x39511);
  not i39645(x39645, x39644);
  not i39647(x39647, x39516);
  not i39650(x39650, x39649);
  not i39652(x39652, x39521);
  not i39655(x39655, x39654);
  not i39657(x39657, x39526);
  not i39660(x39660, x39659);
  not i39662(x39662, x39543);
  not i39665(x39665, x39548);
  not i39668(x39668, x39553);
  not i39671(x39671, x39558);
  not i39674(x39674, x39563);
  not i39677(x39677, x39568);
  not i39680(x39680, x39573);
  not i39683(x39683, x39578);
  not i39686(x39686, x39583);
  not i39689(x39689, x39688);
  not i39691(x39691, x39588);
  not i39694(x39694, x39693);
  not i39696(x39696, x39593);
  not i39699(x39699, x39698);
  not i39701(x39701, x39598);
  not i39704(x39704, x39703);
  not i39706(x39706, x39603);
  not i39709(x39709, x39708);
  not i39711(x39711, x39608);
  not i39714(x39714, x39713);
  not i39716(x39716, x39613);
  not i39719(x39719, x39718);
  not i39721(x39721, x39618);
  not i39724(x39724, x39723);
  not i39726(x39726, x39623);
  not i39729(x39729, x39728);
  not i39731(x39731, x39628);
  not i39734(x39734, x39733);
  not i39736(x39736, x39633);
  not i39739(x39739, x39738);
  not i39741(x39741, x39638);
  not i39744(x39744, x39743);
  not i39746(x39746, x39643);
  not i39749(x39749, x39748);
  not i39751(x39751, x39648);
  not i39754(x39754, x39753);
  not i39756(x39756, x39653);
  not i39759(x39759, x39758);
  not i39761(x39761, x39658);
  not i39764(x39764, x39763);
  not i39766(x39766, x39687);
  not i39769(x39769, x39692);
  not i39772(x39772, x39697);
  not i39775(x39775, x39702);
  not i39778(x39778, x39707);
  not i39781(x39781, x39712);
  not i39784(x39784, x39717);
  not i39787(x39787, x39722);
  not i39790(x39790, x39727);
  not i39793(x39793, x39732);
  not i39796(x39796, x39737);
  not i39799(x39799, x39742);
  not i39802(x39802, x39747);
  not i39805(x39805, x39752);
  not i39808(x39808, x39757);
  not i39811(x39811, x39762);
  not i39815(x39815, x39814);
  not i39817(x39817, x39262);
  not i39820(x39820, x39819);
  not i39822(x39822, x39385);
  not i39825(x39825, x39824);
  not i39827(x39827, x39388);
  not i39830(x39830, x39829);
  not i39832(x39832, x39531);
  not i39835(x39835, x39834);
  not i39837(x39837, x39534);
  not i39840(x39840, x39839);
  not i39842(x39842, x39537);
  not i39845(x39845, x39844);
  not i39847(x39847, x39540);
  not i39850(x39850, x39849);
  not i39852(x39852, x39663);
  not i39855(x39855, x39854);
  not i39857(x39857, x39666);
  not i39860(x39860, x39859);
  not i39862(x39862, x39669);
  not i39865(x39865, x39864);
  not i39867(x39867, x39672);
  not i39870(x39870, x39869);
  not i39872(x39872, x39675);
  not i39875(x39875, x39874);
  not i39877(x39877, x39678);
  not i39880(x39880, x39879);
  not i39882(x39882, x39681);
  not i39885(x39885, x39884);
  not i39887(x39887, x39684);
  not i39890(x39890, x39889);
  not i39892(x39892, x39767);
  not i39895(x39895, x39894);
  not i39897(x39897, x39770);
  not i39900(x39900, x39899);
  not i39902(x39902, x39773);
  not i39905(x39905, x39904);
  not i39907(x39907, x39776);
  not i39910(x39910, x39909);
  not i39912(x39912, x39779);
  not i39915(x39915, x39914);
  not i39917(x39917, x39782);
  not i39920(x39920, x39919);
  not i39922(x39922, x39785);
  not i39925(x39925, x39924);
  not i39927(x39927, x39788);
  not i39930(x39930, x39929);
  not i39932(x39932, x39791);
  not i39935(x39935, x39934);
  not i39937(x39937, x39794);
  not i39940(x39940, x39939);
  not i39942(x39942, x39797);
  not i39945(x39945, x39944);
  not i39947(x39947, x39800);
  not i39950(x39950, x39949);
  not i39952(x39952, x39803);
  not i39955(x39955, x39954);
  not i39957(x39957, x39806);
  not i39960(x39960, x39959);
  not i39962(x39962, x39809);
  not i39965(x39965, x39964);
  not i39967(x39967, x39812);
  not i39970(x39970, x39969);
  not i39973(x39973, x39972);
  not i39975(x39975, x39974);
  not i39977(x39977, x39976);
  not i39979(x39979, x39978);
  not i39981(x39981, x39980);
  not i39983(x39983, x39982);
  not i39985(x39985, x39984);
  not i39987(x39987, x39986);
  not i39990(x39990, x39989);
  not i39992(x39992, x39991);
  not i39994(x39994, x39993);
  not i39996(x39996, x39995);
  not i39998(x39998, x39997);
  not i40000(x40000, x39999);
  not i40002(x40002, x40001);
  not i40004(x40004, x40003);
  not i40006(x40006, x40005);
  not i40008(x40008, x40007);
  not i40010(x40010, x40009);
  not i40012(x40012, x40011);
  not i40014(x40014, x40013);
  not i40016(x40016, x40015);
  not i40018(x40018, x40017);
  not i40020(x40020, x40019);
  not i40022(x40022, x40021);
  not i40025(x40025, x40024);
  not i40027(x40027, x40026);
  not i40029(x40029, x40028);
  not i40031(x40031, x40030);
  not i40033(x40033, x40032);
  not i40035(x40035, x40034);
  not i40037(x40037, x40036);
  not i40039(x40039, x40038);
  not i40041(x40041, x40040);
  not i40043(x40043, x40042);
  not i40045(x40045, x40044);
  not i40047(x40047, x40046);
  not i40049(x40049, x40048);
  not i40051(x40051, x40050);
  not i40053(x40053, x40052);
  not i40055(x40055, x40054);
  not i40057(x40057, x40056);
  not i40059(x40059, x40058);
  not i40061(x40061, x40060);
  not i40063(x40063, x40062);
  not i40065(x40065, x40064);
  not i40067(x40067, x40066);
  not i40069(x40069, x40068);
  not i40071(x40071, x40070);
  not i40073(x40073, x40072);
  not i40075(x40075, x40074);
  not i40078(x40078, x40077);
  not i40080(x40080, x40079);
  not i40082(x40082, x40081);
  not i40084(x40084, x40083);
  not i40086(x40086, x40085);
  not i40088(x40088, x40087);
  not i40090(x40090, x40089);
  not i40092(x40092, x40091);
  not i40094(x40094, x40093);
  not i40096(x40096, x40095);
  not i40098(x40098, x40097);
  not i40100(x40100, x40099);
  not i40102(x40102, x40101);
  not i40104(x40104, x40103);
  not i40106(x40106, x40105);
  not i40108(x40108, x40107);
  not i40110(x40110, x40109);
  not i40112(x40112, x40111);
  not i40114(x40114, x40113);
  not i40116(x40116, x40115);
  not i40118(x40118, x40117);
  not i40120(x40120, x40119);
  not i40122(x40122, x40121);
  not i40124(x40124, x40123);
  not i40126(x40126, x40125);
  not i40128(x40128, x40127);
  not i40130(x40130, x40129);
  not i40132(x40132, x40131);
  not i40134(x40134, x40133);
  not i40136(x40136, x40135);
  not i40138(x40138, x40137);
  not i40140(x40140, x40139);
  not i40142(x40142, x40141);
  not i40144(x40144, x40143);
  not i40146(x40146, x40145);
  not i40149(x40149, x40148);
  not i40151(x40151, x40150);
  not i40153(x40153, x40152);
  not i40155(x40155, x40154);
  not i40157(x40157, x40156);
  not i40159(x40159, x40158);
  not i40161(x40161, x40160);
  not i40163(x40163, x40162);
  not i40165(x40165, x40164);
  not i40167(x40167, x40166);
  not i40169(x40169, x40168);
  not i40171(x40171, x40170);
  not i40173(x40173, x40172);
  not i40175(x40175, x40174);
  not i40177(x40177, x40176);
  not i40179(x40179, x40178);
  not i40181(x40181, x40180);
  not i40183(x40183, x40182);
  not i40185(x40185, x40184);
  not i40187(x40187, x40186);
  not i40189(x40189, x40188);
  not i40191(x40191, x40190);
  not i40193(x40193, x40192);
  not i40195(x40195, x40194);
  not i40197(x40197, x40196);
  not i40199(x40199, x40198);
  not i40201(x40201, x40200);
  not i40203(x40203, x40202);
  not i40205(x40205, x40204);
  not i40207(x40207, x40206);
  not i40209(x40209, x40208);
  not i40211(x40211, x40210);
  not i40213(x40213, x40212);
  not i40215(x40215, x40214);
  not i40217(x40217, x40216);
  not i40219(x40219, x40218);
  not i40221(x40221, x40220);
  not i40223(x40223, x40222);
  not i40225(x40225, x40224);
  not i40227(x40227, x40226);
  not i40229(x40229, x40228);
  not i40231(x40231, x40230);
  not i40233(x40233, x40232);
  not i40235(x40235, x40234);
  not i40238(x40238, x40237);
  not i40240(x40240, x40239);
  not i40242(x40242, x40241);
  not i40244(x40244, x40243);
  not i40246(x40246, x40245);
  not i40248(x40248, x40247);
  not i40250(x40250, x40249);
  not i40252(x40252, x40251);
  not i40254(x40254, x40253);
  not i40256(x40256, x40255);
  not i40258(x40258, x40257);
  not i40260(x40260, x40259);
  not i40262(x40262, x40261);
  not i40264(x40264, x40263);
  not i40266(x40266, x40265);
  not i40268(x40268, x40267);
  not i40270(x40270, x40269);
  not i40272(x40272, x40271);
  not i40274(x40274, x40273);
  not i40276(x40276, x40275);
  not i40278(x40278, x40277);
  not i40280(x40280, x40279);
  not i40282(x40282, x40281);
  not i40284(x40284, x40283);
  not i40286(x40286, x40285);
  not i40288(x40288, x40287);
  not i40290(x40290, x40289);
  not i40292(x40292, x40291);
  not i40294(x40294, x40293);
  not i40296(x40296, x40295);
  not i40298(x40298, x40297);
  not i40300(x40300, x40299);
  not i40302(x40302, x40301);
  not i40304(x40304, x40303);
  not i40306(x40306, x40305);
  not i40308(x40308, x40307);
  not i40310(x40310, x40309);
  not i40312(x40312, x40311);
  not i40314(x40314, x40313);
  not i40316(x40316, x40315);
  not i40318(x40318, x40317);
  not i40320(x40320, x40319);
  not i40322(x40322, x40321);
  not i40324(x40324, x40323);
  not i40326(x40326, x40325);
  not i40328(x40328, x40327);
  not i40330(x40330, x40329);
  not i40332(x40332, x40331);
  not i40334(x40334, x40333);
  not i40336(x40336, x40335);
  not i40338(x40338, x40337);
  not i40340(x40340, x40339);
  not i40342(x40342, x40341);
  not i40345(x40345, x40344);
  not i40347(x40347, x40346);
  not i40349(x40349, x40348);
  not i40351(x40351, x40350);
  not i40353(x40353, x40352);
  not i40355(x40355, x40354);
  not i40357(x40357, x40356);
  not i40359(x40359, x40358);
  not i40361(x40361, x40360);
  not i40363(x40363, x40362);
  not i40365(x40365, x40364);
  not i40367(x40367, x40366);
  not i40369(x40369, x40368);
  not i40371(x40371, x40370);
  not i40373(x40373, x40372);
  not i40375(x40375, x40374);
  not i40377(x40377, x40376);
  not i40379(x40379, x40378);
  not i40381(x40381, x40380);
  not i40383(x40383, x40382);
  not i40385(x40385, x40384);
  not i40387(x40387, x40386);
  not i40389(x40389, x40388);
  not i40391(x40391, x40390);
  not i40393(x40393, x40392);
  not i40395(x40395, x40394);
  not i40397(x40397, x40396);
  not i40399(x40399, x40398);
  not i40401(x40401, x40400);
  not i40403(x40403, x40402);
  not i40405(x40405, x40404);
  not i40407(x40407, x40406);
  not i40409(x40409, x40408);
  not i40411(x40411, x40410);
  not i40413(x40413, x40412);
  not i40415(x40415, x40414);
  not i40417(x40417, x40416);
  not i40419(x40419, x40418);
  not i40421(x40421, x40420);
  not i40423(x40423, x40422);
  not i40425(x40425, x40424);
  not i40427(x40427, x40426);
  not i40429(x40429, x40428);
  not i40431(x40431, x40430);
  not i40433(x40433, x40432);
  not i40435(x40435, x40434);
  not i40437(x40437, x40436);
  not i40439(x40439, x40438);
  not i40441(x40441, x40440);
  not i40443(x40443, x40442);
  not i40445(x40445, x40444);
  not i40447(x40447, x40446);
  not i40449(x40449, x40448);
  not i40451(x40451, x40450);
  not i40453(x40453, x40452);
  not i40455(x40455, x40454);
  not i40457(x40457, x40456);
  not i40459(x40459, x40458);
  not i40461(x40461, x40460);
  not i40463(x40463, x40462);
  not i40465(x40465, x40464);
  not i40467(x40467, x40466);
  not i40470(x40470, x40469);
  not i40472(x40472, x40471);
  not i40474(x40474, x40473);
  not i40476(x40476, x40475);
  not i40478(x40478, x40477);
  not i40480(x40480, x40479);
  not i40482(x40482, x40481);
  not i40484(x40484, x40483);
  not i40486(x40486, x40485);
  not i40488(x40488, x40487);
  not i40490(x40490, x40489);
  not i40492(x40492, x40491);
  not i40494(x40494, x40493);
  not i40496(x40496, x40495);
  not i40498(x40498, x40497);
  not i40500(x40500, x40499);
  not i40502(x40502, x40501);
  not i40504(x40504, x40503);
  not i40506(x40506, x40505);
  not i40508(x40508, x40507);
  not i40510(x40510, x40509);
  not i40512(x40512, x40511);
  not i40514(x40514, x40513);
  not i40516(x40516, x40515);
  not i40518(x40518, x40517);
  not i40520(x40520, x40519);
  not i40522(x40522, x40521);
  not i40524(x40524, x40523);
  not i40526(x40526, x40525);
  not i40528(x40528, x40527);
  not i40530(x40530, x40529);
  not i40532(x40532, x40531);
  not i40534(x40534, x40533);
  not i40536(x40536, x40535);
  not i40538(x40538, x40537);
  not i40540(x40540, x40539);
  not i40542(x40542, x40541);
  not i40544(x40544, x40543);
  not i40546(x40546, x40545);
  not i40548(x40548, x40547);
  not i40550(x40550, x40549);
  not i40552(x40552, x40551);
  not i40554(x40554, x40553);
  not i40556(x40556, x40555);
  not i40558(x40558, x40557);
  not i40560(x40560, x40559);
  not i40562(x40562, x40561);
  not i40564(x40564, x40563);
  not i40566(x40566, x40565);
  not i40568(x40568, x40567);
  not i40570(x40570, x40569);
  not i40572(x40572, x40571);
  not i40574(x40574, x40573);
  not i40576(x40576, x40575);
  not i40578(x40578, x40577);
  not i40580(x40580, x40579);
  not i40582(x40582, x40581);
  not i40584(x40584, x40583);
  not i40586(x40586, x40585);
  not i40588(x40588, x40587);
  not i40590(x40590, x40589);
  not i40592(x40592, x40591);
  not i40594(x40594, x40593);
  not i40596(x40596, x40595);
  not i40598(x40598, x40597);
  not i40600(x40600, x40599);
  not i40602(x40602, x40601);
  not i40604(x40604, x40603);
  not i40606(x40606, x40605);
  not i40608(x40608, x40607);
  not i40610(x40610, x40609);
  not i40613(x40613, x40612);
  not i40615(x40615, x40614);
  not i40617(x40617, x40616);
  not i40619(x40619, x40618);
  not i40621(x40621, x40620);
  not i40623(x40623, x40622);
  not i40625(x40625, x40624);
  not i40627(x40627, x40626);
  not i40629(x40629, x40628);
  not i40631(x40631, x40630);
  not i40633(x40633, x40632);
  not i40635(x40635, x40634);
  not i40637(x40637, x40636);
  not i40639(x40639, x40638);
  not i40641(x40641, x40640);
  not i40643(x40643, x40642);
  not i40645(x40645, x40644);
  not i40647(x40647, x40646);
  not i40649(x40649, x40648);
  not i40651(x40651, x40650);
  not i40653(x40653, x40652);
  not i40655(x40655, x40654);
  not i40657(x40657, x40656);
  not i40659(x40659, x40658);
  not i40661(x40661, x40660);
  not i40663(x40663, x40662);
  not i40665(x40665, x40664);
  not i40667(x40667, x40666);
  not i40669(x40669, x40668);
  not i40671(x40671, x40670);
  not i40673(x40673, x40672);
  not i40675(x40675, x40674);
  not i40677(x40677, x40676);
  not i40679(x40679, x40678);
  not i40681(x40681, x40680);
  not i40683(x40683, x40682);
  not i40685(x40685, x40684);
  not i40687(x40687, x40686);
  not i40689(x40689, x40688);
  not i40691(x40691, x40690);
  not i40693(x40693, x40692);
  not i40695(x40695, x40694);
  not i40697(x40697, x40696);
  not i40699(x40699, x40698);
  not i40701(x40701, x40700);
  not i40703(x40703, x40702);
  not i40705(x40705, x40704);
  not i40707(x40707, x40706);
  not i40709(x40709, x40708);
  not i40711(x40711, x40710);
  not i40713(x40713, x40712);
  not i40715(x40715, x40714);
  not i40717(x40717, x40716);
  not i40719(x40719, x40718);
  not i40721(x40721, x40720);
  not i40723(x40723, x40722);
  not i40725(x40725, x40724);
  not i40727(x40727, x40726);
  not i40729(x40729, x40728);
  not i40731(x40731, x40730);
  not i40733(x40733, x40732);
  not i40735(x40735, x40734);
  not i40737(x40737, x40736);
  not i40739(x40739, x40738);
  not i40741(x40741, x40740);
  not i40743(x40743, x40742);
  not i40745(x40745, x40744);
  not i40747(x40747, x40746);
  not i40749(x40749, x40748);
  not i40751(x40751, x40750);
  not i40753(x40753, x40752);
  not i40755(x40755, x40754);
  not i40757(x40757, x40756);
  not i40759(x40759, x40758);
  not i40761(x40761, x40760);
  not i40763(x40763, x40762);
  not i40765(x40765, x40764);
  not i40767(x40767, x40766);
  not i40769(x40769, x40768);
  not i40771(x40771, x40770);
  not i40774(x40774, x40773);
  not i40776(x40776, x40775);
  not i40778(x40778, x40777);
  not i40780(x40780, x40779);
  not i40782(x40782, x40781);
  not i40784(x40784, x40783);
  not i40786(x40786, x40785);
  not i40788(x40788, x40787);
  not i40790(x40790, x40789);
  not i40792(x40792, x40791);
  not i40794(x40794, x40793);
  not i40796(x40796, x40795);
  not i40798(x40798, x40797);
  not i40800(x40800, x40799);
  not i40802(x40802, x40801);
  not i40804(x40804, x40803);
  not i40806(x40806, x40805);
  not i40808(x40808, x40807);
  not i40810(x40810, x40809);
  not i40812(x40812, x40811);
  not i40814(x40814, x40813);
  not i40816(x40816, x40815);
  not i40818(x40818, x40817);
  not i40820(x40820, x40819);
  not i40822(x40822, x40821);
  not i40824(x40824, x40823);
  not i40826(x40826, x40825);
  not i40828(x40828, x40827);
  not i40830(x40830, x40829);
  not i40832(x40832, x40831);
  not i40834(x40834, x40833);
  not i40836(x40836, x40835);
  not i40838(x40838, x40837);
  not i40840(x40840, x40839);
  not i40842(x40842, x40841);
  not i40844(x40844, x40843);
  not i40846(x40846, x40845);
  not i40848(x40848, x40847);
  not i40850(x40850, x40849);
  not i40852(x40852, x40851);
  not i40854(x40854, x40853);
  not i40856(x40856, x40855);
  not i40858(x40858, x40857);
  not i40860(x40860, x40859);
  not i40862(x40862, x40861);
  not i40864(x40864, x40863);
  not i40866(x40866, x40865);
  not i40868(x40868, x40867);
  not i40870(x40870, x40869);
  not i40872(x40872, x40871);
  not i40874(x40874, x40873);
  not i40876(x40876, x40875);
  not i40878(x40878, x40877);
  not i40880(x40880, x40879);
  not i40882(x40882, x40881);
  not i40884(x40884, x40883);
  not i40886(x40886, x40885);
  not i40888(x40888, x40887);
  not i40890(x40890, x40889);
  not i40892(x40892, x40891);
  not i40894(x40894, x40893);
  not i40896(x40896, x40895);
  not i40898(x40898, x40897);
  not i40900(x40900, x40899);
  not i40902(x40902, x40901);
  not i40904(x40904, x40903);
  not i40906(x40906, x40905);
  not i40908(x40908, x40907);
  not i40910(x40910, x40909);
  not i40912(x40912, x40911);
  not i40914(x40914, x40913);
  not i40916(x40916, x40915);
  not i40918(x40918, x40917);
  not i40920(x40920, x40919);
  not i40922(x40922, x40921);
  not i40924(x40924, x40923);
  not i40926(x40926, x40925);
  not i40928(x40928, x40927);
  not i40930(x40930, x40929);
  not i40932(x40932, x40931);
  not i40934(x40934, x40933);
  not i40936(x40936, x40935);
  not i40938(x40938, x40937);
  not i40940(x40940, x40939);
  not i40942(x40942, x40941);
  not i40944(x40944, x40943);
  not i40946(x40946, x40945);
  not i40948(x40948, x40947);
  not i40950(x40950, x40949);
  not i40953(x40953, x40952);
  not i40955(x40955, x40954);
  not i40957(x40957, x40956);
  not i40959(x40959, x40958);
  not i40961(x40961, x40960);
  not i40963(x40963, x40962);
  not i40965(x40965, x40964);
  not i40967(x40967, x40966);
  not i40969(x40969, x40968);
  not i40971(x40971, x40970);
  not i40973(x40973, x40972);
  not i40975(x40975, x40974);
  not i40977(x40977, x40976);
  not i40979(x40979, x40978);
  not i40981(x40981, x40980);
  not i40983(x40983, x40982);
  not i40985(x40985, x40984);
  not i40987(x40987, x40986);
  not i40989(x40989, x40988);
  not i40991(x40991, x40990);
  not i40993(x40993, x40992);
  not i40995(x40995, x40994);
  not i40997(x40997, x40996);
  not i40999(x40999, x40998);
  not i41001(x41001, x41000);
  not i41003(x41003, x41002);
  not i41005(x41005, x41004);
  not i41007(x41007, x41006);
  not i41009(x41009, x41008);
  not i41011(x41011, x41010);
  not i41013(x41013, x41012);
  not i41015(x41015, x41014);
  not i41022(x41022, x41021);
  not i41030(x41030, x41029);
  not i41038(x41038, x41037);
  not i41049(x41049, x41048);
  not i41057(x41057, x41056);
  not i41065(x41065, x41064);
  not i41073(x41073, x41072);
  not i41077(x41077, x41076);
  not i41082(x41082, x41081);
  not i41090(x41090, x41089);
  not i41094(x41094, x41093);
  not i41102(x41102, x41101);
  not i41110(x41110, x41109);
  not i41114(x41114, x41113);
  not i41119(x41119, x41118);
  not i41123(x41123, x41122);
  not i41128(x41128, x41127);
  not i41136(x41136, x41135);
  not i41140(x41140, x41139);
  not i41145(x41145, x41144);
  not i41149(x41149, x41148);
  not i41154(x41154, x41153);
  not i41162(x41162, x41161);
  not i41166(x41166, x41165);
  not i41171(x41171, x41170);
  not i41175(x41175, x41174);
  not i41183(x41183, x41182);
  not i41191(x41191, x41190);
  not i41195(x41195, x41194);
  not i41200(x41200, x41199);
  not i41204(x41204, x41203);
  not i41209(x41209, x41208);
  not i41213(x41213, x41212);
  not i41218(x41218, x41217);
  not i41226(x41226, x41225);
  not i41230(x41230, x41229);
  not i41235(x41235, x41234);
  not i41239(x41239, x41238);
  not i41244(x41244, x41243);
  not i41248(x41248, x41247);
  not i41253(x41253, x41252);
  not i41261(x41261, x41260);
  not i41265(x41265, x41264);
  not i41270(x41270, x41269);
  not i41274(x41274, x41273);
  not i41279(x41279, x41278);
  not i41283(x41283, x41282);
  not i41291(x41291, x41290);
  not i41299(x41299, x41298);
  not i41303(x41303, x41302);
  not i41308(x41308, x41307);
  not i41312(x41312, x41311);
  not i41317(x41317, x41316);
  not i41321(x41321, x41320);
  not i41326(x41326, x41325);
  not i41334(x41334, x41333);
  not i41342(x41342, x41341);
  not i41346(x41346, x41345);
  not i41351(x41351, x41350);
  not i41355(x41355, x41354);
  not i41360(x41360, x41359);
  not i41364(x41364, x41363);
  not i41369(x41369, x41368);
  not i41373(x41373, x41372);
  not i41378(x41378, x41377);
  not i41386(x41386, x41385);
  not i41390(x41390, x41389);
  not i41395(x41395, x41394);
  not i41399(x41399, x41398);
  not i41404(x41404, x41403);
  not i41408(x41408, x41407);
  not i41413(x41413, x41412);
  not i41417(x41417, x41416);
  not i41425(x41425, x41424);
  not i41433(x41433, x41432);
  not i41437(x41437, x41436);
  not i41442(x41442, x41441);
  not i41446(x41446, x41445);
  not i41451(x41451, x41450);
  not i41455(x41455, x41454);
  not i41460(x41460, x41459);
  not i41464(x41464, x41463);
  not i41469(x41469, x41468);
  not i41473(x41473, x41472);
  not i41478(x41478, x41477);
  not i41486(x41486, x41485);
  not i41490(x41490, x41489);
  not i41495(x41495, x41494);
  not i41499(x41499, x41498);
  not i41504(x41504, x41503);
  not i41508(x41508, x41507);
  not i41513(x41513, x41512);
  not i41517(x41517, x41516);
  not i41522(x41522, x41521);
  not i41526(x41526, x41525);
  not i41531(x41531, x41530);
  not i41539(x41539, x41538);
  not i41543(x41543, x41542);
  not i41548(x41548, x41547);
  not i41552(x41552, x41551);
  not i41557(x41557, x41556);
  not i41561(x41561, x41560);
  not i41566(x41566, x41565);
  not i41570(x41570, x41569);
  not i41575(x41575, x41574);
  not i41579(x41579, x41578);
  not i41587(x41587, x41586);
  not i41595(x41595, x41594);
  not i41599(x41599, x41598);
  not i41604(x41604, x41603);
  not i41608(x41608, x41607);
  not i41613(x41613, x41612);
  not i41617(x41617, x41616);
  not i41622(x41622, x41621);
  not i41626(x41626, x41625);
  not i41631(x41631, x41630);
  not i41635(x41635, x41634);
  not i41640(x41640, x41639);
  not i41644(x41644, x41643);
  not i41649(x41649, x41648);
  not i41657(x41657, x41656);
  not i41661(x41661, x41660);
  not i41666(x41666, x41665);
  not i41670(x41670, x41669);
  not i41675(x41675, x41674);
  not i41679(x41679, x41678);
  not i41684(x41684, x41683);
  not i41688(x41688, x41687);
  not i41693(x41693, x41692);
  not i41697(x41697, x41696);
  not i41702(x41702, x41701);
  not i41706(x41706, x41705);
  not i41711(x41711, x41710);
  not i41719(x41719, x41718);
  not i41723(x41723, x41722);
  not i41728(x41728, x41727);
  not i41732(x41732, x41731);
  not i41737(x41737, x41736);
  not i41741(x41741, x41740);
  not i41746(x41746, x41745);
  not i41750(x41750, x41749);
  not i41755(x41755, x41754);
  not i41759(x41759, x41758);
  not i41764(x41764, x41763);
  not i41768(x41768, x41767);
  not i41776(x41776, x41775);
  not i41784(x41784, x41783);
  not i41788(x41788, x41787);
  not i41793(x41793, x41792);
  not i41797(x41797, x41796);
  not i41802(x41802, x41801);
  not i41806(x41806, x41805);
  not i41811(x41811, x41810);
  not i41815(x41815, x41814);
  not i41820(x41820, x41819);
  not i41824(x41824, x41823);
  not i41829(x41829, x41828);
  not i41833(x41833, x41832);
  not i41838(x41838, x41837);
  not i41846(x41846, x41845);
  not i41854(x41854, x41853);
  not i41858(x41858, x41857);
  not i41863(x41863, x41862);
  not i41867(x41867, x41866);
  not i41872(x41872, x41871);
  not i41876(x41876, x41875);
  not i41881(x41881, x41880);
  not i41885(x41885, x41884);
  not i41890(x41890, x41889);
  not i41894(x41894, x41893);
  not i41899(x41899, x41898);
  not i41903(x41903, x41902);
  not i41908(x41908, x41907);
  not i41912(x41912, x41911);
  not i41917(x41917, x41916);
  not i41925(x41925, x41924);
  not i41929(x41929, x41928);
  not i41934(x41934, x41933);
  not i41938(x41938, x41937);
  not i41943(x41943, x41942);
  not i41947(x41947, x41946);
  not i41952(x41952, x41951);
  not i41956(x41956, x41955);
  not i41961(x41961, x41960);
  not i41965(x41965, x41964);
  not i41970(x41970, x41969);
  not i41974(x41974, x41973);
  not i41979(x41979, x41978);
  not i41983(x41983, x41982);
  not i41991(x41991, x41990);
  not i41999(x41999, x41998);
  not i42003(x42003, x42002);
  not i42008(x42008, x42007);
  not i42012(x42012, x42011);
  not i42017(x42017, x42016);
  not i42021(x42021, x42020);
  not i42026(x42026, x42025);
  not i42030(x42030, x42029);
  not i42035(x42035, x42034);
  not i42039(x42039, x42038);
  not i42044(x42044, x42043);
  not i42048(x42048, x42047);
  not i42053(x42053, x42052);
  not i42057(x42057, x42056);
  not i42062(x42062, x42061);
  not i42066(x42066, x42065);
  not i42071(x42071, x42070);
  not i42079(x42079, x42078);
  not i42083(x42083, x42082);
  not i42088(x42088, x42087);
  not i42092(x42092, x42091);
  not i42097(x42097, x42096);
  not i42101(x42101, x42100);
  not i42106(x42106, x42105);
  not i42110(x42110, x42109);
  not i42115(x42115, x42114);
  not i42119(x42119, x42118);
  not i42124(x42124, x42123);
  not i42128(x42128, x42127);
  not i42133(x42133, x42132);
  not i42137(x42137, x42136);
  not i42142(x42142, x42141);
  not i42146(x42146, x42145);
  not i42151(x42151, x42150);
  not i42159(x42159, x42158);
  not i42163(x42163, x42162);
  not i42168(x42168, x42167);
  not i42172(x42172, x42171);
  not i42177(x42177, x42176);
  not i42181(x42181, x42180);
  not i42186(x42186, x42185);
  not i42190(x42190, x42189);
  not i42195(x42195, x42194);
  not i42199(x42199, x42198);
  not i42204(x42204, x42203);
  not i42208(x42208, x42207);
  not i42213(x42213, x42212);
  not i42217(x42217, x42216);
  not i42222(x42222, x42221);
  not i42226(x42226, x42225);
  not i42234(x42234, x42233);
  not i42238(x42238, x42237);
  not i42243(x42243, x42242);
  not i42247(x42247, x42246);
  not i42252(x42252, x42251);
  not i42256(x42256, x42255);
  not i42261(x42261, x42260);
  not i42265(x42265, x42264);
  not i42270(x42270, x42269);
  not i42274(x42274, x42273);
  not i42279(x42279, x42278);
  not i42283(x42283, x42282);
  not i42288(x42288, x42287);
  not i42292(x42292, x42291);
  not i42297(x42297, x42296);
  not i42301(x42301, x42300);
  not i42306(x42306, x42305);
  not i42310(x42310, x42309);
  not i42315(x42315, x42314);
  not i42319(x42319, x42318);
  not i42324(x42324, x42323);
  not i42328(x42328, x42327);
  not i42333(x42333, x42332);
  not i42337(x42337, x42336);
  not i42342(x42342, x42341);
  not i42346(x42346, x42345);
  not i42351(x42351, x42350);
  not i42355(x42355, x42354);
  not i42360(x42360, x42359);
  not i42364(x42364, x42363);
  not i42369(x42369, x42368);
  not i42373(x42373, x42372);
  not i42378(x42378, x42377);
  not i42382(x42382, x42381);
  not i42387(x42387, x42386);
  not i42391(x42391, x42390);
  not i42396(x42396, x42395);
  not i42400(x42400, x42399);
  not i42405(x42405, x42404);
  not i42409(x42409, x42408);
  not i42414(x42414, x42413);
  not i42418(x42418, x42417);
  not i42422(x42422, x42421);
  not i42426(x42426, x42425);
  not i42430(x42430, x42429);
  not i42434(x42434, x42433);
  not i42438(x42438, x42437);
  not i42442(x42442, x42441);
  not i42446(x42446, x42445);
  not i42450(x42450, x42449);
  not i42454(x42454, x42453);
  not i42458(x42458, x42457);
  not i42462(x42462, x42461);
  not i42466(x42466, x42465);
  not i42470(x42470, x42469);
  not i42474(x42474, x42473);
  not i42478(x42478, x42477);
  not i42482(x42482, x42481);
  not i42486(x42486, x42485);
  not i42490(x42490, x42489);
  not i42494(x42494, x42493);
  not i42495(x42495, x41026);
  not i42496(x42496, x41034);
  not i42498(x42498, x41042);
  not i42502(x42502, x41061);
  not i42503(x42503, x41053);
  not i42510(x42510, x41078);
  not i42511(x42511, x41069);
  not i42518(x42518, x41095);
  not i42519(x42519, x41086);
  not i42522(x42522, x42521);
  not i42531(x42531, x41115);
  not i42532(x42532, x41106);
  not i42535(x42535, x42534);
  not i42537(x42537, x41124);
  not i42544(x42544, x42543);
  not i42548(x42548, x42547);
  not i42551(x42551, x41141);
  not i42552(x42552, x41132);
  not i42555(x42555, x42554);
  not i42557(x42557, x41150);
  not i42564(x42564, x42563);
  not i42568(x42568, x42567);
  not i42571(x42571, x41167);
  not i42572(x42572, x41158);
  not i42575(x42575, x42574);
  not i42577(x42577, x41176);
  not i42584(x42584, x42583);
  not i42588(x42588, x42587);
  not i42591(x42591, x41196);
  not i42592(x42592, x41187);
  not i42595(x42595, x42594);
  not i42597(x42597, x41205);
  not i42601(x42601, x41214);
  not i42605(x42605, x42604);
  not i42609(x42609, x42608);
  not i42612(x42612, x41231);
  not i42613(x42613, x41222);
  not i42616(x42616, x42615);
  not i42618(x42618, x41240);
  not i42622(x42622, x41249);
  not i42626(x42626, x42625);
  not i42630(x42630, x42629);
  not i42633(x42633, x41266);
  not i42634(x42634, x41257);
  not i42637(x42637, x42636);
  not i42639(x42639, x41275);
  not i42644(x42644, x41284);
  not i42650(x42650, x42649);
  not i42654(x42654, x42653);
  not i42657(x42657, x41304);
  not i42658(x42658, x41295);
  not i42661(x42661, x42660);
  not i42663(x42663, x41313);
  not i42668(x42668, x41330);
  not i42669(x42669, x41322);
  not i42675(x42675, x42674);
  not i42679(x42679, x42678);
  not i42685(x42685, x41347);
  not i42686(x42686, x41338);
  not i42689(x42689, x42688);
  not i42691(x42691, x41356);
  not i42696(x42696, x41374);
  not i42697(x42697, x41365);
  not i42703(x42703, x42702);
  not i42707(x42707, x42706);
  not i42713(x42713, x41391);
  not i42714(x42714, x41382);
  not i42717(x42717, x42716);
  not i42719(x42719, x41400);
  not i42724(x42724, x41418);
  not i42725(x42725, x41409);
  not i42728(x42728, x42727);
  not i42732(x42732, x42731);
  not i42737(x42737, x42736);
  not i42741(x42741, x42740);
  not i42747(x42747, x41438);
  not i42748(x42748, x41429);
  not i42751(x42751, x42750);
  not i42753(x42753, x41447);
  not i42758(x42758, x41465);
  not i42759(x42759, x41456);
  not i42762(x42762, x42761);
  not i42764(x42764, x41474);
  not i42767(x42767, x42766);
  not i42772(x42772, x42771);
  not i42776(x42776, x42775);
  not i42781(x42781, x42780);
  not i42787(x42787, x41491);
  not i42788(x42788, x41482);
  not i42791(x42791, x42790);
  not i42793(x42793, x41500);
  not i42798(x42798, x41518);
  not i42799(x42799, x41509);
  not i42802(x42802, x42801);
  not i42804(x42804, x41527);
  not i42807(x42807, x42806);
  not i42812(x42812, x42811);
  not i42816(x42816, x42815);
  not i42821(x42821, x42820);
  not i42827(x42827, x41544);
  not i42828(x42828, x41535);
  not i42831(x42831, x42830);
  not i42833(x42833, x41553);
  not i42838(x42838, x41571);
  not i42839(x42839, x41562);
  not i42842(x42842, x42841);
  not i42844(x42844, x41580);
  not i42847(x42847, x42846);
  not i42852(x42852, x42851);
  not i42856(x42856, x42855);
  not i42861(x42861, x42860);
  not i42867(x42867, x41600);
  not i42868(x42868, x41591);
  not i42871(x42871, x42870);
  not i42873(x42873, x41609);
  not i42878(x42878, x41627);
  not i42879(x42879, x41618);
  not i42882(x42882, x42881);
  not i42884(x42884, x41636);
  not i42887(x42887, x42886);
  not i42889(x42889, x41645);
  not i42893(x42893, x42892);
  not i42897(x42897, x42896);
  not i42902(x42902, x42901);
  not i42906(x42906, x42905);
  not i42909(x42909, x41662);
  not i42910(x42910, x41653);
  not i42913(x42913, x42912);
  not i42915(x42915, x41671);
  not i42920(x42920, x41689);
  not i42921(x42921, x41680);
  not i42924(x42924, x42923);
  not i42926(x42926, x41698);
  not i42929(x42929, x42928);
  not i42931(x42931, x41707);
  not i42935(x42935, x42934);
  not i42939(x42939, x42938);
  not i42944(x42944, x42943);
  not i42948(x42948, x42947);
  not i42951(x42951, x41724);
  not i42952(x42952, x41715);
  not i42955(x42955, x42954);
  not i42957(x42957, x41733);
  not i42962(x42962, x41751);
  not i42963(x42963, x41742);
  not i42966(x42966, x42965);
  not i42968(x42968, x41760);
  not i42971(x42971, x42970);
  not i42974(x42974, x41769);
  not i42980(x42980, x42979);
  not i42984(x42984, x42983);
  not i42989(x42989, x42988);
  not i42993(x42993, x42992);
  not i42996(x42996, x41789);
  not i42997(x42997, x41780);
  not i43000(x43000, x42999);
  not i43002(x43002, x41798);
  not i43007(x43007, x41816);
  not i43008(x43008, x41807);
  not i43011(x43011, x43010);
  not i43013(x43013, x41825);
  not i43016(x43016, x43015);
  not i43019(x43019, x41842);
  not i43020(x43020, x41834);
  not i43026(x43026, x43025);
  not i43030(x43030, x43029);
  not i43035(x43035, x43034);
  not i43039(x43039, x43038);
  not i43045(x43045, x41859);
  not i43046(x43046, x41850);
  not i43049(x43049, x43048);
  not i43051(x43051, x41868);
  not i43054(x43054, x43053);
  not i43057(x43057, x41886);
  not i43058(x43058, x41877);
  not i43061(x43061, x43060);
  not i43063(x43063, x41895);
  not i43066(x43066, x43065);
  not i43069(x43069, x41913);
  not i43070(x43070, x41904);
  not i43076(x43076, x43075);
  not i43080(x43080, x43079);
  not i43085(x43085, x43084);
  not i43089(x43089, x43088);
  not i43095(x43095, x41930);
  not i43096(x43096, x41921);
  not i43099(x43099, x43098);
  not i43101(x43101, x41939);
  not i43104(x43104, x43103);
  not i43107(x43107, x41957);
  not i43108(x43108, x41948);
  not i43111(x43111, x43110);
  not i43113(x43113, x41966);
  not i43116(x43116, x43115);
  not i43119(x43119, x41984);
  not i43120(x43120, x41975);
  not i43123(x43123, x43122);
  not i43127(x43127, x43126);
  not i43132(x43132, x43131);
  not i43136(x43136, x43135);
  not i43141(x43141, x43140);
  not i43145(x43145, x43144);
  not i43151(x43151, x42004);
  not i43152(x43152, x41995);
  not i43155(x43155, x43154);
  not i43157(x43157, x42013);
  not i43160(x43160, x43159);
  not i43163(x43163, x42031);
  not i43164(x43164, x42022);
  not i43167(x43167, x43166);
  not i43169(x43169, x42040);
  not i43172(x43172, x43171);
  not i43175(x43175, x42058);
  not i43176(x43176, x42049);
  not i43179(x43179, x43178);
  not i43181(x43181, x42067);
  not i43184(x43184, x43183);
  not i43189(x43189, x43188);
  not i43193(x43193, x43192);
  not i43198(x43198, x43197);
  not i43202(x43202, x43201);
  not i43207(x43207, x43206);
  not i43211(x43211, x43210);
  not i43214(x43214, x42084);
  not i43215(x43215, x42075);
  not i43218(x43218, x43217);
  not i43220(x43220, x42093);
  not i43223(x43223, x43222);
  not i43226(x43226, x42111);
  not i43227(x43227, x42102);
  not i43230(x43230, x43229);
  not i43232(x43232, x42120);
  not i43235(x43235, x43234);
  not i43238(x43238, x42138);
  not i43239(x43239, x42129);
  not i43242(x43242, x43241);
  not i43244(x43244, x42147);
  not i43247(x43247, x43246);
  not i43252(x43252, x43251);
  not i43256(x43256, x43255);
  not i43261(x43261, x43260);
  not i43265(x43265, x43264);
  not i43270(x43270, x43269);
  not i43274(x43274, x43273);
  not i43277(x43277, x42164);
  not i43278(x43278, x42155);
  not i43281(x43281, x43280);
  not i43283(x43283, x42173);
  not i43286(x43286, x43285);
  not i43289(x43289, x42191);
  not i43290(x43290, x42182);
  not i43293(x43293, x43292);
  not i43295(x43295, x42200);
  not i43298(x43298, x43297);
  not i43301(x43301, x42218);
  not i43302(x43302, x42209);
  not i43305(x43305, x43304);
  not i43307(x43307, x42227);
  not i43310(x43310, x43309);
  not i43315(x43315, x43314);
  not i43319(x43319, x43318);
  not i43323(x43323, x43322);
  not i43328(x43328, x43327);
  not i43332(x43332, x43331);
  not i43337(x43337, x43336);
  not i43341(x43341, x43340);
  not i43344(x43344, x42248);
  not i43345(x43345, x42239);
  not i43348(x43348, x43347);
  not i43350(x43350, x42257);
  not i43353(x43353, x43352);
  not i43356(x43356, x42275);
  not i43357(x43357, x42266);
  not i43360(x43360, x43359);
  not i43362(x43362, x42284);
  not i43365(x43365, x43364);
  not i43368(x43368, x42302);
  not i43369(x43369, x42293);
  not i43372(x43372, x43371);
  not i43374(x43374, x42311);
  not i43377(x43377, x43376);
  not i43379(x43379, x42320);
  not i43383(x43383, x43382);
  not i43387(x43387, x43386);
  not i43391(x43391, x43390);
  not i43396(x43396, x43395);
  not i43400(x43400, x43399);
  not i43405(x43405, x43404);
  not i43409(x43409, x43408);
  not i43412(x43412, x42338);
  not i43413(x43413, x42329);
  not i43416(x43416, x43415);
  not i43418(x43418, x42347);
  not i43421(x43421, x43420);
  not i43423(x43423, x42365);
  not i43424(x43424, x42356);
  not i43427(x43427, x43426);
  not i43429(x43429, x42374);
  not i43432(x43432, x43431);
  not i43434(x43434, x42392);
  not i43435(x43435, x42383);
  not i43438(x43438, x43437);
  not i43440(x43440, x42401);
  not i43443(x43443, x43442);
  not i43444(x43444, x42410);
  not i43448(x43448, x43447);
  not i43452(x43452, x43451);
  not i43456(x43456, x43455);
  not i43460(x43460, x43459);
  not i43464(x43464, x43463);
  not i43468(x43468, x43467);
  not i43472(x43472, x43471);
  not i43476(x43476, x43475);
  not i43480(x43480, x43479);
  not i43484(x43484, x43483);
  not i43488(x43488, x43487);
  not i43492(x43492, x43491);
  not i43496(x43496, x43495);
  not i43497(x43497, x42526);
  not i43501(x43501, x43500);
  not i43502(x43502, x42540);
  not i43503(x43503, x42549);
  not i43507(x43507, x43506);
  not i43508(x43508, x42560);
  not i43509(x43509, x42569);
  not i43513(x43513, x43512);
  not i43517(x43517, x43516);
  not i43518(x43518, x42580);
  not i43519(x43519, x42589);
  not i43523(x43523, x43522);
  not i43527(x43527, x43526);
  not i43528(x43528, x42600);
  not i43529(x43529, x42610);
  not i43533(x43533, x43532);
  not i43537(x43537, x43536);
  not i43538(x43538, x42621);
  not i43539(x43539, x42631);
  not i43543(x43543, x43542);
  not i43547(x43547, x43546);
  not i43549(x43549, x42642);
  not i43552(x43552, x42655);
  not i43556(x43556, x43555);
  not i43560(x43560, x43559);
  not i43562(x43562, x42666);
  not i43565(x43565, x42680);
  not i43569(x43569, x43568);
  not i43573(x43573, x43572);
  not i43577(x43577, x43576);
  not i43579(x43579, x42694);
  not i43582(x43582, x42708);
  not i43586(x43586, x43585);
  not i43590(x43590, x43589);
  not i43594(x43594, x43593);
  not i43596(x43596, x42733);
  not i43597(x43597, x42722);
  not i43600(x43600, x42742);
  not i43604(x43604, x43603);
  not i43608(x43608, x43607);
  not i43612(x43612, x43611);
  not i43614(x43614, x42768);
  not i43615(x43615, x42756);
  not i43618(x43618, x42777);
  not i43620(x43620, x42785);
  not i43623(x43623, x43622);
  not i43627(x43627, x43626);
  not i43631(x43631, x43630);
  not i43633(x43633, x42808);
  not i43634(x43634, x42796);
  not i43637(x43637, x42817);
  not i43639(x43639, x42825);
  not i43642(x43642, x43641);
  not i43646(x43646, x43645);
  not i43650(x43650, x43649);
  not i43654(x43654, x43653);
  not i43657(x43657, x42848);
  not i43658(x43658, x42836);
  not i43661(x43661, x42857);
  not i43663(x43663, x42865);
  not i43666(x43666, x43665);
  not i43670(x43670, x43669);
  not i43674(x43674, x43673);
  not i43678(x43678, x43677);
  not i43684(x43684, x42888);
  not i43685(x43685, x42876);
  not i43688(x43688, x42898);
  not i43690(x43690, x42907);
  not i43693(x43693, x43692);
  not i43697(x43697, x43696);
  not i43701(x43701, x43700);
  not i43705(x43705, x43704);
  not i43711(x43711, x42930);
  not i43712(x43712, x42918);
  not i43715(x43715, x42940);
  not i43717(x43717, x42949);
  not i43720(x43720, x43719);
  not i43724(x43724, x43723);
  not i43728(x43728, x43727);
  not i43732(x43732, x43731);
  not i43738(x43738, x42972);
  not i43739(x43739, x42960);
  not i43742(x43742, x43741);
  not i43746(x43746, x43745);
  not i43748(x43748, x42985);
  not i43750(x43750, x42994);
  not i43753(x43753, x43752);
  not i43757(x43757, x43756);
  not i43761(x43761, x43760);
  not i43765(x43765, x43764);
  not i43771(x43771, x43017);
  not i43772(x43772, x43005);
  not i43775(x43775, x43774);
  not i43779(x43779, x43778);
  not i43781(x43781, x43031);
  not i43783(x43783, x43040);
  not i43786(x43786, x43785);
  not i43790(x43790, x43789);
  not i43794(x43794, x43793);
  not i43799(x43799, x43798);
  not i43803(x43803, x43802);
  not i43809(x43809, x43067);
  not i43810(x43810, x43055);
  not i43813(x43813, x43812);
  not i43817(x43817, x43816);
  not i43819(x43819, x43081);
  not i43821(x43821, x43090);
  not i43824(x43824, x43823);
  not i43828(x43828, x43827);
  not i43832(x43832, x43831);
  not i43837(x43837, x43836);
  not i43841(x43841, x43840);
  not i43847(x43847, x43117);
  not i43848(x43848, x43105);
  not i43851(x43851, x43850);
  not i43853(x43853, x43128);
  not i43856(x43856, x43855);
  not i43858(x43858, x43137);
  not i43860(x43860, x43146);
  not i43863(x43863, x43862);
  not i43867(x43867, x43866);
  not i43871(x43871, x43870);
  not i43876(x43876, x43875);
  not i43880(x43880, x43879);
  not i43886(x43886, x43173);
  not i43887(x43887, x43161);
  not i43890(x43890, x43889);
  not i43892(x43892, x43185);
  not i43895(x43895, x43894);
  not i43897(x43897, x43194);
  not i43899(x43899, x43203);
  not i43902(x43902, x43901);
  not i43904(x43904, x43212);
  not i43907(x43907, x43906);
  not i43911(x43911, x43910);
  not i43916(x43916, x43915);
  not i43920(x43920, x43919);
  not i43926(x43926, x43236);
  not i43927(x43927, x43224);
  not i43930(x43930, x43929);
  not i43932(x43932, x43248);
  not i43935(x43935, x43934);
  not i43937(x43937, x43257);
  not i43939(x43939, x43266);
  not i43942(x43942, x43941);
  not i43944(x43944, x43275);
  not i43947(x43947, x43946);
  not i43951(x43951, x43950);
  not i43956(x43956, x43955);
  not i43960(x43960, x43959);
  not i43966(x43966, x43299);
  not i43967(x43967, x43287);
  not i43970(x43970, x43969);
  not i43972(x43972, x43311);
  not i43975(x43975, x43974);
  not i43978(x43978, x43324);
  not i43981(x43981, x43980);
  not i43983(x43983, x43333);
  not i43986(x43986, x43985);
  not i43989(x43989, x43342);
  not i43992(x43992, x43991);
  not i43996(x43996, x43995);
  not i44001(x44001, x44000);
  not i44005(x44005, x44004);
  not i44010(x44010, x44009);
  not i44014(x44014, x44013);
  not i44017(x44017, x43366);
  not i44018(x44018, x43354);
  not i44021(x44021, x44020);
  not i44023(x44023, x43378);
  not i44026(x44026, x44025);
  not i44028(x44028, x43392);
  not i44031(x44031, x44030);
  not i44033(x44033, x43401);
  not i44036(x44036, x44035);
  not i44038(x44038, x43410);
  not i44041(x44041, x44040);
  not i44045(x44045, x44044);
  not i44049(x44049, x44048);
  not i44053(x44053, x44052);
  not i44057(x44057, x44056);
  not i44061(x44061, x44060);
  not i44071(x44071, x44070);
  not i44075(x44075, x44074);
  not i44082(x44082, x44081);
  not i44089(x44089, x44088);
  not i44093(x44093, x44092);
  not i44101(x44101, x44100);
  not i44105(x44105, x44104);
  not i44113(x44113, x44112);
  not i44117(x44117, x44116);
  not i44125(x44125, x44124);
  not i44129(x44129, x44128);
  not i44137(x44137, x44136);
  not i44141(x44141, x44140);
  not i44146(x44146, x44145);
  not i44150(x44150, x44149);
  not i44154(x44154, x44153);
  not i44159(x44159, x44158);
  not i44163(x44163, x44162);
  not i44167(x44167, x44166);
  not i44172(x44172, x44171);
  not i44176(x44176, x44175);
  not i44180(x44180, x44179);
  not i44185(x44185, x44184);
  not i44189(x44189, x44188);
  not i44193(x44193, x44192);
  not i44198(x44198, x44197);
  not i44202(x44202, x44201);
  not i44206(x44206, x44205);
  not i44210(x44210, x44209);
  not i44215(x44215, x44214);
  not i44219(x44219, x44218);
  not i44224(x44224, x44223);
  not i44228(x44228, x44227);
  not i44232(x44232, x44231);
  not i44237(x44237, x44236);
  not i44241(x44241, x44240);
  not i44246(x44246, x44245);
  not i44250(x44250, x44249);
  not i44254(x44254, x44253);
  not i44259(x44259, x44258);
  not i44263(x44263, x44262);
  not i44268(x44268, x44267);
  not i44272(x44272, x44271);
  not i44276(x44276, x44275);
  not i44281(x44281, x44280);
  not i44285(x44285, x44284);
  not i44290(x44290, x44289);
  not i44294(x44294, x44293);
  not i44298(x44298, x44297);
  not i44303(x44303, x44302);
  not i44307(x44307, x44306);
  not i44309(x44309, x43655);
  not i44313(x44313, x44312);
  not i44317(x44317, x44316);
  not i44321(x44321, x44320);
  not i44326(x44326, x44325);
  not i44330(x44330, x44329);
  not i44333(x44333, x43679);
  not i44336(x44336, x44335);
  not i44340(x44340, x44339);
  not i44345(x44345, x44344);
  not i44349(x44349, x44348);
  not i44354(x44354, x44353);
  not i44358(x44358, x44357);
  not i44361(x44361, x43706);
  not i44364(x44364, x44363);
  not i44368(x44368, x44367);
  not i44373(x44373, x44372);
  not i44377(x44377, x44376);
  not i44382(x44382, x44381);
  not i44386(x44386, x44385);
  not i44389(x44389, x43733);
  not i44392(x44392, x44391);
  not i44396(x44396, x44395);
  not i44401(x44401, x44400);
  not i44405(x44405, x44404);
  not i44408(x44408, x43747);
  not i44411(x44411, x44410);
  not i44415(x44415, x44414);
  not i44418(x44418, x43766);
  not i44421(x44421, x44420);
  not i44425(x44425, x44424);
  not i44430(x44430, x44429);
  not i44434(x44434, x44433);
  not i44437(x44437, x43780);
  not i44440(x44440, x44439);
  not i44442(x44442, x43795);
  not i44445(x44445, x44444);
  not i44448(x44448, x43804);
  not i44451(x44451, x44450);
  not i44455(x44455, x44454);
  not i44460(x44460, x44459);
  not i44464(x44464, x44463);
  not i44467(x44467, x43818);
  not i44470(x44470, x44469);
  not i44472(x44472, x43833);
  not i44475(x44475, x44474);
  not i44478(x44478, x43842);
  not i44481(x44481, x44480);
  not i44485(x44485, x44484);
  not i44490(x44490, x44489);
  not i44494(x44494, x44493);
  not i44497(x44497, x43857);
  not i44500(x44500, x44499);
  not i44502(x44502, x43872);
  not i44505(x44505, x44504);
  not i44508(x44508, x43881);
  not i44511(x44511, x44510);
  not i44515(x44515, x44514);
  not i44520(x44520, x44519);
  not i44524(x44524, x44523);
  not i44527(x44527, x43896);
  not i44530(x44530, x44529);
  not i44532(x44532, x43912);
  not i44535(x44535, x44534);
  not i44538(x44538, x43921);
  not i44541(x44541, x44540);
  not i44545(x44545, x44544);
  not i44550(x44550, x44549);
  not i44554(x44554, x44553);
  not i44557(x44557, x43936);
  not i44560(x44560, x44559);
  not i44562(x44562, x43952);
  not i44565(x44565, x44564);
  not i44568(x44568, x43961);
  not i44571(x44571, x44570);
  not i44575(x44575, x44574);
  not i44580(x44580, x44579);
  not i44584(x44584, x44583);
  not i44587(x44587, x43987);
  not i44588(x44588, x43976);
  not i44591(x44591, x44590);
  not i44593(x44593, x43997);
  not i44596(x44596, x44595);
  not i44598(x44598, x44015);
  not i44599(x44599, x44006);
  not i44602(x44602, x44601);
  not i44606(x44606, x44605);
  not i44610(x44610, x44609);
  not i44614(x44614, x44613);
  not i44627(x44627, x44626);
  not i44632(x44632, x44094);
  not i44635(x44635, x44634);
  not i44640(x44640, x44106);
  not i44643(x44643, x44642);
  not i44648(x44648, x44118);
  not i44651(x44651, x44650);
  not i44656(x44656, x44130);
  not i44659(x44659, x44658);
  not i44664(x44664, x44142);
  not i44667(x44667, x44666);
  not i44671(x44671, x44670);
  not i44675(x44675, x44674);
  not i44678(x44678, x44155);
  not i44681(x44681, x44680);
  not i44685(x44685, x44684);
  not i44689(x44689, x44688);
  not i44692(x44692, x44168);
  not i44695(x44695, x44694);
  not i44699(x44699, x44698);
  not i44703(x44703, x44702);
  not i44706(x44706, x44181);
  not i44709(x44709, x44708);
  not i44713(x44713, x44712);
  not i44717(x44717, x44716);
  not i44720(x44720, x44194);
  not i44723(x44723, x44722);
  not i44727(x44727, x44726);
  not i44731(x44731, x44730);
  not i44736(x44736, x44735);
  not i44738(x44738, x44211);
  not i44741(x44741, x44740);
  not i44746(x44746, x44745);
  not i44750(x44750, x44749);
  not i44753(x44753, x44220);
  not i44756(x44756, x44755);
  not i44758(x44758, x44233);
  not i44761(x44761, x44760);
  not i44766(x44766, x44765);
  not i44770(x44770, x44769);
  not i44773(x44773, x44242);
  not i44776(x44776, x44775);
  not i44778(x44778, x44255);
  not i44781(x44781, x44780);
  not i44786(x44786, x44785);
  not i44790(x44790, x44789);
  not i44793(x44793, x44264);
  not i44796(x44796, x44795);
  not i44798(x44798, x44277);
  not i44801(x44801, x44800);
  not i44806(x44806, x44805);
  not i44810(x44810, x44809);
  not i44813(x44813, x44286);
  not i44816(x44816, x44815);
  not i44818(x44818, x44299);
  not i44821(x44821, x44820);
  not i44826(x44826, x44825);
  not i44830(x44830, x44829);
  not i44833(x44833, x44308);
  not i44836(x44836, x44835);
  not i44838(x44838, x44322);
  not i44841(x44841, x44840);
  not i44846(x44846, x44845);
  not i44850(x44850, x44849);
  not i44853(x44853, x44341);
  not i44854(x44854, x44331);
  not i44857(x44857, x44856);
  not i44859(x44859, x44350);
  not i44862(x44862, x44861);
  not i44867(x44867, x44866);
  not i44871(x44871, x44870);
  not i44874(x44874, x44369);
  not i44875(x44875, x44359);
  not i44878(x44878, x44877);
  not i44880(x44880, x44378);
  not i44883(x44883, x44882);
  not i44888(x44888, x44887);
  not i44892(x44892, x44891);
  not i44895(x44895, x44397);
  not i44896(x44896, x44387);
  not i44899(x44899, x44898);
  not i44901(x44901, x44406);
  not i44904(x44904, x44903);
  not i44909(x44909, x44908);
  not i44913(x44913, x44912);
  not i44916(x44916, x44426);
  not i44917(x44917, x44416);
  not i44920(x44920, x44919);
  not i44922(x44922, x44435);
  not i44925(x44925, x44924);
  not i44930(x44930, x44929);
  not i44934(x44934, x44933);
  not i44937(x44937, x44456);
  not i44938(x44938, x44446);
  not i44941(x44941, x44940);
  not i44943(x44943, x44465);
  not i44946(x44946, x44945);
  not i44951(x44951, x44950);
  not i44955(x44955, x44954);
  not i44958(x44958, x44486);
  not i44959(x44959, x44476);
  not i44962(x44962, x44961);
  not i44964(x44964, x44495);
  not i44967(x44967, x44966);
  not i44972(x44972, x44971);
  not i44976(x44976, x44975);
  not i44979(x44979, x44516);
  not i44980(x44980, x44506);
  not i44983(x44983, x44982);
  not i44985(x44985, x44525);
  not i44988(x44988, x44987);
  not i44993(x44993, x44992);
  not i44997(x44997, x44996);
  not i45000(x45000, x44546);
  not i45001(x45001, x44536);
  not i45004(x45004, x45003);
  not i45006(x45006, x44555);
  not i45009(x45009, x45008);
  not i45014(x45014, x45013);
  not i45018(x45018, x45017);
  not i45021(x45021, x44576);
  not i45022(x45022, x44566);
  not i45025(x45025, x45024);
  not i45027(x45027, x44585);
  not i45030(x45030, x45029);
  not i45034(x45034, x45033);
  not i45038(x45038, x45037);
  not i45045(x45045, x45044);
  not i45049(x45049, x45048);
  not i45053(x45053, x45052);
  not i45057(x45057, x45056);
  not i45062(x45062, x45061);
  not i45066(x45066, x45065);
  not i45071(x45071, x45070);
  not i45075(x45075, x45074);
  not i45080(x45080, x45079);
  not i45084(x45084, x45083);
  not i45089(x45089, x45088);
  not i45093(x45093, x45092);
  not i45098(x45098, x45097);
  not i45099(x45099, x45095);
  not i45101(x45101, x44676);
  not i45104(x45104, x45103);
  not i45108(x45108, x45107);
  not i45113(x45113, x45112);
  not i45114(x45114, x45110);
  not i45116(x45116, x44690);
  not i45119(x45119, x45118);
  not i45123(x45123, x45122);
  not i45128(x45128, x45127);
  not i45129(x45129, x45125);
  not i45131(x45131, x44704);
  not i45134(x45134, x45133);
  not i45138(x45138, x45137);
  not i45143(x45143, x45142);
  not i45144(x45144, x45140);
  not i45146(x45146, x44718);
  not i45149(x45149, x45148);
  not i45153(x45153, x45152);
  not i45158(x45158, x45157);
  not i45159(x45159, x45155);
  not i45161(x45161, x44732);
  not i45164(x45164, x45163);
  not i45168(x45168, x45167);
  not i45173(x45173, x45172);
  not i45174(x45174, x45170);
  not i45176(x45176, x44751);
  not i45177(x45177, x44742);
  not i45180(x45180, x45179);
  not i45184(x45184, x45183);
  not i45189(x45189, x45188);
  not i45190(x45190, x45186);
  not i45192(x45192, x44771);
  not i45193(x45193, x44762);
  not i45196(x45196, x45195);
  not i45200(x45200, x45199);
  not i45205(x45205, x45204);
  not i45206(x45206, x45202);
  not i45208(x45208, x44791);
  not i45209(x45209, x44782);
  not i45212(x45212, x45211);
  not i45216(x45216, x45215);
  not i45221(x45221, x45220);
  not i45222(x45222, x45218);
  not i45224(x45224, x44811);
  not i45225(x45225, x44802);
  not i45228(x45228, x45227);
  not i45232(x45232, x45231);
  not i45237(x45237, x45236);
  not i45238(x45238, x45234);
  not i45240(x45240, x44831);
  not i45241(x45241, x44822);
  not i45244(x45244, x45243);
  not i45248(x45248, x45247);
  not i45253(x45253, x45252);
  not i45254(x45254, x45250);
  not i45256(x45256, x44851);
  not i45257(x45257, x44842);
  not i45260(x45260, x45259);
  not i45264(x45264, x45263);
  not i45269(x45269, x45268);
  not i45270(x45270, x45266);
  not i45272(x45272, x44872);
  not i45273(x45273, x44863);
  not i45276(x45276, x45275);
  not i45280(x45280, x45279);
  not i45285(x45285, x45284);
  not i45286(x45286, x45282);
  not i45288(x45288, x44893);
  not i45289(x45289, x44884);
  not i45292(x45292, x45291);
  not i45296(x45296, x45295);
  not i45301(x45301, x45300);
  not i45302(x45302, x45298);
  not i45304(x45304, x44914);
  not i45305(x45305, x44905);
  not i45308(x45308, x45307);
  not i45312(x45312, x45311);
  not i45317(x45317, x45316);
  not i45318(x45318, x45314);
  not i45320(x45320, x44935);
  not i45321(x45321, x44926);
  not i45324(x45324, x45323);
  not i45328(x45328, x45327);
  not i45333(x45333, x45332);
  not i45334(x45334, x45330);
  not i45336(x45336, x44956);
  not i45337(x45337, x44947);
  not i45340(x45340, x45339);
  not i45344(x45344, x45343);
  not i45349(x45349, x45348);
  not i45350(x45350, x45346);
  not i45352(x45352, x44977);
  not i45353(x45353, x44968);
  not i45356(x45356, x45355);
  not i45360(x45360, x45359);
  not i45365(x45365, x45364);
  not i45366(x45366, x45362);
  not i45368(x45368, x44998);
  not i45369(x45369, x44989);
  not i45372(x45372, x45371);
  not i45376(x45376, x45375);
  not i45381(x45381, x45380);
  not i45382(x45382, x45378);
  not i45384(x45384, x45019);
  not i45385(x45385, x45010);
  not i45388(x45388, x45387);
  not i45392(x45392, x45391);
  not i45396(x45396, x45395);
  not i45406(x45406, x45405);
  not i45410(x45410, x45409);
  not i45411(x45411, x45058);
  not i45415(x45415, x45414);
  not i45416(x45416, x45067);
  not i45420(x45420, x45419);
  not i45421(x45421, x45076);
  not i45425(x45425, x45424);
  not i45426(x45426, x45085);
  not i45430(x45430, x45429);
  not i45432(x45432, x45094);
  not i45435(x45435, x45434);
  not i45439(x45439, x45438);
  not i45442(x45442, x45109);
  not i45445(x45445, x45444);
  not i45449(x45449, x45448);
  not i45452(x45452, x45124);
  not i45455(x45455, x45454);
  not i45459(x45459, x45458);
  not i45462(x45462, x45139);
  not i45465(x45465, x45464);
  not i45469(x45469, x45468);
  not i45472(x45472, x45154);
  not i45475(x45475, x45474);
  not i45479(x45479, x45478);
  not i45482(x45482, x45169);
  not i45485(x45485, x45484);
  not i45489(x45489, x45488);
  not i45492(x45492, x45185);
  not i45495(x45495, x45494);
  not i45499(x45499, x45498);
  not i45502(x45502, x45201);
  not i45505(x45505, x45504);
  not i45509(x45509, x45508);
  not i45512(x45512, x45217);
  not i45515(x45515, x45514);
  not i45519(x45519, x45518);
  not i45522(x45522, x45233);
  not i45525(x45525, x45524);
  not i45529(x45529, x45528);
  not i45532(x45532, x45249);
  not i45535(x45535, x45534);
  not i45539(x45539, x45538);
  not i45542(x45542, x45265);
  not i45545(x45545, x45544);
  not i45549(x45549, x45548);
  not i45552(x45552, x45281);
  not i45555(x45555, x45554);
  not i45559(x45559, x45558);
  not i45562(x45562, x45297);
  not i45565(x45565, x45564);
  not i45569(x45569, x45568);
  not i45572(x45572, x45313);
  not i45575(x45575, x45574);
  not i45579(x45579, x45578);
  not i45582(x45582, x45329);
  not i45585(x45585, x45584);
  not i45589(x45589, x45588);
  not i45592(x45592, x45345);
  not i45595(x45595, x45594);
  not i45599(x45599, x45598);
  not i45602(x45602, x45361);
  not i45605(x45605, x45604);
  not i45609(x45609, x45608);
  not i45612(x45612, x45377);
  not i45615(x45615, x45614);
  not i45619(x45619, x45618);
  not i45623(x45623, x45622);
  not i45631(x45631, x45630);
  not i45635(x45635, x45634);
  not i45639(x45639, x45638);
  not i45643(x45643, x45642);
  not i45648(x45648, x45647);
  not i45652(x45652, x45651);
  not i45657(x45657, x45656);
  not i45661(x45661, x45660);
  not i45666(x45666, x45665);
  not i45670(x45670, x45669);
  not i45675(x45675, x45674);
  not i45679(x45679, x45678);
  not i45684(x45684, x45683);
  not i45688(x45688, x45687);
  not i45693(x45693, x45692);
  not i45697(x45697, x45696);
  not i45700(x45700, x45440);
  not i45703(x45703, x45702);
  not i45707(x45707, x45706);
  not i45710(x45710, x45450);
  not i45713(x45713, x45712);
  not i45717(x45717, x45716);
  not i45720(x45720, x45460);
  not i45723(x45723, x45722);
  not i45727(x45727, x45726);
  not i45730(x45730, x45470);
  not i45733(x45733, x45732);
  not i45737(x45737, x45736);
  not i45740(x45740, x45480);
  not i45743(x45743, x45742);
  not i45747(x45747, x45746);
  not i45750(x45750, x45490);
  not i45753(x45753, x45752);
  not i45757(x45757, x45756);
  not i45760(x45760, x45500);
  not i45763(x45763, x45762);
  not i45767(x45767, x45766);
  not i45770(x45770, x45510);
  not i45773(x45773, x45772);
  not i45777(x45777, x45776);
  not i45780(x45780, x45520);
  not i45783(x45783, x45782);
  not i45787(x45787, x45786);
  not i45790(x45790, x45530);
  not i45793(x45793, x45792);
  not i45797(x45797, x45796);
  not i45800(x45800, x45540);
  not i45803(x45803, x45802);
  not i45807(x45807, x45806);
  not i45810(x45810, x45550);
  not i45813(x45813, x45812);
  not i45817(x45817, x45816);
  not i45820(x45820, x45560);
  not i45823(x45823, x45822);
  not i45827(x45827, x45826);
  not i45830(x45830, x45570);
  not i45833(x45833, x45832);
  not i45837(x45837, x45836);
  not i45840(x45840, x45580);
  not i45843(x45843, x45842);
  not i45847(x45847, x45846);
  not i45850(x45850, x45590);
  not i45853(x45853, x45852);
  not i45857(x45857, x45856);
  not i45860(x45860, x45600);
  not i45863(x45863, x45862);
  not i45867(x45867, x45866);
  not i45870(x45870, x45610);
  not i45873(x45873, x45872);
  not i45877(x45877, x45876);
  not i45879(x45879, x45627);
  not i45885(x45885, x45884);
  not i45889(x45889, x45888);
  not i45891(x45891, x45644);
  not i45894(x45894, x45893);
  not i45896(x45896, x45653);
  not i45899(x45899, x45898);
  not i45901(x45901, x45662);
  not i45904(x45904, x45903);
  not i45906(x45906, x45671);
  not i45909(x45909, x45908);
  not i45911(x45911, x45680);
  not i45914(x45914, x45913);
  not i45916(x45916, x45689);
  not i45919(x45919, x45918);
  not i45921(x45921, x45698);
  not i45924(x45924, x45923);
  not i45926(x45926, x45708);
  not i45929(x45929, x45928);
  not i45931(x45931, x45718);
  not i45934(x45934, x45933);
  not i45936(x45936, x45728);
  not i45939(x45939, x45938);
  not i45941(x45941, x45738);
  not i45944(x45944, x45943);
  not i45946(x45946, x45748);
  not i45949(x45949, x45948);
  not i45951(x45951, x45758);
  not i45954(x45954, x45953);
  not i45956(x45956, x45768);
  not i45959(x45959, x45958);
  not i45961(x45961, x45778);
  not i45964(x45964, x45963);
  not i45966(x45966, x45788);
  not i45969(x45969, x45968);
  not i45971(x45971, x45798);
  not i45974(x45974, x45973);
  not i45976(x45976, x45808);
  not i45979(x45979, x45978);
  not i45981(x45981, x45818);
  not i45984(x45984, x45983);
  not i45986(x45986, x45828);
  not i45989(x45989, x45988);
  not i45991(x45991, x45838);
  not i45994(x45994, x45993);
  not i45996(x45996, x45848);
  not i45999(x45999, x45998);
  not i46001(x46001, x45858);
  not i46004(x46004, x46003);
  not i46006(x46006, x45868);
  not i46009(x46009, x46008);
  not i46010(x46010, x45878);
  not i46011(x46011, x45882);
  not i46012(x46012, x45886);
  not i46013(x46013, x45890);
  not i46014(x46014, x45895);
  not i46015(x46015, x45900);
  not i46016(x46016, x45905);
  not i46017(x46017, x45910);
  not i46018(x46018, x45915);
  not i46019(x46019, x45920);
  not i46020(x46020, x45925);
  not i46021(x46021, x45930);
  not i46022(x46022, x45935);
  not i46023(x46023, x45940);
  not i46024(x46024, x45945);
  not i46025(x46025, x45950);
  not i46026(x46026, x45955);
  not i46027(x46027, x45960);
  not i46028(x46028, x45965);
  not i46029(x46029, x45970);
  not i46030(x46030, x45975);
  not i46031(x46031, x45980);
  not i46032(x46032, x45985);
  not i46033(x46033, x45990);
  not i46034(x46034, x45995);
  not i46040(x46040, x46039);
  not i46044(x46044, x46043);
  not i46048(x46048, x46047);
  not i46052(x46052, x46051);
  not i46056(x46056, x46055);
  not i46060(x46060, x46059);
  not i46064(x46064, x46063);
  not i46068(x46068, x46067);
  not i46072(x46072, x46071);
  not i46076(x46076, x46075);
  not i46080(x46080, x46079);
  not i46084(x46084, x46083);
  not i46088(x46088, x46087);
  not i46092(x46092, x46091);
  not i46096(x46096, x46095);
  not i46100(x46100, x46099);
  not i46104(x46104, x46103);
  not i46108(x46108, x46107);
  not i46112(x46112, x46111);
  not i46116(x46116, x46115);
  not i46120(x46120, x46119);
  not i46124(x46124, x46123);
  not i46128(x46128, x46127);
  not i46132(x46132, x46131);
  not i46133(x46133, x46036);
  not i46135(x46135, x46038);
  not i46138(x46138, x46042);
  not i46141(x46141, x46046);
  not i46144(x46144, x46143);
  not i46146(x46146, x46050);
  not i46149(x46149, x46148);
  not i46151(x46151, x46054);
  not i46154(x46154, x46153);
  not i46156(x46156, x46058);
  not i46159(x46159, x46158);
  not i46161(x46161, x46062);
  not i46164(x46164, x46163);
  not i46166(x46166, x46066);
  not i46169(x46169, x46168);
  not i46171(x46171, x46070);
  not i46174(x46174, x46173);
  not i46176(x46176, x46074);
  not i46179(x46179, x46178);
  not i46181(x46181, x46078);
  not i46184(x46184, x46183);
  not i46186(x46186, x46082);
  not i46189(x46189, x46188);
  not i46191(x46191, x46086);
  not i46194(x46194, x46193);
  not i46196(x46196, x46090);
  not i46199(x46199, x46198);
  not i46201(x46201, x46094);
  not i46204(x46204, x46203);
  not i46206(x46206, x46098);
  not i46209(x46209, x46208);
  not i46211(x46211, x46102);
  not i46214(x46214, x46213);
  not i46216(x46216, x46106);
  not i46219(x46219, x46218);
  not i46221(x46221, x46110);
  not i46224(x46224, x46223);
  not i46226(x46226, x46114);
  not i46229(x46229, x46228);
  not i46231(x46231, x46118);
  not i46234(x46234, x46233);
  not i46236(x46236, x46122);
  not i46239(x46239, x46238);
  not i46241(x46241, x46126);
  not i46244(x46244, x46243);
  not i46246(x46246, x46130);
  not i46249(x46249, x46248);
  not i46250(x46250, x46136);
  not i46251(x46251, x46139);
  not i46253(x46253, x46142);
  not i46256(x46256, x46147);
  not i46259(x46259, x46152);
  not i46262(x46262, x46157);
  not i46265(x46265, x46162);
  not i46268(x46268, x46267);
  not i46270(x46270, x46167);
  not i46273(x46273, x46272);
  not i46275(x46275, x46172);
  not i46278(x46278, x46277);
  not i46280(x46280, x46177);
  not i46283(x46283, x46282);
  not i46285(x46285, x46182);
  not i46288(x46288, x46287);
  not i46290(x46290, x46187);
  not i46293(x46293, x46292);
  not i46295(x46295, x46192);
  not i46298(x46298, x46297);
  not i46300(x46300, x46197);
  not i46303(x46303, x46302);
  not i46305(x46305, x46202);
  not i46308(x46308, x46307);
  not i46310(x46310, x46207);
  not i46313(x46313, x46312);
  not i46315(x46315, x46212);
  not i46318(x46318, x46317);
  not i46320(x46320, x46217);
  not i46323(x46323, x46322);
  not i46325(x46325, x46222);
  not i46328(x46328, x46327);
  not i46330(x46330, x46227);
  not i46333(x46333, x46332);
  not i46335(x46335, x46232);
  not i46338(x46338, x46337);
  not i46340(x46340, x46237);
  not i46343(x46343, x46342);
  not i46345(x46345, x46242);
  not i46348(x46348, x46347);
  not i46350(x46350, x46247);
  not i46353(x46353, x46352);
  not i46354(x46354, x46254);
  not i46355(x46355, x46257);
  not i46356(x46356, x46260);
  not i46357(x46357, x46263);
  not i46359(x46359, x46266);
  not i46362(x46362, x46271);
  not i46365(x46365, x46276);
  not i46368(x46368, x46281);
  not i46371(x46371, x46286);
  not i46374(x46374, x46291);
  not i46377(x46377, x46296);
  not i46380(x46380, x46301);
  not i46383(x46383, x46306);
  not i46386(x46386, x46385);
  not i46388(x46388, x46311);
  not i46391(x46391, x46390);
  not i46393(x46393, x46316);
  not i46396(x46396, x46395);
  not i46398(x46398, x46321);
  not i46401(x46401, x46400);
  not i46403(x46403, x46326);
  not i46406(x46406, x46405);
  not i46408(x46408, x46331);
  not i46411(x46411, x46410);
  not i46413(x46413, x46336);
  not i46416(x46416, x46415);
  not i46418(x46418, x46341);
  not i46421(x46421, x46420);
  not i46423(x46423, x46346);
  not i46426(x46426, x46425);
  not i46428(x46428, x46351);
  not i46431(x46431, x46430);
  not i46432(x46432, x46366);
  not i46433(x46433, x46369);
  not i46434(x46434, x46372);
  not i46435(x46435, x46375);
  not i46436(x46436, x46378);
  not i46437(x46437, x46381);
  not i46439(x46439, x46384);
  not i46442(x46442, x46389);
  not i46445(x46445, x46394);
  not i46448(x46448, x46399);
  not i46451(x46451, x46404);
  not i46454(x46454, x46409);
  not i46457(x46457, x46414);
  not i46460(x46460, x46419);
  not i46463(x46463, x46424);
  not i46466(x46466, x46429);
  not i46470(x46470, x46469);
  not i46474(x46474, x46473);
  not i46478(x46478, x46477);
  not i46482(x46482, x46481);
  not i46486(x46486, x46485);
  not i46490(x46490, x46489);
  not i46494(x46494, x46493);
  not i46498(x46498, x46497);
  not i46500(x46500, x46360);
  not i46503(x46503, x46502);
  not i46505(x46505, x46363);
  not i46508(x46508, x46507);
  not i46512(x46512, x46511);
  not i46516(x46516, x46515);
  not i46520(x46520, x46519);
  not i46524(x46524, x46523);
  not i46528(x46528, x46527);
  not i46532(x46532, x46531);
  not i46534(x46534, x46440);
  not i46537(x46537, x46536);
  not i46539(x46539, x46443);
  not i46542(x46542, x46541);
  not i46544(x46544, x46446);
  not i46547(x46547, x46546);
  not i46549(x46549, x46449);
  not i46552(x46552, x46551);
  not i46554(x46554, x46452);
  not i46557(x46557, x46556);
  not i46559(x46559, x46455);
  not i46562(x46562, x46561);
  not i46564(x46564, x46458);
  not i46567(x46567, x46566);
  not i46569(x46569, x46461);
  not i46572(x46572, x46571);
  not i46574(x46574, x46464);
  not i46577(x46577, x46576);
  not i46579(x46579, x46467);
  not i46582(x46582, x46581);
  not i46584(x46584, x46583);
  not i46586(x46586, x46585);
  not i46588(x46588, x46587);
  not i46590(x46590, x46589);
  not i46592(x46592, x46591);
  not i46594(x46594, x46593);
  not i46596(x46596, x46595);
  not i46598(x46598, x46597);
  not i46600(x46600, x46599);
  not i46602(x46602, x46601);
  not i46604(x46604, x46603);
  not i46606(x46606, x46605);
  not i46608(x46608, x46607);
  not i46610(x46610, x46609);
  not i46612(x46612, x46611);
  not i46614(x46614, x46613);
  not i46616(x46616, x46615);
  not i46618(x46618, x46617);
  not i46620(x46620, x46619);
  not i46622(x46622, x46621);
  not i46624(x46624, x46623);
  not i46626(x46626, x46625);
  not i46628(x46628, x46627);
  not i46630(x46630, x46629);
  not i46632(x46632, x46631);
  not i46634(x46634, x46633);
  not i46636(x46636, x46635);
  not i46638(x46638, x46637);
  not i46640(x46640, x46639);
  not i46642(x46642, x46641);
  not i46645(x46645, x46644);
  not i46647(x46647, x46646);
  not i46649(x46649, x46648);
  not i46651(x46651, x46650);
  not i46653(x46653, x46652);
  not i46655(x46655, x46654);
  not i46657(x46657, x46656);
  not i46659(x46659, x46658);
  not i46661(x46661, x46660);
  not i46663(x46663, x46662);
  not i46665(x46665, x46664);
  not i46667(x46667, x46666);
  not i46669(x46669, x46668);
  not i46671(x46671, x46670);
  not i46673(x46673, x46672);
  not i46675(x46675, x46674);
  not i46677(x46677, x46676);
  not i46679(x46679, x46678);
  not i46681(x46681, x46680);
  not i46683(x46683, x46682);
  not i46685(x46685, x46684);
  not i46687(x46687, x46686);
  not i46689(x46689, x46688);
  not i46691(x46691, x46690);
  not i46693(x46693, x46692);
  not i46695(x46695, x46694);
  not i46697(x46697, x46696);
  not i46699(x46699, x46698);
  not i46704(x46704, x46703);
  not i46706(x46706, x46705);
  not i46708(x46708, x46707);
  not i46710(x46710, x46709);
  not i46712(x46712, x46711);
  not i46714(x46714, x46713);
  not i46716(x46716, x46715);
  not i46718(x46718, x46717);
  not i46720(x46720, x46719);
  not i46722(x46722, x46721);
  not i46724(x46724, x46723);
  not i46726(x46726, x46725);
  not i46728(x46728, x46727);
  not i46730(x46730, x46729);
  not i46732(x46732, x46731);
  not i46734(x46734, x46733);
  not i46736(x46736, x46735);
  not i46738(x46738, x46737);
  not i46740(x46740, x46739);
  not i46742(x46742, x46741);
  not i46744(x46744, x46743);
  not i46746(x46746, x46745);
  not i46748(x46748, x46747);
  not i46750(x46750, x46749);
  not i46760(x46760, x46759);
  not i46762(x46762, x46761);
  not i46764(x46764, x46763);
  not i46766(x46766, x46765);
  not i46768(x46768, x46767);
  not i46770(x46770, x46769);
  not i46772(x46772, x46771);
  not i46774(x46774, x46773);
  not i46776(x46776, x46775);
  not i46778(x46778, x46777);
  not i46780(x46780, x46779);
  not i46782(x46782, x46781);
  not i46784(x46784, x46783);
  not i46786(x46786, x46785);
  not i46788(x46788, x46787);
  not i46806(x46806, x46805);
  not i46810(x46810, x46809);
  not i46814(x46814, x46813);
  not i46818(x46818, x46817);
  not i46822(x46822, x46821);
  not i46826(x46826, x46825);
  not i46830(x46830, x46829);
  not i46834(x46834, x46833);
  not i46838(x46838, x46837);
  not i46842(x46842, x46841);
  not i46846(x46846, x46845);
  not i46850(x46850, x46849);
  not i46854(x46854, x46853);
  not i46858(x46858, x46857);
  not i46862(x46862, x46861);
  not i46866(x46866, x46865);
  not i46870(x46870, x46869);
  not i46874(x46874, x46873);
  not i46878(x46878, x46877);
  not i46882(x46882, x46881);
  not i46886(x46886, x46885);
  not i46890(x46890, x46889);
  not i46894(x46894, x46893);
  not i46898(x46898, x46897);
  not i46902(x46902, x46901);
  not i46906(x46906, x46905);
  not i46910(x46910, x46909);
  not i46914(x46914, x46913);
  not i46918(x46918, x46917);
  not i46922(x46922, x46921);
  not i46926(x46926, x46925);
  not i46927(x46927, x39971);
  not i46929(x46929, x46928);
  not i46931(x46931, x46930);
  not i46933(x46933, x46932);
  not i46935(x46935, x46934);
  not i46937(x46937, x46936);
  not i46939(x46939, x46938);
  not i46941(x46941, x46940);
  not i46943(x46943, x46942);
  not i46945(x46945, x46944);
  not i46947(x46947, x46946);
  not i46949(x46949, x46948);
  not i46951(x46951, x46950);
  not i46953(x46953, x46952);
  not i46955(x46955, x46954);
  not i46957(x46957, x46956);
  not i46959(x46959, x46958);
  not i46993(x46993, x46992);
  not i46995(x46995, x46994);
  not i46997(x46997, x46996);
  not i46999(x46999, x46998);
  not i47001(x47001, x47000);
  not i47003(x47003, x47002);
  not i47005(x47005, x47004);
  not i47007(x47007, x47006);
  not i47009(x47009, x47008);
  not i47011(x47011, x47010);
  not i47013(x47013, x47012);
  not i47015(x47015, x47014);
  not i47017(x47017, x47016);
  not i47019(x47019, x47018);
  not i47021(x47021, x47020);
  not i47023(x47023, x47022);
  not i47025(x47025, x47024);
  not i47027(x47027, x47026);
  not i47029(x47029, x47028);
  not i47031(x47031, x47030);
  not i47033(x47033, x47032);
  not i47035(x47035, x47034);
  not i47037(x47037, x47036);
  not i47039(x47039, x47038);
  not i47041(x47041, x47040);
  not i47043(x47043, x47042);
  not i47045(x47045, x47044);
  not i47047(x47047, x47046);
  not i47049(x47049, x47048);
  not i47051(x47051, x47050);
  not i47053(x47053, x47052);
  not i47055(x47055, x47054);
  not i49878(x49878, x49815);
  not i49879(x49879, x49817);
  not i49880(x49880, x49819);
  not i49881(x49881, x49821);
  not i49882(x49882, x49823);
  not i49883(x49883, x49825);
  not i49884(x49884, x49827);
  not i49885(x49885, x49829);
  not i49886(x49886, x49831);
  not i49887(x49887, x49833);
  not i49888(x49888, x49835);
  not i49889(x49889, x49837);
  not i49890(x49890, x49839);
  not i49891(x49891, x49841);
  not i49892(x49892, x49843);
  not i49893(x49893, x49845);
  not i49894(x49894, x49847);
  not i49895(x49895, x49849);
  not i49896(x49896, x49851);
  not i49897(x49897, x49853);
  not i49898(x49898, x49855);
  not i49899(x49899, x49857);
  not i49900(x49900, x49859);
  not i49901(x49901, x49861);
  not i49902(x49902, x49863);
  not i49903(x49903, x49865);
  not i49904(x49904, x49867);
  not i49905(x49905, x49869);
  not i49906(x49906, x49871);
  not i49907(x49907, x49873);
  not i49908(x49908, x49875);
  not i49909(x49909, x49877);
  not i50007(x50007, x49912);
  not i50008(x50008, x73517);
  not i50011(x50011, x50010);
  not i50013(x50013, x49915);
  not i50014(x50014, x73522);
  not i50017(x50017, x50016);
  not i50019(x50019, x49918);
  not i50020(x50020, x73527);
  not i50023(x50023, x50022);
  not i50025(x50025, x49921);
  not i50026(x50026, x73532);
  not i50029(x50029, x50028);
  not i50031(x50031, x49924);
  not i50032(x50032, x73537);
  not i50035(x50035, x50034);
  not i50037(x50037, x49927);
  not i50038(x50038, x73542);
  not i50041(x50041, x50040);
  not i50043(x50043, x49930);
  not i50044(x50044, x73547);
  not i50047(x50047, x50046);
  not i50049(x50049, x49933);
  not i50050(x50050, x73552);
  not i50053(x50053, x50052);
  not i50055(x50055, x49936);
  not i50056(x50056, x73557);
  not i50059(x50059, x50058);
  not i50061(x50061, x49939);
  not i50062(x50062, x73562);
  not i50065(x50065, x50064);
  not i50067(x50067, x49942);
  not i50068(x50068, x73567);
  not i50071(x50071, x50070);
  not i50073(x50073, x49945);
  not i50074(x50074, x73572);
  not i50077(x50077, x50076);
  not i50079(x50079, x49948);
  not i50080(x50080, x73577);
  not i50083(x50083, x50082);
  not i50085(x50085, x49951);
  not i50086(x50086, x73582);
  not i50089(x50089, x50088);
  not i50091(x50091, x49954);
  not i50092(x50092, x73587);
  not i50095(x50095, x50094);
  not i50097(x50097, x49957);
  not i50098(x50098, x73592);
  not i50101(x50101, x50100);
  not i50103(x50103, x49960);
  not i50104(x50104, x73597);
  not i50107(x50107, x50106);
  not i50109(x50109, x49963);
  not i50110(x50110, x73602);
  not i50113(x50113, x50112);
  not i50115(x50115, x49966);
  not i50116(x50116, x73607);
  not i50119(x50119, x50118);
  not i50121(x50121, x49969);
  not i50122(x50122, x73612);
  not i50125(x50125, x50124);
  not i50127(x50127, x49972);
  not i50128(x50128, x73617);
  not i50131(x50131, x50130);
  not i50133(x50133, x49975);
  not i50134(x50134, x73622);
  not i50137(x50137, x50136);
  not i50139(x50139, x49978);
  not i50140(x50140, x73627);
  not i50143(x50143, x50142);
  not i50145(x50145, x49981);
  not i50146(x50146, x73632);
  not i50149(x50149, x50148);
  not i50151(x50151, x49984);
  not i50152(x50152, x73637);
  not i50155(x50155, x50154);
  not i50157(x50157, x49987);
  not i50158(x50158, x73642);
  not i50161(x50161, x50160);
  not i50163(x50163, x49990);
  not i50164(x50164, x73647);
  not i50167(x50167, x50166);
  not i50169(x50169, x49993);
  not i50170(x50170, x73652);
  not i50173(x50173, x50172);
  not i50175(x50175, x49996);
  not i50176(x50176, x73657);
  not i50179(x50179, x50178);
  not i50181(x50181, x49999);
  not i50182(x50182, x73662);
  not i50185(x50185, x50184);
  not i50187(x50187, x50002);
  not i50188(x50188, x73667);
  not i50191(x50191, x50190);
  not i50193(x50193, x50005);
  not i50194(x50194, x73672);
  not i50197(x50197, x50196);
  not i50198(x50198, x50006);
  not i50199(x50199, x50012);
  not i50200(x50200, x50018);
  not i50201(x50201, x50024);
  not i50202(x50202, x50030);
  not i50203(x50203, x50036);
  not i50204(x50204, x50042);
  not i50205(x50205, x50048);
  not i50206(x50206, x50054);
  not i50207(x50207, x50060);
  not i50208(x50208, x50066);
  not i50209(x50209, x50072);
  not i50210(x50210, x50078);
  not i50211(x50211, x50084);
  not i50212(x50212, x50090);
  not i50213(x50213, x50096);
  not i50214(x50214, x50102);
  not i50215(x50215, x50108);
  not i50216(x50216, x50114);
  not i50217(x50217, x50120);
  not i50218(x50218, x50126);
  not i50219(x50219, x50132);
  not i50220(x50220, x50138);
  not i50221(x50221, x50144);
  not i50222(x50222, x50150);
  not i50223(x50223, x50156);
  not i50224(x50224, x50162);
  not i50225(x50225, x50168);
  not i50226(x50226, x50174);
  not i50227(x50227, x50180);
  not i50233(x50233, x50232);
  not i50237(x50237, x50236);
  not i50241(x50241, x50240);
  not i50245(x50245, x50244);
  not i50249(x50249, x50248);
  not i50253(x50253, x50252);
  not i50257(x50257, x50256);
  not i50261(x50261, x50260);
  not i50265(x50265, x50264);
  not i50269(x50269, x50268);
  not i50273(x50273, x50272);
  not i50277(x50277, x50276);
  not i50281(x50281, x50280);
  not i50285(x50285, x50284);
  not i50289(x50289, x50288);
  not i50293(x50293, x50292);
  not i50297(x50297, x50296);
  not i50301(x50301, x50300);
  not i50305(x50305, x50304);
  not i50309(x50309, x50308);
  not i50313(x50313, x50312);
  not i50317(x50317, x50316);
  not i50321(x50321, x50320);
  not i50325(x50325, x50324);
  not i50329(x50329, x50328);
  not i50333(x50333, x50332);
  not i50337(x50337, x50336);
  not i50341(x50341, x50340);
  not i50345(x50345, x50344);
  not i50349(x50349, x50348);
  not i50351(x50351, x50231);
  not i50354(x50354, x50235);
  not i50357(x50357, x50239);
  not i50360(x50360, x50359);
  not i50362(x50362, x50243);
  not i50365(x50365, x50364);
  not i50367(x50367, x50247);
  not i50370(x50370, x50369);
  not i50372(x50372, x50251);
  not i50375(x50375, x50374);
  not i50377(x50377, x50255);
  not i50380(x50380, x50379);
  not i50382(x50382, x50259);
  not i50385(x50385, x50384);
  not i50387(x50387, x50263);
  not i50390(x50390, x50389);
  not i50392(x50392, x50267);
  not i50395(x50395, x50394);
  not i50397(x50397, x50271);
  not i50400(x50400, x50399);
  not i50402(x50402, x50275);
  not i50405(x50405, x50404);
  not i50407(x50407, x50279);
  not i50410(x50410, x50409);
  not i50412(x50412, x50283);
  not i50415(x50415, x50414);
  not i50417(x50417, x50287);
  not i50420(x50420, x50419);
  not i50422(x50422, x50291);
  not i50425(x50425, x50424);
  not i50427(x50427, x50295);
  not i50430(x50430, x50429);
  not i50432(x50432, x50299);
  not i50435(x50435, x50434);
  not i50437(x50437, x50303);
  not i50440(x50440, x50439);
  not i50442(x50442, x50307);
  not i50445(x50445, x50444);
  not i50447(x50447, x50311);
  not i50450(x50450, x50449);
  not i50452(x50452, x50315);
  not i50455(x50455, x50454);
  not i50457(x50457, x50319);
  not i50460(x50460, x50459);
  not i50462(x50462, x50323);
  not i50465(x50465, x50464);
  not i50467(x50467, x50327);
  not i50470(x50470, x50469);
  not i50472(x50472, x50331);
  not i50475(x50475, x50474);
  not i50477(x50477, x50335);
  not i50480(x50480, x50479);
  not i50482(x50482, x50339);
  not i50485(x50485, x50484);
  not i50487(x50487, x50343);
  not i50490(x50490, x50489);
  not i50492(x50492, x50347);
  not i50495(x50495, x50494);
  not i50497(x50497, x50358);
  not i50500(x50500, x50363);
  not i50503(x50503, x50368);
  not i50506(x50506, x50373);
  not i50509(x50509, x50378);
  not i50512(x50512, x50511);
  not i50514(x50514, x50383);
  not i50517(x50517, x50516);
  not i50519(x50519, x50388);
  not i50522(x50522, x50521);
  not i50524(x50524, x50393);
  not i50527(x50527, x50526);
  not i50529(x50529, x50398);
  not i50532(x50532, x50531);
  not i50534(x50534, x50403);
  not i50537(x50537, x50536);
  not i50539(x50539, x50408);
  not i50542(x50542, x50541);
  not i50544(x50544, x50413);
  not i50547(x50547, x50546);
  not i50549(x50549, x50418);
  not i50552(x50552, x50551);
  not i50554(x50554, x50423);
  not i50557(x50557, x50556);
  not i50559(x50559, x50428);
  not i50562(x50562, x50561);
  not i50564(x50564, x50433);
  not i50567(x50567, x50566);
  not i50569(x50569, x50438);
  not i50572(x50572, x50571);
  not i50574(x50574, x50443);
  not i50577(x50577, x50576);
  not i50579(x50579, x50448);
  not i50582(x50582, x50581);
  not i50584(x50584, x50453);
  not i50587(x50587, x50586);
  not i50589(x50589, x50458);
  not i50592(x50592, x50591);
  not i50594(x50594, x50463);
  not i50597(x50597, x50596);
  not i50599(x50599, x50468);
  not i50602(x50602, x50601);
  not i50604(x50604, x50473);
  not i50607(x50607, x50606);
  not i50609(x50609, x50478);
  not i50612(x50612, x50611);
  not i50614(x50614, x50483);
  not i50617(x50617, x50616);
  not i50619(x50619, x50488);
  not i50622(x50622, x50621);
  not i50624(x50624, x50493);
  not i50627(x50627, x50626);
  not i50629(x50629, x50510);
  not i50632(x50632, x50515);
  not i50635(x50635, x50520);
  not i50638(x50638, x50525);
  not i50641(x50641, x50530);
  not i50644(x50644, x50535);
  not i50647(x50647, x50540);
  not i50650(x50650, x50545);
  not i50653(x50653, x50550);
  not i50656(x50656, x50655);
  not i50658(x50658, x50555);
  not i50661(x50661, x50660);
  not i50663(x50663, x50560);
  not i50666(x50666, x50665);
  not i50668(x50668, x50565);
  not i50671(x50671, x50670);
  not i50673(x50673, x50570);
  not i50676(x50676, x50675);
  not i50678(x50678, x50575);
  not i50681(x50681, x50680);
  not i50683(x50683, x50580);
  not i50686(x50686, x50685);
  not i50688(x50688, x50585);
  not i50691(x50691, x50690);
  not i50693(x50693, x50590);
  not i50696(x50696, x50695);
  not i50698(x50698, x50595);
  not i50701(x50701, x50700);
  not i50703(x50703, x50600);
  not i50706(x50706, x50705);
  not i50708(x50708, x50605);
  not i50711(x50711, x50710);
  not i50713(x50713, x50610);
  not i50716(x50716, x50715);
  not i50718(x50718, x50615);
  not i50721(x50721, x50720);
  not i50723(x50723, x50620);
  not i50726(x50726, x50725);
  not i50728(x50728, x50625);
  not i50731(x50731, x50730);
  not i50733(x50733, x50654);
  not i50736(x50736, x50659);
  not i50739(x50739, x50664);
  not i50742(x50742, x50669);
  not i50745(x50745, x50674);
  not i50748(x50748, x50679);
  not i50751(x50751, x50684);
  not i50754(x50754, x50689);
  not i50757(x50757, x50694);
  not i50760(x50760, x50699);
  not i50763(x50763, x50704);
  not i50766(x50766, x50709);
  not i50769(x50769, x50714);
  not i50772(x50772, x50719);
  not i50775(x50775, x50724);
  not i50778(x50778, x50729);
  not i50782(x50782, x50781);
  not i50784(x50784, x50229);
  not i50787(x50787, x50786);
  not i50789(x50789, x50352);
  not i50792(x50792, x50791);
  not i50794(x50794, x50355);
  not i50797(x50797, x50796);
  not i50799(x50799, x50498);
  not i50802(x50802, x50801);
  not i50804(x50804, x50501);
  not i50807(x50807, x50806);
  not i50809(x50809, x50504);
  not i50812(x50812, x50811);
  not i50814(x50814, x50507);
  not i50817(x50817, x50816);
  not i50819(x50819, x50630);
  not i50822(x50822, x50821);
  not i50824(x50824, x50633);
  not i50827(x50827, x50826);
  not i50829(x50829, x50636);
  not i50832(x50832, x50831);
  not i50834(x50834, x50639);
  not i50837(x50837, x50836);
  not i50839(x50839, x50642);
  not i50842(x50842, x50841);
  not i50844(x50844, x50645);
  not i50847(x50847, x50846);
  not i50849(x50849, x50648);
  not i50852(x50852, x50851);
  not i50854(x50854, x50651);
  not i50857(x50857, x50856);
  not i50859(x50859, x50734);
  not i50862(x50862, x50861);
  not i50864(x50864, x50737);
  not i50867(x50867, x50866);
  not i50869(x50869, x50740);
  not i50872(x50872, x50871);
  not i50874(x50874, x50743);
  not i50877(x50877, x50876);
  not i50879(x50879, x50746);
  not i50882(x50882, x50881);
  not i50884(x50884, x50749);
  not i50887(x50887, x50886);
  not i50889(x50889, x50752);
  not i50892(x50892, x50891);
  not i50894(x50894, x50755);
  not i50897(x50897, x50896);
  not i50899(x50899, x50758);
  not i50902(x50902, x50901);
  not i50904(x50904, x50761);
  not i50907(x50907, x50906);
  not i50909(x50909, x50764);
  not i50912(x50912, x50911);
  not i50914(x50914, x50767);
  not i50917(x50917, x50916);
  not i50919(x50919, x50770);
  not i50922(x50922, x50921);
  not i50924(x50924, x50773);
  not i50927(x50927, x50926);
  not i50929(x50929, x50776);
  not i50932(x50932, x50931);
  not i50934(x50934, x50779);
  not i50937(x50937, x50936);
  not i50940(x50940, x50939);
  not i50942(x50942, x50941);
  not i50944(x50944, x50943);
  not i50946(x50946, x50945);
  not i50948(x50948, x50947);
  not i50950(x50950, x50949);
  not i50952(x50952, x50951);
  not i50954(x50954, x50953);
  not i50957(x50957, x50956);
  not i50959(x50959, x50958);
  not i50961(x50961, x50960);
  not i50963(x50963, x50962);
  not i50965(x50965, x50964);
  not i50967(x50967, x50966);
  not i50969(x50969, x50968);
  not i50971(x50971, x50970);
  not i50973(x50973, x50972);
  not i50975(x50975, x50974);
  not i50977(x50977, x50976);
  not i50979(x50979, x50978);
  not i50981(x50981, x50980);
  not i50983(x50983, x50982);
  not i50985(x50985, x50984);
  not i50987(x50987, x50986);
  not i50989(x50989, x50988);
  not i50992(x50992, x50991);
  not i50994(x50994, x50993);
  not i50996(x50996, x50995);
  not i50998(x50998, x50997);
  not i51000(x51000, x50999);
  not i51002(x51002, x51001);
  not i51004(x51004, x51003);
  not i51006(x51006, x51005);
  not i51008(x51008, x51007);
  not i51010(x51010, x51009);
  not i51012(x51012, x51011);
  not i51014(x51014, x51013);
  not i51016(x51016, x51015);
  not i51018(x51018, x51017);
  not i51020(x51020, x51019);
  not i51022(x51022, x51021);
  not i51024(x51024, x51023);
  not i51026(x51026, x51025);
  not i51028(x51028, x51027);
  not i51030(x51030, x51029);
  not i51032(x51032, x51031);
  not i51034(x51034, x51033);
  not i51036(x51036, x51035);
  not i51038(x51038, x51037);
  not i51040(x51040, x51039);
  not i51042(x51042, x51041);
  not i51045(x51045, x51044);
  not i51047(x51047, x51046);
  not i51049(x51049, x51048);
  not i51051(x51051, x51050);
  not i51053(x51053, x51052);
  not i51055(x51055, x51054);
  not i51057(x51057, x51056);
  not i51059(x51059, x51058);
  not i51061(x51061, x51060);
  not i51063(x51063, x51062);
  not i51065(x51065, x51064);
  not i51067(x51067, x51066);
  not i51069(x51069, x51068);
  not i51071(x51071, x51070);
  not i51073(x51073, x51072);
  not i51075(x51075, x51074);
  not i51077(x51077, x51076);
  not i51079(x51079, x51078);
  not i51081(x51081, x51080);
  not i51083(x51083, x51082);
  not i51085(x51085, x51084);
  not i51087(x51087, x51086);
  not i51089(x51089, x51088);
  not i51091(x51091, x51090);
  not i51093(x51093, x51092);
  not i51095(x51095, x51094);
  not i51097(x51097, x51096);
  not i51099(x51099, x51098);
  not i51101(x51101, x51100);
  not i51103(x51103, x51102);
  not i51105(x51105, x51104);
  not i51107(x51107, x51106);
  not i51109(x51109, x51108);
  not i51111(x51111, x51110);
  not i51113(x51113, x51112);
  not i51116(x51116, x51115);
  not i51118(x51118, x51117);
  not i51120(x51120, x51119);
  not i51122(x51122, x51121);
  not i51124(x51124, x51123);
  not i51126(x51126, x51125);
  not i51128(x51128, x51127);
  not i51130(x51130, x51129);
  not i51132(x51132, x51131);
  not i51134(x51134, x51133);
  not i51136(x51136, x51135);
  not i51138(x51138, x51137);
  not i51140(x51140, x51139);
  not i51142(x51142, x51141);
  not i51144(x51144, x51143);
  not i51146(x51146, x51145);
  not i51148(x51148, x51147);
  not i51150(x51150, x51149);
  not i51152(x51152, x51151);
  not i51154(x51154, x51153);
  not i51156(x51156, x51155);
  not i51158(x51158, x51157);
  not i51160(x51160, x51159);
  not i51162(x51162, x51161);
  not i51164(x51164, x51163);
  not i51166(x51166, x51165);
  not i51168(x51168, x51167);
  not i51170(x51170, x51169);
  not i51172(x51172, x51171);
  not i51174(x51174, x51173);
  not i51176(x51176, x51175);
  not i51178(x51178, x51177);
  not i51180(x51180, x51179);
  not i51182(x51182, x51181);
  not i51184(x51184, x51183);
  not i51186(x51186, x51185);
  not i51188(x51188, x51187);
  not i51190(x51190, x51189);
  not i51192(x51192, x51191);
  not i51194(x51194, x51193);
  not i51196(x51196, x51195);
  not i51198(x51198, x51197);
  not i51200(x51200, x51199);
  not i51202(x51202, x51201);
  not i51205(x51205, x51204);
  not i51207(x51207, x51206);
  not i51209(x51209, x51208);
  not i51211(x51211, x51210);
  not i51213(x51213, x51212);
  not i51215(x51215, x51214);
  not i51217(x51217, x51216);
  not i51219(x51219, x51218);
  not i51221(x51221, x51220);
  not i51223(x51223, x51222);
  not i51225(x51225, x51224);
  not i51227(x51227, x51226);
  not i51229(x51229, x51228);
  not i51231(x51231, x51230);
  not i51233(x51233, x51232);
  not i51235(x51235, x51234);
  not i51237(x51237, x51236);
  not i51239(x51239, x51238);
  not i51241(x51241, x51240);
  not i51243(x51243, x51242);
  not i51245(x51245, x51244);
  not i51247(x51247, x51246);
  not i51249(x51249, x51248);
  not i51251(x51251, x51250);
  not i51253(x51253, x51252);
  not i51255(x51255, x51254);
  not i51257(x51257, x51256);
  not i51259(x51259, x51258);
  not i51261(x51261, x51260);
  not i51263(x51263, x51262);
  not i51265(x51265, x51264);
  not i51267(x51267, x51266);
  not i51269(x51269, x51268);
  not i51271(x51271, x51270);
  not i51273(x51273, x51272);
  not i51275(x51275, x51274);
  not i51277(x51277, x51276);
  not i51279(x51279, x51278);
  not i51281(x51281, x51280);
  not i51283(x51283, x51282);
  not i51285(x51285, x51284);
  not i51287(x51287, x51286);
  not i51289(x51289, x51288);
  not i51291(x51291, x51290);
  not i51293(x51293, x51292);
  not i51295(x51295, x51294);
  not i51297(x51297, x51296);
  not i51299(x51299, x51298);
  not i51301(x51301, x51300);
  not i51303(x51303, x51302);
  not i51305(x51305, x51304);
  not i51307(x51307, x51306);
  not i51309(x51309, x51308);
  not i51312(x51312, x51311);
  not i51314(x51314, x51313);
  not i51316(x51316, x51315);
  not i51318(x51318, x51317);
  not i51320(x51320, x51319);
  not i51322(x51322, x51321);
  not i51324(x51324, x51323);
  not i51326(x51326, x51325);
  not i51328(x51328, x51327);
  not i51330(x51330, x51329);
  not i51332(x51332, x51331);
  not i51334(x51334, x51333);
  not i51336(x51336, x51335);
  not i51338(x51338, x51337);
  not i51340(x51340, x51339);
  not i51342(x51342, x51341);
  not i51344(x51344, x51343);
  not i51346(x51346, x51345);
  not i51348(x51348, x51347);
  not i51350(x51350, x51349);
  not i51352(x51352, x51351);
  not i51354(x51354, x51353);
  not i51356(x51356, x51355);
  not i51358(x51358, x51357);
  not i51360(x51360, x51359);
  not i51362(x51362, x51361);
  not i51364(x51364, x51363);
  not i51366(x51366, x51365);
  not i51368(x51368, x51367);
  not i51370(x51370, x51369);
  not i51372(x51372, x51371);
  not i51374(x51374, x51373);
  not i51376(x51376, x51375);
  not i51378(x51378, x51377);
  not i51380(x51380, x51379);
  not i51382(x51382, x51381);
  not i51384(x51384, x51383);
  not i51386(x51386, x51385);
  not i51388(x51388, x51387);
  not i51390(x51390, x51389);
  not i51392(x51392, x51391);
  not i51394(x51394, x51393);
  not i51396(x51396, x51395);
  not i51398(x51398, x51397);
  not i51400(x51400, x51399);
  not i51402(x51402, x51401);
  not i51404(x51404, x51403);
  not i51406(x51406, x51405);
  not i51408(x51408, x51407);
  not i51410(x51410, x51409);
  not i51412(x51412, x51411);
  not i51414(x51414, x51413);
  not i51416(x51416, x51415);
  not i51418(x51418, x51417);
  not i51420(x51420, x51419);
  not i51422(x51422, x51421);
  not i51424(x51424, x51423);
  not i51426(x51426, x51425);
  not i51428(x51428, x51427);
  not i51430(x51430, x51429);
  not i51432(x51432, x51431);
  not i51434(x51434, x51433);
  not i51437(x51437, x51436);
  not i51439(x51439, x51438);
  not i51441(x51441, x51440);
  not i51443(x51443, x51442);
  not i51445(x51445, x51444);
  not i51447(x51447, x51446);
  not i51449(x51449, x51448);
  not i51451(x51451, x51450);
  not i51453(x51453, x51452);
  not i51455(x51455, x51454);
  not i51457(x51457, x51456);
  not i51459(x51459, x51458);
  not i51461(x51461, x51460);
  not i51463(x51463, x51462);
  not i51465(x51465, x51464);
  not i51467(x51467, x51466);
  not i51469(x51469, x51468);
  not i51471(x51471, x51470);
  not i51473(x51473, x51472);
  not i51475(x51475, x51474);
  not i51477(x51477, x51476);
  not i51479(x51479, x51478);
  not i51481(x51481, x51480);
  not i51483(x51483, x51482);
  not i51485(x51485, x51484);
  not i51487(x51487, x51486);
  not i51489(x51489, x51488);
  not i51491(x51491, x51490);
  not i51493(x51493, x51492);
  not i51495(x51495, x51494);
  not i51497(x51497, x51496);
  not i51499(x51499, x51498);
  not i51501(x51501, x51500);
  not i51503(x51503, x51502);
  not i51505(x51505, x51504);
  not i51507(x51507, x51506);
  not i51509(x51509, x51508);
  not i51511(x51511, x51510);
  not i51513(x51513, x51512);
  not i51515(x51515, x51514);
  not i51517(x51517, x51516);
  not i51519(x51519, x51518);
  not i51521(x51521, x51520);
  not i51523(x51523, x51522);
  not i51525(x51525, x51524);
  not i51527(x51527, x51526);
  not i51529(x51529, x51528);
  not i51531(x51531, x51530);
  not i51533(x51533, x51532);
  not i51535(x51535, x51534);
  not i51537(x51537, x51536);
  not i51539(x51539, x51538);
  not i51541(x51541, x51540);
  not i51543(x51543, x51542);
  not i51545(x51545, x51544);
  not i51547(x51547, x51546);
  not i51549(x51549, x51548);
  not i51551(x51551, x51550);
  not i51553(x51553, x51552);
  not i51555(x51555, x51554);
  not i51557(x51557, x51556);
  not i51559(x51559, x51558);
  not i51561(x51561, x51560);
  not i51563(x51563, x51562);
  not i51565(x51565, x51564);
  not i51567(x51567, x51566);
  not i51569(x51569, x51568);
  not i51571(x51571, x51570);
  not i51573(x51573, x51572);
  not i51575(x51575, x51574);
  not i51577(x51577, x51576);
  not i51580(x51580, x51579);
  not i51582(x51582, x51581);
  not i51584(x51584, x51583);
  not i51586(x51586, x51585);
  not i51588(x51588, x51587);
  not i51590(x51590, x51589);
  not i51592(x51592, x51591);
  not i51594(x51594, x51593);
  not i51596(x51596, x51595);
  not i51598(x51598, x51597);
  not i51600(x51600, x51599);
  not i51602(x51602, x51601);
  not i51604(x51604, x51603);
  not i51606(x51606, x51605);
  not i51608(x51608, x51607);
  not i51610(x51610, x51609);
  not i51612(x51612, x51611);
  not i51614(x51614, x51613);
  not i51616(x51616, x51615);
  not i51618(x51618, x51617);
  not i51620(x51620, x51619);
  not i51622(x51622, x51621);
  not i51624(x51624, x51623);
  not i51626(x51626, x51625);
  not i51628(x51628, x51627);
  not i51630(x51630, x51629);
  not i51632(x51632, x51631);
  not i51634(x51634, x51633);
  not i51636(x51636, x51635);
  not i51638(x51638, x51637);
  not i51640(x51640, x51639);
  not i51642(x51642, x51641);
  not i51644(x51644, x51643);
  not i51646(x51646, x51645);
  not i51648(x51648, x51647);
  not i51650(x51650, x51649);
  not i51652(x51652, x51651);
  not i51654(x51654, x51653);
  not i51656(x51656, x51655);
  not i51658(x51658, x51657);
  not i51660(x51660, x51659);
  not i51662(x51662, x51661);
  not i51664(x51664, x51663);
  not i51666(x51666, x51665);
  not i51668(x51668, x51667);
  not i51670(x51670, x51669);
  not i51672(x51672, x51671);
  not i51674(x51674, x51673);
  not i51676(x51676, x51675);
  not i51678(x51678, x51677);
  not i51680(x51680, x51679);
  not i51682(x51682, x51681);
  not i51684(x51684, x51683);
  not i51686(x51686, x51685);
  not i51688(x51688, x51687);
  not i51690(x51690, x51689);
  not i51692(x51692, x51691);
  not i51694(x51694, x51693);
  not i51696(x51696, x51695);
  not i51698(x51698, x51697);
  not i51700(x51700, x51699);
  not i51702(x51702, x51701);
  not i51704(x51704, x51703);
  not i51706(x51706, x51705);
  not i51708(x51708, x51707);
  not i51710(x51710, x51709);
  not i51712(x51712, x51711);
  not i51714(x51714, x51713);
  not i51716(x51716, x51715);
  not i51718(x51718, x51717);
  not i51720(x51720, x51719);
  not i51722(x51722, x51721);
  not i51724(x51724, x51723);
  not i51726(x51726, x51725);
  not i51728(x51728, x51727);
  not i51730(x51730, x51729);
  not i51732(x51732, x51731);
  not i51734(x51734, x51733);
  not i51736(x51736, x51735);
  not i51738(x51738, x51737);
  not i51741(x51741, x51740);
  not i51743(x51743, x51742);
  not i51745(x51745, x51744);
  not i51747(x51747, x51746);
  not i51749(x51749, x51748);
  not i51751(x51751, x51750);
  not i51753(x51753, x51752);
  not i51755(x51755, x51754);
  not i51757(x51757, x51756);
  not i51759(x51759, x51758);
  not i51761(x51761, x51760);
  not i51763(x51763, x51762);
  not i51765(x51765, x51764);
  not i51767(x51767, x51766);
  not i51769(x51769, x51768);
  not i51771(x51771, x51770);
  not i51773(x51773, x51772);
  not i51775(x51775, x51774);
  not i51777(x51777, x51776);
  not i51779(x51779, x51778);
  not i51781(x51781, x51780);
  not i51783(x51783, x51782);
  not i51785(x51785, x51784);
  not i51787(x51787, x51786);
  not i51789(x51789, x51788);
  not i51791(x51791, x51790);
  not i51793(x51793, x51792);
  not i51795(x51795, x51794);
  not i51797(x51797, x51796);
  not i51799(x51799, x51798);
  not i51801(x51801, x51800);
  not i51803(x51803, x51802);
  not i51805(x51805, x51804);
  not i51807(x51807, x51806);
  not i51809(x51809, x51808);
  not i51811(x51811, x51810);
  not i51813(x51813, x51812);
  not i51815(x51815, x51814);
  not i51817(x51817, x51816);
  not i51819(x51819, x51818);
  not i51821(x51821, x51820);
  not i51823(x51823, x51822);
  not i51825(x51825, x51824);
  not i51827(x51827, x51826);
  not i51829(x51829, x51828);
  not i51831(x51831, x51830);
  not i51833(x51833, x51832);
  not i51835(x51835, x51834);
  not i51837(x51837, x51836);
  not i51839(x51839, x51838);
  not i51841(x51841, x51840);
  not i51843(x51843, x51842);
  not i51845(x51845, x51844);
  not i51847(x51847, x51846);
  not i51849(x51849, x51848);
  not i51851(x51851, x51850);
  not i51853(x51853, x51852);
  not i51855(x51855, x51854);
  not i51857(x51857, x51856);
  not i51859(x51859, x51858);
  not i51861(x51861, x51860);
  not i51863(x51863, x51862);
  not i51865(x51865, x51864);
  not i51867(x51867, x51866);
  not i51869(x51869, x51868);
  not i51871(x51871, x51870);
  not i51873(x51873, x51872);
  not i51875(x51875, x51874);
  not i51877(x51877, x51876);
  not i51879(x51879, x51878);
  not i51881(x51881, x51880);
  not i51883(x51883, x51882);
  not i51885(x51885, x51884);
  not i51887(x51887, x51886);
  not i51889(x51889, x51888);
  not i51891(x51891, x51890);
  not i51893(x51893, x51892);
  not i51895(x51895, x51894);
  not i51897(x51897, x51896);
  not i51899(x51899, x51898);
  not i51901(x51901, x51900);
  not i51903(x51903, x51902);
  not i51905(x51905, x51904);
  not i51907(x51907, x51906);
  not i51909(x51909, x51908);
  not i51911(x51911, x51910);
  not i51913(x51913, x51912);
  not i51915(x51915, x51914);
  not i51917(x51917, x51916);
  not i51920(x51920, x51919);
  not i51922(x51922, x51921);
  not i51924(x51924, x51923);
  not i51926(x51926, x51925);
  not i51928(x51928, x51927);
  not i51930(x51930, x51929);
  not i51932(x51932, x51931);
  not i51934(x51934, x51933);
  not i51936(x51936, x51935);
  not i51938(x51938, x51937);
  not i51940(x51940, x51939);
  not i51942(x51942, x51941);
  not i51944(x51944, x51943);
  not i51946(x51946, x51945);
  not i51948(x51948, x51947);
  not i51950(x51950, x51949);
  not i51952(x51952, x51951);
  not i51954(x51954, x51953);
  not i51956(x51956, x51955);
  not i51958(x51958, x51957);
  not i51960(x51960, x51959);
  not i51962(x51962, x51961);
  not i51964(x51964, x51963);
  not i51966(x51966, x51965);
  not i51968(x51968, x51967);
  not i51970(x51970, x51969);
  not i51972(x51972, x51971);
  not i51974(x51974, x51973);
  not i51976(x51976, x51975);
  not i51978(x51978, x51977);
  not i51980(x51980, x51979);
  not i51982(x51982, x51981);
  not i51989(x51989, x51988);
  not i51997(x51997, x51996);
  not i52005(x52005, x52004);
  not i52016(x52016, x52015);
  not i52024(x52024, x52023);
  not i52032(x52032, x52031);
  not i52040(x52040, x52039);
  not i52044(x52044, x52043);
  not i52049(x52049, x52048);
  not i52057(x52057, x52056);
  not i52061(x52061, x52060);
  not i52069(x52069, x52068);
  not i52077(x52077, x52076);
  not i52081(x52081, x52080);
  not i52086(x52086, x52085);
  not i52090(x52090, x52089);
  not i52095(x52095, x52094);
  not i52103(x52103, x52102);
  not i52107(x52107, x52106);
  not i52112(x52112, x52111);
  not i52116(x52116, x52115);
  not i52121(x52121, x52120);
  not i52129(x52129, x52128);
  not i52133(x52133, x52132);
  not i52138(x52138, x52137);
  not i52142(x52142, x52141);
  not i52150(x52150, x52149);
  not i52158(x52158, x52157);
  not i52162(x52162, x52161);
  not i52167(x52167, x52166);
  not i52171(x52171, x52170);
  not i52176(x52176, x52175);
  not i52180(x52180, x52179);
  not i52185(x52185, x52184);
  not i52193(x52193, x52192);
  not i52197(x52197, x52196);
  not i52202(x52202, x52201);
  not i52206(x52206, x52205);
  not i52211(x52211, x52210);
  not i52215(x52215, x52214);
  not i52220(x52220, x52219);
  not i52228(x52228, x52227);
  not i52232(x52232, x52231);
  not i52237(x52237, x52236);
  not i52241(x52241, x52240);
  not i52246(x52246, x52245);
  not i52250(x52250, x52249);
  not i52258(x52258, x52257);
  not i52266(x52266, x52265);
  not i52270(x52270, x52269);
  not i52275(x52275, x52274);
  not i52279(x52279, x52278);
  not i52284(x52284, x52283);
  not i52288(x52288, x52287);
  not i52293(x52293, x52292);
  not i52301(x52301, x52300);
  not i52309(x52309, x52308);
  not i52313(x52313, x52312);
  not i52318(x52318, x52317);
  not i52322(x52322, x52321);
  not i52327(x52327, x52326);
  not i52331(x52331, x52330);
  not i52336(x52336, x52335);
  not i52340(x52340, x52339);
  not i52345(x52345, x52344);
  not i52353(x52353, x52352);
  not i52357(x52357, x52356);
  not i52362(x52362, x52361);
  not i52366(x52366, x52365);
  not i52371(x52371, x52370);
  not i52375(x52375, x52374);
  not i52380(x52380, x52379);
  not i52384(x52384, x52383);
  not i52392(x52392, x52391);
  not i52400(x52400, x52399);
  not i52404(x52404, x52403);
  not i52409(x52409, x52408);
  not i52413(x52413, x52412);
  not i52418(x52418, x52417);
  not i52422(x52422, x52421);
  not i52427(x52427, x52426);
  not i52431(x52431, x52430);
  not i52436(x52436, x52435);
  not i52440(x52440, x52439);
  not i52445(x52445, x52444);
  not i52453(x52453, x52452);
  not i52457(x52457, x52456);
  not i52462(x52462, x52461);
  not i52466(x52466, x52465);
  not i52471(x52471, x52470);
  not i52475(x52475, x52474);
  not i52480(x52480, x52479);
  not i52484(x52484, x52483);
  not i52489(x52489, x52488);
  not i52493(x52493, x52492);
  not i52498(x52498, x52497);
  not i52506(x52506, x52505);
  not i52510(x52510, x52509);
  not i52515(x52515, x52514);
  not i52519(x52519, x52518);
  not i52524(x52524, x52523);
  not i52528(x52528, x52527);
  not i52533(x52533, x52532);
  not i52537(x52537, x52536);
  not i52542(x52542, x52541);
  not i52546(x52546, x52545);
  not i52554(x52554, x52553);
  not i52562(x52562, x52561);
  not i52566(x52566, x52565);
  not i52571(x52571, x52570);
  not i52575(x52575, x52574);
  not i52580(x52580, x52579);
  not i52584(x52584, x52583);
  not i52589(x52589, x52588);
  not i52593(x52593, x52592);
  not i52598(x52598, x52597);
  not i52602(x52602, x52601);
  not i52607(x52607, x52606);
  not i52611(x52611, x52610);
  not i52616(x52616, x52615);
  not i52624(x52624, x52623);
  not i52628(x52628, x52627);
  not i52633(x52633, x52632);
  not i52637(x52637, x52636);
  not i52642(x52642, x52641);
  not i52646(x52646, x52645);
  not i52651(x52651, x52650);
  not i52655(x52655, x52654);
  not i52660(x52660, x52659);
  not i52664(x52664, x52663);
  not i52669(x52669, x52668);
  not i52673(x52673, x52672);
  not i52678(x52678, x52677);
  not i52686(x52686, x52685);
  not i52690(x52690, x52689);
  not i52695(x52695, x52694);
  not i52699(x52699, x52698);
  not i52704(x52704, x52703);
  not i52708(x52708, x52707);
  not i52713(x52713, x52712);
  not i52717(x52717, x52716);
  not i52722(x52722, x52721);
  not i52726(x52726, x52725);
  not i52731(x52731, x52730);
  not i52735(x52735, x52734);
  not i52743(x52743, x52742);
  not i52751(x52751, x52750);
  not i52755(x52755, x52754);
  not i52760(x52760, x52759);
  not i52764(x52764, x52763);
  not i52769(x52769, x52768);
  not i52773(x52773, x52772);
  not i52778(x52778, x52777);
  not i52782(x52782, x52781);
  not i52787(x52787, x52786);
  not i52791(x52791, x52790);
  not i52796(x52796, x52795);
  not i52800(x52800, x52799);
  not i52805(x52805, x52804);
  not i52813(x52813, x52812);
  not i52821(x52821, x52820);
  not i52825(x52825, x52824);
  not i52830(x52830, x52829);
  not i52834(x52834, x52833);
  not i52839(x52839, x52838);
  not i52843(x52843, x52842);
  not i52848(x52848, x52847);
  not i52852(x52852, x52851);
  not i52857(x52857, x52856);
  not i52861(x52861, x52860);
  not i52866(x52866, x52865);
  not i52870(x52870, x52869);
  not i52875(x52875, x52874);
  not i52879(x52879, x52878);
  not i52884(x52884, x52883);
  not i52892(x52892, x52891);
  not i52896(x52896, x52895);
  not i52901(x52901, x52900);
  not i52905(x52905, x52904);
  not i52910(x52910, x52909);
  not i52914(x52914, x52913);
  not i52919(x52919, x52918);
  not i52923(x52923, x52922);
  not i52928(x52928, x52927);
  not i52932(x52932, x52931);
  not i52937(x52937, x52936);
  not i52941(x52941, x52940);
  not i52946(x52946, x52945);
  not i52950(x52950, x52949);
  not i52958(x52958, x52957);
  not i52966(x52966, x52965);
  not i52970(x52970, x52969);
  not i52975(x52975, x52974);
  not i52979(x52979, x52978);
  not i52984(x52984, x52983);
  not i52988(x52988, x52987);
  not i52993(x52993, x52992);
  not i52997(x52997, x52996);
  not i53002(x53002, x53001);
  not i53006(x53006, x53005);
  not i53011(x53011, x53010);
  not i53015(x53015, x53014);
  not i53020(x53020, x53019);
  not i53024(x53024, x53023);
  not i53029(x53029, x53028);
  not i53033(x53033, x53032);
  not i53038(x53038, x53037);
  not i53046(x53046, x53045);
  not i53050(x53050, x53049);
  not i53055(x53055, x53054);
  not i53059(x53059, x53058);
  not i53064(x53064, x53063);
  not i53068(x53068, x53067);
  not i53073(x53073, x53072);
  not i53077(x53077, x53076);
  not i53082(x53082, x53081);
  not i53086(x53086, x53085);
  not i53091(x53091, x53090);
  not i53095(x53095, x53094);
  not i53100(x53100, x53099);
  not i53104(x53104, x53103);
  not i53109(x53109, x53108);
  not i53113(x53113, x53112);
  not i53118(x53118, x53117);
  not i53126(x53126, x53125);
  not i53130(x53130, x53129);
  not i53135(x53135, x53134);
  not i53139(x53139, x53138);
  not i53144(x53144, x53143);
  not i53148(x53148, x53147);
  not i53153(x53153, x53152);
  not i53157(x53157, x53156);
  not i53162(x53162, x53161);
  not i53166(x53166, x53165);
  not i53171(x53171, x53170);
  not i53175(x53175, x53174);
  not i53180(x53180, x53179);
  not i53184(x53184, x53183);
  not i53189(x53189, x53188);
  not i53193(x53193, x53192);
  not i53201(x53201, x53200);
  not i53205(x53205, x53204);
  not i53210(x53210, x53209);
  not i53214(x53214, x53213);
  not i53219(x53219, x53218);
  not i53223(x53223, x53222);
  not i53228(x53228, x53227);
  not i53232(x53232, x53231);
  not i53237(x53237, x53236);
  not i53241(x53241, x53240);
  not i53246(x53246, x53245);
  not i53250(x53250, x53249);
  not i53255(x53255, x53254);
  not i53259(x53259, x53258);
  not i53264(x53264, x53263);
  not i53268(x53268, x53267);
  not i53273(x53273, x53272);
  not i53277(x53277, x53276);
  not i53282(x53282, x53281);
  not i53286(x53286, x53285);
  not i53291(x53291, x53290);
  not i53295(x53295, x53294);
  not i53300(x53300, x53299);
  not i53304(x53304, x53303);
  not i53309(x53309, x53308);
  not i53313(x53313, x53312);
  not i53318(x53318, x53317);
  not i53322(x53322, x53321);
  not i53327(x53327, x53326);
  not i53331(x53331, x53330);
  not i53336(x53336, x53335);
  not i53340(x53340, x53339);
  not i53345(x53345, x53344);
  not i53349(x53349, x53348);
  not i53354(x53354, x53353);
  not i53358(x53358, x53357);
  not i53363(x53363, x53362);
  not i53367(x53367, x53366);
  not i53372(x53372, x53371);
  not i53376(x53376, x53375);
  not i53381(x53381, x53380);
  not i53385(x53385, x53384);
  not i53389(x53389, x53388);
  not i53393(x53393, x53392);
  not i53397(x53397, x53396);
  not i53401(x53401, x53400);
  not i53405(x53405, x53404);
  not i53409(x53409, x53408);
  not i53413(x53413, x53412);
  not i53417(x53417, x53416);
  not i53421(x53421, x53420);
  not i53425(x53425, x53424);
  not i53429(x53429, x53428);
  not i53433(x53433, x53432);
  not i53437(x53437, x53436);
  not i53441(x53441, x53440);
  not i53445(x53445, x53444);
  not i53449(x53449, x53448);
  not i53453(x53453, x53452);
  not i53457(x53457, x53456);
  not i53461(x53461, x53460);
  not i53462(x53462, x51993);
  not i53463(x53463, x52001);
  not i53465(x53465, x52009);
  not i53469(x53469, x52028);
  not i53470(x53470, x52020);
  not i53477(x53477, x52045);
  not i53478(x53478, x52036);
  not i53485(x53485, x52062);
  not i53486(x53486, x52053);
  not i53489(x53489, x53488);
  not i53498(x53498, x52082);
  not i53499(x53499, x52073);
  not i53502(x53502, x53501);
  not i53504(x53504, x52091);
  not i53511(x53511, x53510);
  not i53515(x53515, x53514);
  not i53518(x53518, x52108);
  not i53519(x53519, x52099);
  not i53522(x53522, x53521);
  not i53524(x53524, x52117);
  not i53531(x53531, x53530);
  not i53535(x53535, x53534);
  not i53538(x53538, x52134);
  not i53539(x53539, x52125);
  not i53542(x53542, x53541);
  not i53544(x53544, x52143);
  not i53551(x53551, x53550);
  not i53555(x53555, x53554);
  not i53558(x53558, x52163);
  not i53559(x53559, x52154);
  not i53562(x53562, x53561);
  not i53564(x53564, x52172);
  not i53568(x53568, x52181);
  not i53572(x53572, x53571);
  not i53576(x53576, x53575);
  not i53579(x53579, x52198);
  not i53580(x53580, x52189);
  not i53583(x53583, x53582);
  not i53585(x53585, x52207);
  not i53589(x53589, x52216);
  not i53593(x53593, x53592);
  not i53597(x53597, x53596);
  not i53600(x53600, x52233);
  not i53601(x53601, x52224);
  not i53604(x53604, x53603);
  not i53606(x53606, x52242);
  not i53611(x53611, x52251);
  not i53617(x53617, x53616);
  not i53621(x53621, x53620);
  not i53624(x53624, x52271);
  not i53625(x53625, x52262);
  not i53628(x53628, x53627);
  not i53630(x53630, x52280);
  not i53635(x53635, x52297);
  not i53636(x53636, x52289);
  not i53642(x53642, x53641);
  not i53646(x53646, x53645);
  not i53652(x53652, x52314);
  not i53653(x53653, x52305);
  not i53656(x53656, x53655);
  not i53658(x53658, x52323);
  not i53663(x53663, x52341);
  not i53664(x53664, x52332);
  not i53670(x53670, x53669);
  not i53674(x53674, x53673);
  not i53680(x53680, x52358);
  not i53681(x53681, x52349);
  not i53684(x53684, x53683);
  not i53686(x53686, x52367);
  not i53691(x53691, x52385);
  not i53692(x53692, x52376);
  not i53695(x53695, x53694);
  not i53699(x53699, x53698);
  not i53704(x53704, x53703);
  not i53708(x53708, x53707);
  not i53714(x53714, x52405);
  not i53715(x53715, x52396);
  not i53718(x53718, x53717);
  not i53720(x53720, x52414);
  not i53725(x53725, x52432);
  not i53726(x53726, x52423);
  not i53729(x53729, x53728);
  not i53731(x53731, x52441);
  not i53734(x53734, x53733);
  not i53739(x53739, x53738);
  not i53743(x53743, x53742);
  not i53748(x53748, x53747);
  not i53754(x53754, x52458);
  not i53755(x53755, x52449);
  not i53758(x53758, x53757);
  not i53760(x53760, x52467);
  not i53765(x53765, x52485);
  not i53766(x53766, x52476);
  not i53769(x53769, x53768);
  not i53771(x53771, x52494);
  not i53774(x53774, x53773);
  not i53779(x53779, x53778);
  not i53783(x53783, x53782);
  not i53788(x53788, x53787);
  not i53794(x53794, x52511);
  not i53795(x53795, x52502);
  not i53798(x53798, x53797);
  not i53800(x53800, x52520);
  not i53805(x53805, x52538);
  not i53806(x53806, x52529);
  not i53809(x53809, x53808);
  not i53811(x53811, x52547);
  not i53814(x53814, x53813);
  not i53819(x53819, x53818);
  not i53823(x53823, x53822);
  not i53828(x53828, x53827);
  not i53834(x53834, x52567);
  not i53835(x53835, x52558);
  not i53838(x53838, x53837);
  not i53840(x53840, x52576);
  not i53845(x53845, x52594);
  not i53846(x53846, x52585);
  not i53849(x53849, x53848);
  not i53851(x53851, x52603);
  not i53854(x53854, x53853);
  not i53856(x53856, x52612);
  not i53860(x53860, x53859);
  not i53864(x53864, x53863);
  not i53869(x53869, x53868);
  not i53873(x53873, x53872);
  not i53876(x53876, x52629);
  not i53877(x53877, x52620);
  not i53880(x53880, x53879);
  not i53882(x53882, x52638);
  not i53887(x53887, x52656);
  not i53888(x53888, x52647);
  not i53891(x53891, x53890);
  not i53893(x53893, x52665);
  not i53896(x53896, x53895);
  not i53898(x53898, x52674);
  not i53902(x53902, x53901);
  not i53906(x53906, x53905);
  not i53911(x53911, x53910);
  not i53915(x53915, x53914);
  not i53918(x53918, x52691);
  not i53919(x53919, x52682);
  not i53922(x53922, x53921);
  not i53924(x53924, x52700);
  not i53929(x53929, x52718);
  not i53930(x53930, x52709);
  not i53933(x53933, x53932);
  not i53935(x53935, x52727);
  not i53938(x53938, x53937);
  not i53941(x53941, x52736);
  not i53947(x53947, x53946);
  not i53951(x53951, x53950);
  not i53956(x53956, x53955);
  not i53960(x53960, x53959);
  not i53963(x53963, x52756);
  not i53964(x53964, x52747);
  not i53967(x53967, x53966);
  not i53969(x53969, x52765);
  not i53974(x53974, x52783);
  not i53975(x53975, x52774);
  not i53978(x53978, x53977);
  not i53980(x53980, x52792);
  not i53983(x53983, x53982);
  not i53986(x53986, x52809);
  not i53987(x53987, x52801);
  not i53993(x53993, x53992);
  not i53997(x53997, x53996);
  not i54002(x54002, x54001);
  not i54006(x54006, x54005);
  not i54012(x54012, x52826);
  not i54013(x54013, x52817);
  not i54016(x54016, x54015);
  not i54018(x54018, x52835);
  not i54021(x54021, x54020);
  not i54024(x54024, x52853);
  not i54025(x54025, x52844);
  not i54028(x54028, x54027);
  not i54030(x54030, x52862);
  not i54033(x54033, x54032);
  not i54036(x54036, x52880);
  not i54037(x54037, x52871);
  not i54043(x54043, x54042);
  not i54047(x54047, x54046);
  not i54052(x54052, x54051);
  not i54056(x54056, x54055);
  not i54062(x54062, x52897);
  not i54063(x54063, x52888);
  not i54066(x54066, x54065);
  not i54068(x54068, x52906);
  not i54071(x54071, x54070);
  not i54074(x54074, x52924);
  not i54075(x54075, x52915);
  not i54078(x54078, x54077);
  not i54080(x54080, x52933);
  not i54083(x54083, x54082);
  not i54086(x54086, x52951);
  not i54087(x54087, x52942);
  not i54090(x54090, x54089);
  not i54094(x54094, x54093);
  not i54099(x54099, x54098);
  not i54103(x54103, x54102);
  not i54108(x54108, x54107);
  not i54112(x54112, x54111);
  not i54118(x54118, x52971);
  not i54119(x54119, x52962);
  not i54122(x54122, x54121);
  not i54124(x54124, x52980);
  not i54127(x54127, x54126);
  not i54130(x54130, x52998);
  not i54131(x54131, x52989);
  not i54134(x54134, x54133);
  not i54136(x54136, x53007);
  not i54139(x54139, x54138);
  not i54142(x54142, x53025);
  not i54143(x54143, x53016);
  not i54146(x54146, x54145);
  not i54148(x54148, x53034);
  not i54151(x54151, x54150);
  not i54156(x54156, x54155);
  not i54160(x54160, x54159);
  not i54165(x54165, x54164);
  not i54169(x54169, x54168);
  not i54174(x54174, x54173);
  not i54178(x54178, x54177);
  not i54181(x54181, x53051);
  not i54182(x54182, x53042);
  not i54185(x54185, x54184);
  not i54187(x54187, x53060);
  not i54190(x54190, x54189);
  not i54193(x54193, x53078);
  not i54194(x54194, x53069);
  not i54197(x54197, x54196);
  not i54199(x54199, x53087);
  not i54202(x54202, x54201);
  not i54205(x54205, x53105);
  not i54206(x54206, x53096);
  not i54209(x54209, x54208);
  not i54211(x54211, x53114);
  not i54214(x54214, x54213);
  not i54219(x54219, x54218);
  not i54223(x54223, x54222);
  not i54228(x54228, x54227);
  not i54232(x54232, x54231);
  not i54237(x54237, x54236);
  not i54241(x54241, x54240);
  not i54244(x54244, x53131);
  not i54245(x54245, x53122);
  not i54248(x54248, x54247);
  not i54250(x54250, x53140);
  not i54253(x54253, x54252);
  not i54256(x54256, x53158);
  not i54257(x54257, x53149);
  not i54260(x54260, x54259);
  not i54262(x54262, x53167);
  not i54265(x54265, x54264);
  not i54268(x54268, x53185);
  not i54269(x54269, x53176);
  not i54272(x54272, x54271);
  not i54274(x54274, x53194);
  not i54277(x54277, x54276);
  not i54282(x54282, x54281);
  not i54286(x54286, x54285);
  not i54290(x54290, x54289);
  not i54295(x54295, x54294);
  not i54299(x54299, x54298);
  not i54304(x54304, x54303);
  not i54308(x54308, x54307);
  not i54311(x54311, x53215);
  not i54312(x54312, x53206);
  not i54315(x54315, x54314);
  not i54317(x54317, x53224);
  not i54320(x54320, x54319);
  not i54323(x54323, x53242);
  not i54324(x54324, x53233);
  not i54327(x54327, x54326);
  not i54329(x54329, x53251);
  not i54332(x54332, x54331);
  not i54335(x54335, x53269);
  not i54336(x54336, x53260);
  not i54339(x54339, x54338);
  not i54341(x54341, x53278);
  not i54344(x54344, x54343);
  not i54346(x54346, x53287);
  not i54350(x54350, x54349);
  not i54354(x54354, x54353);
  not i54358(x54358, x54357);
  not i54363(x54363, x54362);
  not i54367(x54367, x54366);
  not i54372(x54372, x54371);
  not i54376(x54376, x54375);
  not i54379(x54379, x53305);
  not i54380(x54380, x53296);
  not i54383(x54383, x54382);
  not i54385(x54385, x53314);
  not i54388(x54388, x54387);
  not i54390(x54390, x53332);
  not i54391(x54391, x53323);
  not i54394(x54394, x54393);
  not i54396(x54396, x53341);
  not i54399(x54399, x54398);
  not i54401(x54401, x53359);
  not i54402(x54402, x53350);
  not i54405(x54405, x54404);
  not i54407(x54407, x53368);
  not i54410(x54410, x54409);
  not i54411(x54411, x53377);
  not i54415(x54415, x54414);
  not i54419(x54419, x54418);
  not i54423(x54423, x54422);
  not i54427(x54427, x54426);
  not i54431(x54431, x54430);
  not i54435(x54435, x54434);
  not i54439(x54439, x54438);
  not i54443(x54443, x54442);
  not i54447(x54447, x54446);
  not i54451(x54451, x54450);
  not i54455(x54455, x54454);
  not i54459(x54459, x54458);
  not i54463(x54463, x54462);
  not i54464(x54464, x53493);
  not i54468(x54468, x54467);
  not i54469(x54469, x53507);
  not i54470(x54470, x53516);
  not i54474(x54474, x54473);
  not i54475(x54475, x53527);
  not i54476(x54476, x53536);
  not i54480(x54480, x54479);
  not i54484(x54484, x54483);
  not i54485(x54485, x53547);
  not i54486(x54486, x53556);
  not i54490(x54490, x54489);
  not i54494(x54494, x54493);
  not i54495(x54495, x53567);
  not i54496(x54496, x53577);
  not i54500(x54500, x54499);
  not i54504(x54504, x54503);
  not i54505(x54505, x53588);
  not i54506(x54506, x53598);
  not i54510(x54510, x54509);
  not i54514(x54514, x54513);
  not i54516(x54516, x53609);
  not i54519(x54519, x53622);
  not i54523(x54523, x54522);
  not i54527(x54527, x54526);
  not i54529(x54529, x53633);
  not i54532(x54532, x53647);
  not i54536(x54536, x54535);
  not i54540(x54540, x54539);
  not i54544(x54544, x54543);
  not i54546(x54546, x53661);
  not i54549(x54549, x53675);
  not i54553(x54553, x54552);
  not i54557(x54557, x54556);
  not i54561(x54561, x54560);
  not i54563(x54563, x53700);
  not i54564(x54564, x53689);
  not i54567(x54567, x53709);
  not i54571(x54571, x54570);
  not i54575(x54575, x54574);
  not i54579(x54579, x54578);
  not i54581(x54581, x53735);
  not i54582(x54582, x53723);
  not i54585(x54585, x53744);
  not i54587(x54587, x53752);
  not i54590(x54590, x54589);
  not i54594(x54594, x54593);
  not i54598(x54598, x54597);
  not i54600(x54600, x53775);
  not i54601(x54601, x53763);
  not i54604(x54604, x53784);
  not i54606(x54606, x53792);
  not i54609(x54609, x54608);
  not i54613(x54613, x54612);
  not i54617(x54617, x54616);
  not i54621(x54621, x54620);
  not i54624(x54624, x53815);
  not i54625(x54625, x53803);
  not i54628(x54628, x53824);
  not i54630(x54630, x53832);
  not i54633(x54633, x54632);
  not i54637(x54637, x54636);
  not i54641(x54641, x54640);
  not i54645(x54645, x54644);
  not i54651(x54651, x53855);
  not i54652(x54652, x53843);
  not i54655(x54655, x53865);
  not i54657(x54657, x53874);
  not i54660(x54660, x54659);
  not i54664(x54664, x54663);
  not i54668(x54668, x54667);
  not i54672(x54672, x54671);
  not i54678(x54678, x53897);
  not i54679(x54679, x53885);
  not i54682(x54682, x53907);
  not i54684(x54684, x53916);
  not i54687(x54687, x54686);
  not i54691(x54691, x54690);
  not i54695(x54695, x54694);
  not i54699(x54699, x54698);
  not i54705(x54705, x53939);
  not i54706(x54706, x53927);
  not i54709(x54709, x54708);
  not i54713(x54713, x54712);
  not i54715(x54715, x53952);
  not i54717(x54717, x53961);
  not i54720(x54720, x54719);
  not i54724(x54724, x54723);
  not i54728(x54728, x54727);
  not i54732(x54732, x54731);
  not i54738(x54738, x53984);
  not i54739(x54739, x53972);
  not i54742(x54742, x54741);
  not i54746(x54746, x54745);
  not i54748(x54748, x53998);
  not i54750(x54750, x54007);
  not i54753(x54753, x54752);
  not i54757(x54757, x54756);
  not i54761(x54761, x54760);
  not i54766(x54766, x54765);
  not i54770(x54770, x54769);
  not i54776(x54776, x54034);
  not i54777(x54777, x54022);
  not i54780(x54780, x54779);
  not i54784(x54784, x54783);
  not i54786(x54786, x54048);
  not i54788(x54788, x54057);
  not i54791(x54791, x54790);
  not i54795(x54795, x54794);
  not i54799(x54799, x54798);
  not i54804(x54804, x54803);
  not i54808(x54808, x54807);
  not i54814(x54814, x54084);
  not i54815(x54815, x54072);
  not i54818(x54818, x54817);
  not i54820(x54820, x54095);
  not i54823(x54823, x54822);
  not i54825(x54825, x54104);
  not i54827(x54827, x54113);
  not i54830(x54830, x54829);
  not i54834(x54834, x54833);
  not i54838(x54838, x54837);
  not i54843(x54843, x54842);
  not i54847(x54847, x54846);
  not i54853(x54853, x54140);
  not i54854(x54854, x54128);
  not i54857(x54857, x54856);
  not i54859(x54859, x54152);
  not i54862(x54862, x54861);
  not i54864(x54864, x54161);
  not i54866(x54866, x54170);
  not i54869(x54869, x54868);
  not i54871(x54871, x54179);
  not i54874(x54874, x54873);
  not i54878(x54878, x54877);
  not i54883(x54883, x54882);
  not i54887(x54887, x54886);
  not i54893(x54893, x54203);
  not i54894(x54894, x54191);
  not i54897(x54897, x54896);
  not i54899(x54899, x54215);
  not i54902(x54902, x54901);
  not i54904(x54904, x54224);
  not i54906(x54906, x54233);
  not i54909(x54909, x54908);
  not i54911(x54911, x54242);
  not i54914(x54914, x54913);
  not i54918(x54918, x54917);
  not i54923(x54923, x54922);
  not i54927(x54927, x54926);
  not i54933(x54933, x54266);
  not i54934(x54934, x54254);
  not i54937(x54937, x54936);
  not i54939(x54939, x54278);
  not i54942(x54942, x54941);
  not i54945(x54945, x54291);
  not i54948(x54948, x54947);
  not i54950(x54950, x54300);
  not i54953(x54953, x54952);
  not i54956(x54956, x54309);
  not i54959(x54959, x54958);
  not i54963(x54963, x54962);
  not i54968(x54968, x54967);
  not i54972(x54972, x54971);
  not i54977(x54977, x54976);
  not i54981(x54981, x54980);
  not i54984(x54984, x54333);
  not i54985(x54985, x54321);
  not i54988(x54988, x54987);
  not i54990(x54990, x54345);
  not i54993(x54993, x54992);
  not i54995(x54995, x54359);
  not i54998(x54998, x54997);
  not i55000(x55000, x54368);
  not i55003(x55003, x55002);
  not i55005(x55005, x54377);
  not i55008(x55008, x55007);
  not i55012(x55012, x55011);
  not i55016(x55016, x55015);
  not i55020(x55020, x55019);
  not i55024(x55024, x55023);
  not i55028(x55028, x55027);
  not i55038(x55038, x55037);
  not i55042(x55042, x55041);
  not i55049(x55049, x55048);
  not i55056(x55056, x55055);
  not i55060(x55060, x55059);
  not i55068(x55068, x55067);
  not i55072(x55072, x55071);
  not i55080(x55080, x55079);
  not i55084(x55084, x55083);
  not i55092(x55092, x55091);
  not i55096(x55096, x55095);
  not i55104(x55104, x55103);
  not i55108(x55108, x55107);
  not i55113(x55113, x55112);
  not i55117(x55117, x55116);
  not i55121(x55121, x55120);
  not i55126(x55126, x55125);
  not i55130(x55130, x55129);
  not i55134(x55134, x55133);
  not i55139(x55139, x55138);
  not i55143(x55143, x55142);
  not i55147(x55147, x55146);
  not i55152(x55152, x55151);
  not i55156(x55156, x55155);
  not i55160(x55160, x55159);
  not i55165(x55165, x55164);
  not i55169(x55169, x55168);
  not i55173(x55173, x55172);
  not i55177(x55177, x55176);
  not i55182(x55182, x55181);
  not i55186(x55186, x55185);
  not i55191(x55191, x55190);
  not i55195(x55195, x55194);
  not i55199(x55199, x55198);
  not i55204(x55204, x55203);
  not i55208(x55208, x55207);
  not i55213(x55213, x55212);
  not i55217(x55217, x55216);
  not i55221(x55221, x55220);
  not i55226(x55226, x55225);
  not i55230(x55230, x55229);
  not i55235(x55235, x55234);
  not i55239(x55239, x55238);
  not i55243(x55243, x55242);
  not i55248(x55248, x55247);
  not i55252(x55252, x55251);
  not i55257(x55257, x55256);
  not i55261(x55261, x55260);
  not i55265(x55265, x55264);
  not i55270(x55270, x55269);
  not i55274(x55274, x55273);
  not i55276(x55276, x54622);
  not i55280(x55280, x55279);
  not i55284(x55284, x55283);
  not i55288(x55288, x55287);
  not i55293(x55293, x55292);
  not i55297(x55297, x55296);
  not i55300(x55300, x54646);
  not i55303(x55303, x55302);
  not i55307(x55307, x55306);
  not i55312(x55312, x55311);
  not i55316(x55316, x55315);
  not i55321(x55321, x55320);
  not i55325(x55325, x55324);
  not i55328(x55328, x54673);
  not i55331(x55331, x55330);
  not i55335(x55335, x55334);
  not i55340(x55340, x55339);
  not i55344(x55344, x55343);
  not i55349(x55349, x55348);
  not i55353(x55353, x55352);
  not i55356(x55356, x54700);
  not i55359(x55359, x55358);
  not i55363(x55363, x55362);
  not i55368(x55368, x55367);
  not i55372(x55372, x55371);
  not i55375(x55375, x54714);
  not i55378(x55378, x55377);
  not i55382(x55382, x55381);
  not i55385(x55385, x54733);
  not i55388(x55388, x55387);
  not i55392(x55392, x55391);
  not i55397(x55397, x55396);
  not i55401(x55401, x55400);
  not i55404(x55404, x54747);
  not i55407(x55407, x55406);
  not i55409(x55409, x54762);
  not i55412(x55412, x55411);
  not i55415(x55415, x54771);
  not i55418(x55418, x55417);
  not i55422(x55422, x55421);
  not i55427(x55427, x55426);
  not i55431(x55431, x55430);
  not i55434(x55434, x54785);
  not i55437(x55437, x55436);
  not i55439(x55439, x54800);
  not i55442(x55442, x55441);
  not i55445(x55445, x54809);
  not i55448(x55448, x55447);
  not i55452(x55452, x55451);
  not i55457(x55457, x55456);
  not i55461(x55461, x55460);
  not i55464(x55464, x54824);
  not i55467(x55467, x55466);
  not i55469(x55469, x54839);
  not i55472(x55472, x55471);
  not i55475(x55475, x54848);
  not i55478(x55478, x55477);
  not i55482(x55482, x55481);
  not i55487(x55487, x55486);
  not i55491(x55491, x55490);
  not i55494(x55494, x54863);
  not i55497(x55497, x55496);
  not i55499(x55499, x54879);
  not i55502(x55502, x55501);
  not i55505(x55505, x54888);
  not i55508(x55508, x55507);
  not i55512(x55512, x55511);
  not i55517(x55517, x55516);
  not i55521(x55521, x55520);
  not i55524(x55524, x54903);
  not i55527(x55527, x55526);
  not i55529(x55529, x54919);
  not i55532(x55532, x55531);
  not i55535(x55535, x54928);
  not i55538(x55538, x55537);
  not i55542(x55542, x55541);
  not i55547(x55547, x55546);
  not i55551(x55551, x55550);
  not i55554(x55554, x54954);
  not i55555(x55555, x54943);
  not i55558(x55558, x55557);
  not i55560(x55560, x54964);
  not i55563(x55563, x55562);
  not i55565(x55565, x54982);
  not i55566(x55566, x54973);
  not i55569(x55569, x55568);
  not i55573(x55573, x55572);
  not i55577(x55577, x55576);
  not i55581(x55581, x55580);
  not i55594(x55594, x55593);
  not i55599(x55599, x55061);
  not i55602(x55602, x55601);
  not i55607(x55607, x55073);
  not i55610(x55610, x55609);
  not i55615(x55615, x55085);
  not i55618(x55618, x55617);
  not i55623(x55623, x55097);
  not i55626(x55626, x55625);
  not i55631(x55631, x55109);
  not i55634(x55634, x55633);
  not i55638(x55638, x55637);
  not i55642(x55642, x55641);
  not i55645(x55645, x55122);
  not i55648(x55648, x55647);
  not i55652(x55652, x55651);
  not i55656(x55656, x55655);
  not i55659(x55659, x55135);
  not i55662(x55662, x55661);
  not i55666(x55666, x55665);
  not i55670(x55670, x55669);
  not i55673(x55673, x55148);
  not i55676(x55676, x55675);
  not i55680(x55680, x55679);
  not i55684(x55684, x55683);
  not i55687(x55687, x55161);
  not i55690(x55690, x55689);
  not i55694(x55694, x55693);
  not i55698(x55698, x55697);
  not i55703(x55703, x55702);
  not i55705(x55705, x55178);
  not i55708(x55708, x55707);
  not i55713(x55713, x55712);
  not i55717(x55717, x55716);
  not i55720(x55720, x55187);
  not i55723(x55723, x55722);
  not i55725(x55725, x55200);
  not i55728(x55728, x55727);
  not i55733(x55733, x55732);
  not i55737(x55737, x55736);
  not i55740(x55740, x55209);
  not i55743(x55743, x55742);
  not i55745(x55745, x55222);
  not i55748(x55748, x55747);
  not i55753(x55753, x55752);
  not i55757(x55757, x55756);
  not i55760(x55760, x55231);
  not i55763(x55763, x55762);
  not i55765(x55765, x55244);
  not i55768(x55768, x55767);
  not i55773(x55773, x55772);
  not i55777(x55777, x55776);
  not i55780(x55780, x55253);
  not i55783(x55783, x55782);
  not i55785(x55785, x55266);
  not i55788(x55788, x55787);
  not i55793(x55793, x55792);
  not i55797(x55797, x55796);
  not i55800(x55800, x55275);
  not i55803(x55803, x55802);
  not i55805(x55805, x55289);
  not i55808(x55808, x55807);
  not i55813(x55813, x55812);
  not i55817(x55817, x55816);
  not i55820(x55820, x55308);
  not i55821(x55821, x55298);
  not i55824(x55824, x55823);
  not i55826(x55826, x55317);
  not i55829(x55829, x55828);
  not i55834(x55834, x55833);
  not i55838(x55838, x55837);
  not i55841(x55841, x55336);
  not i55842(x55842, x55326);
  not i55845(x55845, x55844);
  not i55847(x55847, x55345);
  not i55850(x55850, x55849);
  not i55855(x55855, x55854);
  not i55859(x55859, x55858);
  not i55862(x55862, x55364);
  not i55863(x55863, x55354);
  not i55866(x55866, x55865);
  not i55868(x55868, x55373);
  not i55871(x55871, x55870);
  not i55876(x55876, x55875);
  not i55880(x55880, x55879);
  not i55883(x55883, x55393);
  not i55884(x55884, x55383);
  not i55887(x55887, x55886);
  not i55889(x55889, x55402);
  not i55892(x55892, x55891);
  not i55897(x55897, x55896);
  not i55901(x55901, x55900);
  not i55904(x55904, x55423);
  not i55905(x55905, x55413);
  not i55908(x55908, x55907);
  not i55910(x55910, x55432);
  not i55913(x55913, x55912);
  not i55918(x55918, x55917);
  not i55922(x55922, x55921);
  not i55925(x55925, x55453);
  not i55926(x55926, x55443);
  not i55929(x55929, x55928);
  not i55931(x55931, x55462);
  not i55934(x55934, x55933);
  not i55939(x55939, x55938);
  not i55943(x55943, x55942);
  not i55946(x55946, x55483);
  not i55947(x55947, x55473);
  not i55950(x55950, x55949);
  not i55952(x55952, x55492);
  not i55955(x55955, x55954);
  not i55960(x55960, x55959);
  not i55964(x55964, x55963);
  not i55967(x55967, x55513);
  not i55968(x55968, x55503);
  not i55971(x55971, x55970);
  not i55973(x55973, x55522);
  not i55976(x55976, x55975);
  not i55981(x55981, x55980);
  not i55985(x55985, x55984);
  not i55988(x55988, x55543);
  not i55989(x55989, x55533);
  not i55992(x55992, x55991);
  not i55994(x55994, x55552);
  not i55997(x55997, x55996);
  not i56001(x56001, x56000);
  not i56005(x56005, x56004);
  not i56012(x56012, x56011);
  not i56016(x56016, x56015);
  not i56020(x56020, x56019);
  not i56024(x56024, x56023);
  not i56029(x56029, x56028);
  not i56033(x56033, x56032);
  not i56038(x56038, x56037);
  not i56042(x56042, x56041);
  not i56047(x56047, x56046);
  not i56051(x56051, x56050);
  not i56056(x56056, x56055);
  not i56060(x56060, x56059);
  not i56065(x56065, x56064);
  not i56066(x56066, x56062);
  not i56068(x56068, x55643);
  not i56071(x56071, x56070);
  not i56075(x56075, x56074);
  not i56080(x56080, x56079);
  not i56081(x56081, x56077);
  not i56083(x56083, x55657);
  not i56086(x56086, x56085);
  not i56090(x56090, x56089);
  not i56095(x56095, x56094);
  not i56096(x56096, x56092);
  not i56098(x56098, x55671);
  not i56101(x56101, x56100);
  not i56105(x56105, x56104);
  not i56110(x56110, x56109);
  not i56111(x56111, x56107);
  not i56113(x56113, x55685);
  not i56116(x56116, x56115);
  not i56120(x56120, x56119);
  not i56125(x56125, x56124);
  not i56126(x56126, x56122);
  not i56128(x56128, x55699);
  not i56131(x56131, x56130);
  not i56135(x56135, x56134);
  not i56140(x56140, x56139);
  not i56141(x56141, x56137);
  not i56143(x56143, x55718);
  not i56144(x56144, x55709);
  not i56147(x56147, x56146);
  not i56151(x56151, x56150);
  not i56156(x56156, x56155);
  not i56157(x56157, x56153);
  not i56159(x56159, x55738);
  not i56160(x56160, x55729);
  not i56163(x56163, x56162);
  not i56167(x56167, x56166);
  not i56172(x56172, x56171);
  not i56173(x56173, x56169);
  not i56175(x56175, x55758);
  not i56176(x56176, x55749);
  not i56179(x56179, x56178);
  not i56183(x56183, x56182);
  not i56188(x56188, x56187);
  not i56189(x56189, x56185);
  not i56191(x56191, x55778);
  not i56192(x56192, x55769);
  not i56195(x56195, x56194);
  not i56199(x56199, x56198);
  not i56204(x56204, x56203);
  not i56205(x56205, x56201);
  not i56207(x56207, x55798);
  not i56208(x56208, x55789);
  not i56211(x56211, x56210);
  not i56215(x56215, x56214);
  not i56220(x56220, x56219);
  not i56221(x56221, x56217);
  not i56223(x56223, x55818);
  not i56224(x56224, x55809);
  not i56227(x56227, x56226);
  not i56231(x56231, x56230);
  not i56236(x56236, x56235);
  not i56237(x56237, x56233);
  not i56239(x56239, x55839);
  not i56240(x56240, x55830);
  not i56243(x56243, x56242);
  not i56247(x56247, x56246);
  not i56252(x56252, x56251);
  not i56253(x56253, x56249);
  not i56255(x56255, x55860);
  not i56256(x56256, x55851);
  not i56259(x56259, x56258);
  not i56263(x56263, x56262);
  not i56268(x56268, x56267);
  not i56269(x56269, x56265);
  not i56271(x56271, x55881);
  not i56272(x56272, x55872);
  not i56275(x56275, x56274);
  not i56279(x56279, x56278);
  not i56284(x56284, x56283);
  not i56285(x56285, x56281);
  not i56287(x56287, x55902);
  not i56288(x56288, x55893);
  not i56291(x56291, x56290);
  not i56295(x56295, x56294);
  not i56300(x56300, x56299);
  not i56301(x56301, x56297);
  not i56303(x56303, x55923);
  not i56304(x56304, x55914);
  not i56307(x56307, x56306);
  not i56311(x56311, x56310);
  not i56316(x56316, x56315);
  not i56317(x56317, x56313);
  not i56319(x56319, x55944);
  not i56320(x56320, x55935);
  not i56323(x56323, x56322);
  not i56327(x56327, x56326);
  not i56332(x56332, x56331);
  not i56333(x56333, x56329);
  not i56335(x56335, x55965);
  not i56336(x56336, x55956);
  not i56339(x56339, x56338);
  not i56343(x56343, x56342);
  not i56348(x56348, x56347);
  not i56349(x56349, x56345);
  not i56351(x56351, x55986);
  not i56352(x56352, x55977);
  not i56355(x56355, x56354);
  not i56359(x56359, x56358);
  not i56363(x56363, x56362);
  not i56373(x56373, x56372);
  not i56377(x56377, x56376);
  not i56378(x56378, x56025);
  not i56382(x56382, x56381);
  not i56383(x56383, x56034);
  not i56387(x56387, x56386);
  not i56388(x56388, x56043);
  not i56392(x56392, x56391);
  not i56393(x56393, x56052);
  not i56397(x56397, x56396);
  not i56399(x56399, x56061);
  not i56402(x56402, x56401);
  not i56406(x56406, x56405);
  not i56409(x56409, x56076);
  not i56412(x56412, x56411);
  not i56416(x56416, x56415);
  not i56419(x56419, x56091);
  not i56422(x56422, x56421);
  not i56426(x56426, x56425);
  not i56429(x56429, x56106);
  not i56432(x56432, x56431);
  not i56436(x56436, x56435);
  not i56439(x56439, x56121);
  not i56442(x56442, x56441);
  not i56446(x56446, x56445);
  not i56449(x56449, x56136);
  not i56452(x56452, x56451);
  not i56456(x56456, x56455);
  not i56459(x56459, x56152);
  not i56462(x56462, x56461);
  not i56466(x56466, x56465);
  not i56469(x56469, x56168);
  not i56472(x56472, x56471);
  not i56476(x56476, x56475);
  not i56479(x56479, x56184);
  not i56482(x56482, x56481);
  not i56486(x56486, x56485);
  not i56489(x56489, x56200);
  not i56492(x56492, x56491);
  not i56496(x56496, x56495);
  not i56499(x56499, x56216);
  not i56502(x56502, x56501);
  not i56506(x56506, x56505);
  not i56509(x56509, x56232);
  not i56512(x56512, x56511);
  not i56516(x56516, x56515);
  not i56519(x56519, x56248);
  not i56522(x56522, x56521);
  not i56526(x56526, x56525);
  not i56529(x56529, x56264);
  not i56532(x56532, x56531);
  not i56536(x56536, x56535);
  not i56539(x56539, x56280);
  not i56542(x56542, x56541);
  not i56546(x56546, x56545);
  not i56549(x56549, x56296);
  not i56552(x56552, x56551);
  not i56556(x56556, x56555);
  not i56559(x56559, x56312);
  not i56562(x56562, x56561);
  not i56566(x56566, x56565);
  not i56569(x56569, x56328);
  not i56572(x56572, x56571);
  not i56576(x56576, x56575);
  not i56579(x56579, x56344);
  not i56582(x56582, x56581);
  not i56586(x56586, x56585);
  not i56590(x56590, x56589);
  not i56598(x56598, x56597);
  not i56602(x56602, x56601);
  not i56606(x56606, x56605);
  not i56610(x56610, x56609);
  not i56615(x56615, x56614);
  not i56619(x56619, x56618);
  not i56624(x56624, x56623);
  not i56628(x56628, x56627);
  not i56633(x56633, x56632);
  not i56637(x56637, x56636);
  not i56642(x56642, x56641);
  not i56646(x56646, x56645);
  not i56651(x56651, x56650);
  not i56655(x56655, x56654);
  not i56660(x56660, x56659);
  not i56664(x56664, x56663);
  not i56667(x56667, x56407);
  not i56670(x56670, x56669);
  not i56674(x56674, x56673);
  not i56677(x56677, x56417);
  not i56680(x56680, x56679);
  not i56684(x56684, x56683);
  not i56687(x56687, x56427);
  not i56690(x56690, x56689);
  not i56694(x56694, x56693);
  not i56697(x56697, x56437);
  not i56700(x56700, x56699);
  not i56704(x56704, x56703);
  not i56707(x56707, x56447);
  not i56710(x56710, x56709);
  not i56714(x56714, x56713);
  not i56717(x56717, x56457);
  not i56720(x56720, x56719);
  not i56724(x56724, x56723);
  not i56727(x56727, x56467);
  not i56730(x56730, x56729);
  not i56734(x56734, x56733);
  not i56737(x56737, x56477);
  not i56740(x56740, x56739);
  not i56744(x56744, x56743);
  not i56747(x56747, x56487);
  not i56750(x56750, x56749);
  not i56754(x56754, x56753);
  not i56757(x56757, x56497);
  not i56760(x56760, x56759);
  not i56764(x56764, x56763);
  not i56767(x56767, x56507);
  not i56770(x56770, x56769);
  not i56774(x56774, x56773);
  not i56777(x56777, x56517);
  not i56780(x56780, x56779);
  not i56784(x56784, x56783);
  not i56787(x56787, x56527);
  not i56790(x56790, x56789);
  not i56794(x56794, x56793);
  not i56797(x56797, x56537);
  not i56800(x56800, x56799);
  not i56804(x56804, x56803);
  not i56807(x56807, x56547);
  not i56810(x56810, x56809);
  not i56814(x56814, x56813);
  not i56817(x56817, x56557);
  not i56820(x56820, x56819);
  not i56824(x56824, x56823);
  not i56827(x56827, x56567);
  not i56830(x56830, x56829);
  not i56834(x56834, x56833);
  not i56837(x56837, x56577);
  not i56840(x56840, x56839);
  not i56844(x56844, x56843);
  not i56846(x56846, x56594);
  not i56852(x56852, x56851);
  not i56856(x56856, x56855);
  not i56858(x56858, x56611);
  not i56861(x56861, x56860);
  not i56863(x56863, x56620);
  not i56866(x56866, x56865);
  not i56868(x56868, x56629);
  not i56871(x56871, x56870);
  not i56873(x56873, x56638);
  not i56876(x56876, x56875);
  not i56878(x56878, x56647);
  not i56881(x56881, x56880);
  not i56883(x56883, x56656);
  not i56886(x56886, x56885);
  not i56888(x56888, x56665);
  not i56891(x56891, x56890);
  not i56893(x56893, x56675);
  not i56896(x56896, x56895);
  not i56898(x56898, x56685);
  not i56901(x56901, x56900);
  not i56903(x56903, x56695);
  not i56906(x56906, x56905);
  not i56908(x56908, x56705);
  not i56911(x56911, x56910);
  not i56913(x56913, x56715);
  not i56916(x56916, x56915);
  not i56918(x56918, x56725);
  not i56921(x56921, x56920);
  not i56923(x56923, x56735);
  not i56926(x56926, x56925);
  not i56928(x56928, x56745);
  not i56931(x56931, x56930);
  not i56933(x56933, x56755);
  not i56936(x56936, x56935);
  not i56938(x56938, x56765);
  not i56941(x56941, x56940);
  not i56943(x56943, x56775);
  not i56946(x56946, x56945);
  not i56948(x56948, x56785);
  not i56951(x56951, x56950);
  not i56953(x56953, x56795);
  not i56956(x56956, x56955);
  not i56958(x56958, x56805);
  not i56961(x56961, x56960);
  not i56963(x56963, x56815);
  not i56966(x56966, x56965);
  not i56968(x56968, x56825);
  not i56971(x56971, x56970);
  not i56973(x56973, x56835);
  not i56976(x56976, x56975);
  not i56977(x56977, x56845);
  not i56978(x56978, x56849);
  not i56979(x56979, x56853);
  not i56980(x56980, x56857);
  not i56981(x56981, x56862);
  not i56982(x56982, x56867);
  not i56983(x56983, x56872);
  not i56984(x56984, x56877);
  not i56985(x56985, x56882);
  not i56986(x56986, x56887);
  not i56987(x56987, x56892);
  not i56988(x56988, x56897);
  not i56989(x56989, x56902);
  not i56990(x56990, x56907);
  not i56991(x56991, x56912);
  not i56992(x56992, x56917);
  not i56993(x56993, x56922);
  not i56994(x56994, x56927);
  not i56995(x56995, x56932);
  not i56996(x56996, x56937);
  not i56997(x56997, x56942);
  not i56998(x56998, x56947);
  not i56999(x56999, x56952);
  not i57000(x57000, x56957);
  not i57001(x57001, x56962);
  not i57007(x57007, x57006);
  not i57011(x57011, x57010);
  not i57015(x57015, x57014);
  not i57019(x57019, x57018);
  not i57023(x57023, x57022);
  not i57027(x57027, x57026);
  not i57031(x57031, x57030);
  not i57035(x57035, x57034);
  not i57039(x57039, x57038);
  not i57043(x57043, x57042);
  not i57047(x57047, x57046);
  not i57051(x57051, x57050);
  not i57055(x57055, x57054);
  not i57059(x57059, x57058);
  not i57063(x57063, x57062);
  not i57067(x57067, x57066);
  not i57071(x57071, x57070);
  not i57075(x57075, x57074);
  not i57079(x57079, x57078);
  not i57083(x57083, x57082);
  not i57087(x57087, x57086);
  not i57091(x57091, x57090);
  not i57095(x57095, x57094);
  not i57099(x57099, x57098);
  not i57100(x57100, x57003);
  not i57102(x57102, x57005);
  not i57105(x57105, x57009);
  not i57108(x57108, x57013);
  not i57111(x57111, x57110);
  not i57113(x57113, x57017);
  not i57116(x57116, x57115);
  not i57118(x57118, x57021);
  not i57121(x57121, x57120);
  not i57123(x57123, x57025);
  not i57126(x57126, x57125);
  not i57128(x57128, x57029);
  not i57131(x57131, x57130);
  not i57133(x57133, x57033);
  not i57136(x57136, x57135);
  not i57138(x57138, x57037);
  not i57141(x57141, x57140);
  not i57143(x57143, x57041);
  not i57146(x57146, x57145);
  not i57148(x57148, x57045);
  not i57151(x57151, x57150);
  not i57153(x57153, x57049);
  not i57156(x57156, x57155);
  not i57158(x57158, x57053);
  not i57161(x57161, x57160);
  not i57163(x57163, x57057);
  not i57166(x57166, x57165);
  not i57168(x57168, x57061);
  not i57171(x57171, x57170);
  not i57173(x57173, x57065);
  not i57176(x57176, x57175);
  not i57178(x57178, x57069);
  not i57181(x57181, x57180);
  not i57183(x57183, x57073);
  not i57186(x57186, x57185);
  not i57188(x57188, x57077);
  not i57191(x57191, x57190);
  not i57193(x57193, x57081);
  not i57196(x57196, x57195);
  not i57198(x57198, x57085);
  not i57201(x57201, x57200);
  not i57203(x57203, x57089);
  not i57206(x57206, x57205);
  not i57208(x57208, x57093);
  not i57211(x57211, x57210);
  not i57213(x57213, x57097);
  not i57216(x57216, x57215);
  not i57217(x57217, x57103);
  not i57218(x57218, x57106);
  not i57220(x57220, x57109);
  not i57223(x57223, x57114);
  not i57226(x57226, x57119);
  not i57229(x57229, x57124);
  not i57232(x57232, x57129);
  not i57235(x57235, x57234);
  not i57237(x57237, x57134);
  not i57240(x57240, x57239);
  not i57242(x57242, x57139);
  not i57245(x57245, x57244);
  not i57247(x57247, x57144);
  not i57250(x57250, x57249);
  not i57252(x57252, x57149);
  not i57255(x57255, x57254);
  not i57257(x57257, x57154);
  not i57260(x57260, x57259);
  not i57262(x57262, x57159);
  not i57265(x57265, x57264);
  not i57267(x57267, x57164);
  not i57270(x57270, x57269);
  not i57272(x57272, x57169);
  not i57275(x57275, x57274);
  not i57277(x57277, x57174);
  not i57280(x57280, x57279);
  not i57282(x57282, x57179);
  not i57285(x57285, x57284);
  not i57287(x57287, x57184);
  not i57290(x57290, x57289);
  not i57292(x57292, x57189);
  not i57295(x57295, x57294);
  not i57297(x57297, x57194);
  not i57300(x57300, x57299);
  not i57302(x57302, x57199);
  not i57305(x57305, x57304);
  not i57307(x57307, x57204);
  not i57310(x57310, x57309);
  not i57312(x57312, x57209);
  not i57315(x57315, x57314);
  not i57317(x57317, x57214);
  not i57320(x57320, x57319);
  not i57321(x57321, x57221);
  not i57322(x57322, x57224);
  not i57323(x57323, x57227);
  not i57324(x57324, x57230);
  not i57326(x57326, x57233);
  not i57329(x57329, x57238);
  not i57332(x57332, x57243);
  not i57335(x57335, x57248);
  not i57338(x57338, x57253);
  not i57341(x57341, x57258);
  not i57344(x57344, x57263);
  not i57347(x57347, x57268);
  not i57350(x57350, x57273);
  not i57353(x57353, x57352);
  not i57355(x57355, x57278);
  not i57358(x57358, x57357);
  not i57360(x57360, x57283);
  not i57363(x57363, x57362);
  not i57365(x57365, x57288);
  not i57368(x57368, x57367);
  not i57370(x57370, x57293);
  not i57373(x57373, x57372);
  not i57375(x57375, x57298);
  not i57378(x57378, x57377);
  not i57380(x57380, x57303);
  not i57383(x57383, x57382);
  not i57385(x57385, x57308);
  not i57388(x57388, x57387);
  not i57390(x57390, x57313);
  not i57393(x57393, x57392);
  not i57395(x57395, x57318);
  not i57398(x57398, x57397);
  not i57399(x57399, x57333);
  not i57400(x57400, x57336);
  not i57401(x57401, x57339);
  not i57402(x57402, x57342);
  not i57403(x57403, x57345);
  not i57404(x57404, x57348);
  not i57406(x57406, x57351);
  not i57409(x57409, x57356);
  not i57412(x57412, x57361);
  not i57415(x57415, x57366);
  not i57418(x57418, x57371);
  not i57421(x57421, x57376);
  not i57424(x57424, x57381);
  not i57427(x57427, x57386);
  not i57430(x57430, x57391);
  not i57433(x57433, x57396);
  not i57437(x57437, x57436);
  not i57441(x57441, x57440);
  not i57445(x57445, x57444);
  not i57449(x57449, x57448);
  not i57453(x57453, x57452);
  not i57457(x57457, x57456);
  not i57461(x57461, x57460);
  not i57465(x57465, x57464);
  not i57467(x57467, x57327);
  not i57470(x57470, x57469);
  not i57472(x57472, x57330);
  not i57475(x57475, x57474);
  not i57479(x57479, x57478);
  not i57483(x57483, x57482);
  not i57487(x57487, x57486);
  not i57491(x57491, x57490);
  not i57495(x57495, x57494);
  not i57499(x57499, x57498);
  not i57501(x57501, x57407);
  not i57504(x57504, x57503);
  not i57506(x57506, x57410);
  not i57509(x57509, x57508);
  not i57511(x57511, x57413);
  not i57514(x57514, x57513);
  not i57516(x57516, x57416);
  not i57519(x57519, x57518);
  not i57521(x57521, x57419);
  not i57524(x57524, x57523);
  not i57526(x57526, x57422);
  not i57529(x57529, x57528);
  not i57531(x57531, x57425);
  not i57534(x57534, x57533);
  not i57536(x57536, x57428);
  not i57539(x57539, x57538);
  not i57541(x57541, x57431);
  not i57544(x57544, x57543);
  not i57546(x57546, x57434);
  not i57549(x57549, x57548);
  not i57551(x57551, x57550);
  not i57553(x57553, x57552);
  not i57555(x57555, x57554);
  not i57557(x57557, x57556);
  not i57559(x57559, x57558);
  not i57561(x57561, x57560);
  not i57563(x57563, x57562);
  not i57565(x57565, x57564);
  not i57567(x57567, x57566);
  not i57569(x57569, x57568);
  not i57571(x57571, x57570);
  not i57573(x57573, x57572);
  not i57575(x57575, x57574);
  not i57577(x57577, x57576);
  not i57579(x57579, x57578);
  not i57581(x57581, x57580);
  not i57583(x57583, x57582);
  not i57585(x57585, x57584);
  not i57587(x57587, x57586);
  not i57589(x57589, x57588);
  not i57591(x57591, x57590);
  not i57593(x57593, x57592);
  not i57595(x57595, x57594);
  not i57597(x57597, x57596);
  not i57599(x57599, x57598);
  not i57601(x57601, x57600);
  not i57603(x57603, x57602);
  not i57605(x57605, x57604);
  not i57607(x57607, x57606);
  not i57609(x57609, x57608);
  not i57612(x57612, x57611);
  not i57614(x57614, x57613);
  not i57616(x57616, x57615);
  not i57618(x57618, x57617);
  not i57620(x57620, x57619);
  not i57622(x57622, x57621);
  not i57624(x57624, x57623);
  not i57626(x57626, x57625);
  not i57628(x57628, x57627);
  not i57630(x57630, x57629);
  not i57632(x57632, x57631);
  not i57634(x57634, x57633);
  not i57636(x57636, x57635);
  not i57638(x57638, x57637);
  not i57640(x57640, x57639);
  not i57642(x57642, x57641);
  not i57644(x57644, x57643);
  not i57646(x57646, x57645);
  not i57648(x57648, x57647);
  not i57650(x57650, x57649);
  not i57652(x57652, x57651);
  not i57654(x57654, x57653);
  not i57656(x57656, x57655);
  not i57658(x57658, x57657);
  not i57660(x57660, x57659);
  not i57662(x57662, x57661);
  not i57664(x57664, x57663);
  not i57666(x57666, x57665);
  not i57671(x57671, x57670);
  not i57673(x57673, x57672);
  not i57675(x57675, x57674);
  not i57677(x57677, x57676);
  not i57679(x57679, x57678);
  not i57681(x57681, x57680);
  not i57683(x57683, x57682);
  not i57685(x57685, x57684);
  not i57687(x57687, x57686);
  not i57689(x57689, x57688);
  not i57691(x57691, x57690);
  not i57693(x57693, x57692);
  not i57695(x57695, x57694);
  not i57697(x57697, x57696);
  not i57699(x57699, x57698);
  not i57701(x57701, x57700);
  not i57703(x57703, x57702);
  not i57705(x57705, x57704);
  not i57707(x57707, x57706);
  not i57709(x57709, x57708);
  not i57711(x57711, x57710);
  not i57713(x57713, x57712);
  not i57715(x57715, x57714);
  not i57717(x57717, x57716);
  not i57727(x57727, x57726);
  not i57729(x57729, x57728);
  not i57731(x57731, x57730);
  not i57733(x57733, x57732);
  not i57735(x57735, x57734);
  not i57737(x57737, x57736);
  not i57739(x57739, x57738);
  not i57741(x57741, x57740);
  not i57743(x57743, x57742);
  not i57745(x57745, x57744);
  not i57747(x57747, x57746);
  not i57749(x57749, x57748);
  not i57751(x57751, x57750);
  not i57753(x57753, x57752);
  not i57755(x57755, x57754);
  not i57773(x57773, x57772);
  not i57777(x57777, x57776);
  not i57781(x57781, x57780);
  not i57785(x57785, x57784);
  not i57789(x57789, x57788);
  not i57793(x57793, x57792);
  not i57797(x57797, x57796);
  not i57801(x57801, x57800);
  not i57805(x57805, x57804);
  not i57809(x57809, x57808);
  not i57813(x57813, x57812);
  not i57817(x57817, x57816);
  not i57821(x57821, x57820);
  not i57825(x57825, x57824);
  not i57829(x57829, x57828);
  not i57833(x57833, x57832);
  not i57837(x57837, x57836);
  not i57841(x57841, x57840);
  not i57845(x57845, x57844);
  not i57849(x57849, x57848);
  not i57853(x57853, x57852);
  not i57857(x57857, x57856);
  not i57861(x57861, x57860);
  not i57865(x57865, x57864);
  not i57869(x57869, x57868);
  not i57873(x57873, x57872);
  not i57877(x57877, x57876);
  not i57881(x57881, x57880);
  not i57885(x57885, x57884);
  not i57889(x57889, x57888);
  not i57893(x57893, x57892);
  not i57894(x57894, x50938);
  not i57896(x57896, x57895);
  not i57898(x57898, x57897);
  not i57900(x57900, x57899);
  not i57902(x57902, x57901);
  not i57904(x57904, x57903);
  not i57906(x57906, x57905);
  not i57908(x57908, x57907);
  not i57910(x57910, x57909);
  not i57912(x57912, x57911);
  not i57914(x57914, x57913);
  not i57916(x57916, x57915);
  not i57918(x57918, x57917);
  not i57920(x57920, x57919);
  not i57922(x57922, x57921);
  not i57924(x57924, x57923);
  not i57926(x57926, x57925);
  not i57960(x57960, x57959);
  not i57962(x57962, x57961);
  not i57964(x57964, x57963);
  not i57966(x57966, x57965);
  not i57968(x57968, x57967);
  not i57970(x57970, x57969);
  not i57972(x57972, x57971);
  not i57974(x57974, x57973);
  not i57976(x57976, x57975);
  not i57978(x57978, x57977);
  not i57980(x57980, x57979);
  not i57982(x57982, x57981);
  not i57984(x57984, x57983);
  not i57986(x57986, x57985);
  not i57988(x57988, x57987);
  not i57990(x57990, x57989);
  not i57992(x57992, x57991);
  not i57994(x57994, x57993);
  not i57996(x57996, x57995);
  not i57998(x57998, x57997);
  not i58000(x58000, x57999);
  not i58002(x58002, x58001);
  not i58004(x58004, x58003);
  not i58006(x58006, x58005);
  not i58008(x58008, x58007);
  not i58010(x58010, x58009);
  not i58012(x58012, x58011);
  not i58014(x58014, x58013);
  not i58016(x58016, x58015);
  not i58018(x58018, x58017);
  not i58020(x58020, x58019);
  not i58022(x58022, x58021);
  not i60842(x60842, x68739);
  not i60843(x60843, x74257);
  not i60844(x60844, x74254);
  not i60846(x60846, x74251);
  not i60847(x60847, x74248);
  not i60849(x60849, x74245);
  not i60850(x60850, x74242);
  not i60852(x60852, x74239);
  not i60853(x60853, x74236);
  not i60855(x60855, x74233);
  not i60856(x60856, x74230);
  not i60858(x60858, x74227);
  not i60859(x60859, x74224);
  not i60861(x60861, x74221);
  not i60862(x60862, x74218);
  not i60864(x60864, x74215);
  not i60865(x60865, x74212);
  not i60867(x60867, x74209);
  not i60868(x60868, x74206);
  not i60870(x60870, x74203);
  not i60871(x60871, x74200);
  not i60873(x60873, x74197);
  not i60874(x60874, x74194);
  not i60876(x60876, x74191);
  not i60877(x60877, x74188);
  not i60879(x60879, x74185);
  not i60880(x60880, x74182);
  not i60882(x60882, x74179);
  not i60883(x60883, x74176);
  not i60885(x60885, x74173);
  not i60886(x60886, x74170);
  not i60888(x60888, x74167);
  not i60889(x60889, x74164);
  not i60891(x60891, x60845);
  not i60892(x60892, x60848);
  not i60894(x60894, x60851);
  not i60895(x60895, x60854);
  not i60897(x60897, x60857);
  not i60898(x60898, x60860);
  not i60900(x60900, x60863);
  not i60901(x60901, x60866);
  not i60903(x60903, x60869);
  not i60904(x60904, x60872);
  not i60906(x60906, x60875);
  not i60907(x60907, x60878);
  not i60909(x60909, x60881);
  not i60910(x60910, x60884);
  not i60912(x60912, x60887);
  not i60913(x60913, x60890);
  not i60915(x60915, x60893);
  not i60916(x60916, x60896);
  not i60918(x60918, x60899);
  not i60919(x60919, x60902);
  not i60921(x60921, x60905);
  not i60922(x60922, x60908);
  not i60924(x60924, x60911);
  not i60925(x60925, x60914);
  not i60927(x60927, x60917);
  not i60928(x60928, x60920);
  not i60930(x60930, x60923);
  not i60931(x60931, x60926);
  not i60933(x60933, x60929);
  not i60934(x60934, x60932);
  not i60937(x60937, x60936);
  not i60938(x60938, x74455);
  not i60939(x60939, x74452);
  not i60942(x60942, x60941);
  not i60943(x60943, x60935);
  not i60944(x60944, x74122);
  not i60955(x60955, x74125);
  not i60962(x60962, x74128);
  not i60967(x60967, x74131);
  not i60970(x60970, x74134);
  not i60977(x60977, x74551);
  not i60978(x60978, x74548);
  not i60980(x60980, x74545);
  not i60981(x60981, x74542);
  not i60983(x60983, x74539);
  not i60984(x60984, x74536);
  not i60986(x60986, x74533);
  not i60987(x60987, x74530);
  not i60989(x60989, x74527);
  not i60990(x60990, x74524);
  not i60992(x60992, x74521);
  not i60993(x60993, x74518);
  not i60995(x60995, x74515);
  not i60996(x60996, x74512);
  not i60998(x60998, x74509);
  not i60999(x60999, x74506);
  not i61001(x61001, x74503);
  not i61002(x61002, x74500);
  not i61004(x61004, x74497);
  not i61005(x61005, x74494);
  not i61007(x61007, x74491);
  not i61008(x61008, x74488);
  not i61010(x61010, x74485);
  not i61011(x61011, x74482);
  not i61013(x61013, x74479);
  not i61014(x61014, x74476);
  not i61016(x61016, x74473);
  not i61017(x61017, x74470);
  not i61019(x61019, x74467);
  not i61020(x61020, x74464);
  not i61022(x61022, x74461);
  not i61023(x61023, x74458);
  not i61025(x61025, x60979);
  not i61026(x61026, x60982);
  not i61028(x61028, x60985);
  not i61029(x61029, x60988);
  not i61031(x61031, x60991);
  not i61032(x61032, x60994);
  not i61034(x61034, x60997);
  not i61035(x61035, x61000);
  not i61037(x61037, x61003);
  not i61038(x61038, x61006);
  not i61040(x61040, x61009);
  not i61041(x61041, x61012);
  not i61043(x61043, x61015);
  not i61044(x61044, x61018);
  not i61046(x61046, x61021);
  not i61047(x61047, x61024);
  not i61049(x61049, x61027);
  not i61050(x61050, x61030);
  not i61052(x61052, x61033);
  not i61053(x61053, x61036);
  not i61055(x61055, x61039);
  not i61056(x61056, x61042);
  not i61058(x61058, x61045);
  not i61059(x61059, x61048);
  not i61061(x61061, x61051);
  not i61062(x61062, x61054);
  not i61064(x61064, x61057);
  not i61065(x61065, x61060);
  not i61067(x61067, x61063);
  not i61068(x61068, x61066);
  not i61071(x61071, x61070);
  not i61072(x61072, x74749);
  not i61073(x61073, x74746);
  not i61076(x61076, x61075);
  not i61077(x61077, x61069);
  not i61106(x61106, x74845);
  not i61107(x61107, x74842);
  not i61109(x61109, x74839);
  not i61110(x61110, x74836);
  not i61112(x61112, x74833);
  not i61113(x61113, x74830);
  not i61115(x61115, x74827);
  not i61116(x61116, x74824);
  not i61118(x61118, x74821);
  not i61119(x61119, x74818);
  not i61121(x61121, x74815);
  not i61122(x61122, x74812);
  not i61124(x61124, x74809);
  not i61125(x61125, x74806);
  not i61127(x61127, x74803);
  not i61128(x61128, x74800);
  not i61130(x61130, x74797);
  not i61131(x61131, x74794);
  not i61133(x61133, x74791);
  not i61134(x61134, x74788);
  not i61136(x61136, x74785);
  not i61137(x61137, x74782);
  not i61139(x61139, x74779);
  not i61140(x61140, x74776);
  not i61142(x61142, x74773);
  not i61143(x61143, x74770);
  not i61145(x61145, x74767);
  not i61146(x61146, x74764);
  not i61148(x61148, x74761);
  not i61149(x61149, x74758);
  not i61151(x61151, x74755);
  not i61152(x61152, x74752);
  not i61154(x61154, x61108);
  not i61155(x61155, x61111);
  not i61157(x61157, x61114);
  not i61158(x61158, x61117);
  not i61160(x61160, x61120);
  not i61161(x61161, x61123);
  not i61163(x61163, x61126);
  not i61164(x61164, x61129);
  not i61166(x61166, x61132);
  not i61167(x61167, x61135);
  not i61169(x61169, x61138);
  not i61170(x61170, x61141);
  not i61172(x61172, x61144);
  not i61173(x61173, x61147);
  not i61175(x61175, x61150);
  not i61176(x61176, x61153);
  not i61178(x61178, x61156);
  not i61179(x61179, x61159);
  not i61181(x61181, x61162);
  not i61182(x61182, x61165);
  not i61184(x61184, x61168);
  not i61185(x61185, x61171);
  not i61187(x61187, x61174);
  not i61188(x61188, x61177);
  not i61190(x61190, x61180);
  not i61191(x61191, x61183);
  not i61193(x61193, x61186);
  not i61194(x61194, x61189);
  not i61196(x61196, x61192);
  not i61197(x61197, x61195);
  not i61200(x61200, x61199);
  not i61201(x61201, x75043);
  not i61202(x61202, x75040);
  not i61205(x61205, x61204);
  not i61206(x61206, x61198);
  not i61235(x61235, x75139);
  not i61236(x61236, x75136);
  not i61238(x61238, x75133);
  not i61239(x61239, x75130);
  not i61241(x61241, x75127);
  not i61242(x61242, x75124);
  not i61244(x61244, x75121);
  not i61245(x61245, x75118);
  not i61247(x61247, x75115);
  not i61248(x61248, x75112);
  not i61250(x61250, x75109);
  not i61251(x61251, x75106);
  not i61253(x61253, x75103);
  not i61254(x61254, x75100);
  not i61256(x61256, x75097);
  not i61257(x61257, x75094);
  not i61259(x61259, x75091);
  not i61260(x61260, x75088);
  not i61262(x61262, x75085);
  not i61263(x61263, x75082);
  not i61265(x61265, x75079);
  not i61266(x61266, x75076);
  not i61268(x61268, x75073);
  not i61269(x61269, x75070);
  not i61271(x61271, x75067);
  not i61272(x61272, x75064);
  not i61274(x61274, x75061);
  not i61275(x61275, x75058);
  not i61277(x61277, x75055);
  not i61278(x61278, x75052);
  not i61280(x61280, x75049);
  not i61281(x61281, x75046);
  not i61283(x61283, x61237);
  not i61284(x61284, x61240);
  not i61286(x61286, x61243);
  not i61287(x61287, x61246);
  not i61289(x61289, x61249);
  not i61290(x61290, x61252);
  not i61292(x61292, x61255);
  not i61293(x61293, x61258);
  not i61295(x61295, x61261);
  not i61296(x61296, x61264);
  not i61298(x61298, x61267);
  not i61299(x61299, x61270);
  not i61301(x61301, x61273);
  not i61302(x61302, x61276);
  not i61304(x61304, x61279);
  not i61305(x61305, x61282);
  not i61307(x61307, x61285);
  not i61308(x61308, x61288);
  not i61310(x61310, x61291);
  not i61311(x61311, x61294);
  not i61313(x61313, x61297);
  not i61314(x61314, x61300);
  not i61316(x61316, x61303);
  not i61317(x61317, x61306);
  not i61319(x61319, x61309);
  not i61320(x61320, x61312);
  not i61322(x61322, x61315);
  not i61323(x61323, x61318);
  not i61325(x61325, x61321);
  not i61326(x61326, x61324);
  not i61329(x61329, x61328);
  not i61330(x61330, x75337);
  not i61331(x61331, x75334);
  not i61334(x61334, x61333);
  not i61335(x61335, x61327);
  not i61425(x61425, x68740);
  not i61427(x61427, x61426);
  not i61686(x61686, x75436);
  not i61975(x61975, x75457);
  not i62931(x62931, x68741);
  not i62933(x62933, x76792);
  not i63027(x63027, x62935);
  not i63028(x63028, x76675);
  not i63032(x63032, x62938);
  not i63033(x63033, x76678);
  not i63036(x63036, x63035);
  not i63038(x63038, x62941);
  not i63039(x63039, x76681);
  not i63042(x63042, x63041);
  not i63044(x63044, x62944);
  not i63045(x63045, x76684);
  not i63048(x63048, x63047);
  not i63050(x63050, x62947);
  not i63051(x63051, x76687);
  not i63054(x63054, x63053);
  not i63056(x63056, x62950);
  not i63057(x63057, x76690);
  not i63060(x63060, x63059);
  not i63062(x63062, x62953);
  not i63063(x63063, x76693);
  not i63066(x63066, x63065);
  not i63068(x63068, x62956);
  not i63069(x63069, x76696);
  not i63072(x63072, x63071);
  not i63074(x63074, x62959);
  not i63075(x63075, x76699);
  not i63078(x63078, x63077);
  not i63080(x63080, x62962);
  not i63081(x63081, x76702);
  not i63084(x63084, x63083);
  not i63086(x63086, x62965);
  not i63087(x63087, x76705);
  not i63090(x63090, x63089);
  not i63092(x63092, x62968);
  not i63093(x63093, x76708);
  not i63096(x63096, x63095);
  not i63098(x63098, x62971);
  not i63099(x63099, x76711);
  not i63102(x63102, x63101);
  not i63104(x63104, x62974);
  not i63105(x63105, x76714);
  not i63108(x63108, x63107);
  not i63110(x63110, x62977);
  not i63111(x63111, x76717);
  not i63114(x63114, x63113);
  not i63116(x63116, x62980);
  not i63117(x63117, x76720);
  not i63120(x63120, x63119);
  not i63122(x63122, x62983);
  not i63123(x63123, x76723);
  not i63126(x63126, x63125);
  not i63128(x63128, x62986);
  not i63129(x63129, x76726);
  not i63132(x63132, x63131);
  not i63134(x63134, x62989);
  not i63135(x63135, x76729);
  not i63138(x63138, x63137);
  not i63140(x63140, x62992);
  not i63141(x63141, x76732);
  not i63144(x63144, x63143);
  not i63146(x63146, x62995);
  not i63147(x63147, x76735);
  not i63150(x63150, x63149);
  not i63152(x63152, x62998);
  not i63153(x63153, x76738);
  not i63156(x63156, x63155);
  not i63158(x63158, x63001);
  not i63159(x63159, x76741);
  not i63162(x63162, x63161);
  not i63164(x63164, x63004);
  not i63165(x63165, x76744);
  not i63168(x63168, x63167);
  not i63170(x63170, x63007);
  not i63171(x63171, x76747);
  not i63174(x63174, x63173);
  not i63176(x63176, x63010);
  not i63177(x63177, x76750);
  not i63180(x63180, x63179);
  not i63182(x63182, x63013);
  not i63183(x63183, x76753);
  not i63186(x63186, x63185);
  not i63188(x63188, x63016);
  not i63189(x63189, x76756);
  not i63192(x63192, x63191);
  not i63194(x63194, x63019);
  not i63195(x63195, x76759);
  not i63198(x63198, x63197);
  not i63200(x63200, x63022);
  not i63201(x63201, x76762);
  not i63204(x63204, x63203);
  not i63206(x63206, x63025);
  not i63207(x63207, x76765);
  not i63210(x63210, x63209);
  not i63211(x63211, x63026);
  not i63212(x63212, x63031);
  not i63213(x63213, x63037);
  not i63214(x63214, x63043);
  not i63215(x63215, x63049);
  not i63216(x63216, x63055);
  not i63217(x63217, x63061);
  not i63218(x63218, x63067);
  not i63219(x63219, x63073);
  not i63220(x63220, x63079);
  not i63221(x63221, x63085);
  not i63222(x63222, x63091);
  not i63223(x63223, x63097);
  not i63224(x63224, x63103);
  not i63225(x63225, x63109);
  not i63226(x63226, x63115);
  not i63227(x63227, x63121);
  not i63228(x63228, x63127);
  not i63229(x63229, x63133);
  not i63230(x63230, x63139);
  not i63231(x63231, x63145);
  not i63232(x63232, x63151);
  not i63233(x63233, x63157);
  not i63234(x63234, x63163);
  not i63235(x63235, x63169);
  not i63236(x63236, x63175);
  not i63237(x63237, x63181);
  not i63238(x63238, x63187);
  not i63239(x63239, x63193);
  not i63245(x63245, x63244);
  not i63249(x63249, x63248);
  not i63253(x63253, x63252);
  not i63257(x63257, x63256);
  not i63261(x63261, x63260);
  not i63265(x63265, x63264);
  not i63269(x63269, x63268);
  not i63273(x63273, x63272);
  not i63277(x63277, x63276);
  not i63281(x63281, x63280);
  not i63285(x63285, x63284);
  not i63289(x63289, x63288);
  not i63293(x63293, x63292);
  not i63297(x63297, x63296);
  not i63301(x63301, x63300);
  not i63305(x63305, x63304);
  not i63309(x63309, x63308);
  not i63313(x63313, x63312);
  not i63317(x63317, x63316);
  not i63321(x63321, x63320);
  not i63325(x63325, x63324);
  not i63329(x63329, x63328);
  not i63333(x63333, x63332);
  not i63337(x63337, x63336);
  not i63341(x63341, x63340);
  not i63345(x63345, x63344);
  not i63349(x63349, x63348);
  not i63353(x63353, x63352);
  not i63354(x63354, x63241);
  not i63356(x63356, x63243);
  not i63359(x63359, x63247);
  not i63362(x63362, x63251);
  not i63365(x63365, x63364);
  not i63367(x63367, x63255);
  not i63370(x63370, x63369);
  not i63372(x63372, x63259);
  not i63375(x63375, x63374);
  not i63377(x63377, x63263);
  not i63380(x63380, x63379);
  not i63382(x63382, x63267);
  not i63385(x63385, x63384);
  not i63387(x63387, x63271);
  not i63390(x63390, x63389);
  not i63392(x63392, x63275);
  not i63395(x63395, x63394);
  not i63397(x63397, x63279);
  not i63400(x63400, x63399);
  not i63402(x63402, x63283);
  not i63405(x63405, x63404);
  not i63407(x63407, x63287);
  not i63410(x63410, x63409);
  not i63412(x63412, x63291);
  not i63415(x63415, x63414);
  not i63417(x63417, x63295);
  not i63420(x63420, x63419);
  not i63422(x63422, x63299);
  not i63425(x63425, x63424);
  not i63427(x63427, x63303);
  not i63430(x63430, x63429);
  not i63432(x63432, x63307);
  not i63435(x63435, x63434);
  not i63437(x63437, x63311);
  not i63440(x63440, x63439);
  not i63442(x63442, x63315);
  not i63445(x63445, x63444);
  not i63447(x63447, x63319);
  not i63450(x63450, x63449);
  not i63452(x63452, x63323);
  not i63455(x63455, x63454);
  not i63457(x63457, x63327);
  not i63460(x63460, x63459);
  not i63462(x63462, x63331);
  not i63465(x63465, x63464);
  not i63467(x63467, x63335);
  not i63470(x63470, x63469);
  not i63472(x63472, x63339);
  not i63475(x63475, x63474);
  not i63477(x63477, x63343);
  not i63480(x63480, x63479);
  not i63482(x63482, x63347);
  not i63485(x63485, x63484);
  not i63487(x63487, x63351);
  not i63490(x63490, x63489);
  not i63491(x63491, x63360);
  not i63493(x63493, x63363);
  not i63496(x63496, x63368);
  not i63499(x63499, x63373);
  not i63502(x63502, x63378);
  not i63505(x63505, x63383);
  not i63508(x63508, x63507);
  not i63510(x63510, x63388);
  not i63513(x63513, x63512);
  not i63515(x63515, x63393);
  not i63518(x63518, x63517);
  not i63520(x63520, x63398);
  not i63523(x63523, x63522);
  not i63525(x63525, x63403);
  not i63528(x63528, x63527);
  not i63530(x63530, x63408);
  not i63533(x63533, x63532);
  not i63535(x63535, x63413);
  not i63538(x63538, x63537);
  not i63540(x63540, x63418);
  not i63543(x63543, x63542);
  not i63545(x63545, x63423);
  not i63548(x63548, x63547);
  not i63550(x63550, x63428);
  not i63553(x63553, x63552);
  not i63555(x63555, x63433);
  not i63558(x63558, x63557);
  not i63560(x63560, x63438);
  not i63563(x63563, x63562);
  not i63565(x63565, x63443);
  not i63568(x63568, x63567);
  not i63570(x63570, x63448);
  not i63573(x63573, x63572);
  not i63575(x63575, x63453);
  not i63578(x63578, x63577);
  not i63580(x63580, x63458);
  not i63583(x63583, x63582);
  not i63585(x63585, x63463);
  not i63588(x63588, x63587);
  not i63590(x63590, x63468);
  not i63593(x63593, x63592);
  not i63595(x63595, x63473);
  not i63598(x63598, x63597);
  not i63600(x63600, x63478);
  not i63603(x63603, x63602);
  not i63605(x63605, x63483);
  not i63608(x63608, x63607);
  not i63610(x63610, x63488);
  not i63613(x63613, x63612);
  not i63614(x63614, x63503);
  not i63616(x63616, x63506);
  not i63619(x63619, x63511);
  not i63622(x63622, x63516);
  not i63625(x63625, x63521);
  not i63628(x63628, x63526);
  not i63631(x63631, x63531);
  not i63634(x63634, x63536);
  not i63637(x63637, x63541);
  not i63640(x63640, x63546);
  not i63643(x63643, x63642);
  not i63645(x63645, x63551);
  not i63648(x63648, x63647);
  not i63650(x63650, x63556);
  not i63653(x63653, x63652);
  not i63655(x63655, x63561);
  not i63658(x63658, x63657);
  not i63660(x63660, x63566);
  not i63663(x63663, x63662);
  not i63665(x63665, x63571);
  not i63668(x63668, x63667);
  not i63670(x63670, x63576);
  not i63673(x63673, x63672);
  not i63675(x63675, x63581);
  not i63678(x63678, x63677);
  not i63680(x63680, x63586);
  not i63683(x63683, x63682);
  not i63685(x63685, x63591);
  not i63688(x63688, x63687);
  not i63690(x63690, x63596);
  not i63693(x63693, x63692);
  not i63695(x63695, x63601);
  not i63698(x63698, x63697);
  not i63700(x63700, x63606);
  not i63703(x63703, x63702);
  not i63705(x63705, x63611);
  not i63708(x63708, x63707);
  not i63709(x63709, x63638);
  not i63711(x63711, x63641);
  not i63714(x63714, x63646);
  not i63717(x63717, x63651);
  not i63720(x63720, x63656);
  not i63723(x63723, x63661);
  not i63726(x63726, x63666);
  not i63729(x63729, x63671);
  not i63732(x63732, x63676);
  not i63735(x63735, x63681);
  not i63738(x63738, x63686);
  not i63741(x63741, x63691);
  not i63744(x63744, x63696);
  not i63747(x63747, x63701);
  not i63750(x63750, x63706);
  not i63757(x63757, x63756);
  not i63759(x63759, x63357);
  not i63762(x63762, x63761);
  not i63766(x63766, x63765);
  not i63768(x63768, x63494);
  not i63771(x63771, x63770);
  not i63773(x63773, x63497);
  not i63776(x63776, x63775);
  not i63778(x63778, x63500);
  not i63781(x63781, x63780);
  not i63785(x63785, x63784);
  not i63787(x63787, x63617);
  not i63790(x63790, x63789);
  not i63792(x63792, x63620);
  not i63796(x63796, x63623);
  not i63800(x63800, x63626);
  not i63804(x63804, x63629);
  not i63808(x63808, x63632);
  not i63812(x63812, x63635);
  not i63819(x63819, x63712);
  not i63823(x63823, x63715);
  not i63827(x63827, x63718);
  not i63831(x63831, x63721);
  not i63835(x63835, x63724);
  not i63839(x63839, x63727);
  not i63843(x63843, x63730);
  not i63847(x63847, x63733);
  not i63851(x63851, x63736);
  not i63855(x63855, x63739);
  not i63859(x63859, x63742);
  not i63863(x63863, x63745);
  not i63867(x63867, x63748);
  not i63871(x63871, x63751);
  not i63875(x63875, x63874);
  not i63914(x63914, x63908);
  not i64009(x64009, x63909);
  not i64102(x64102, x63910);
  not i64191(x64191, x63911);
  not i64272(x64272, x63912);
  not i64337(x64337, x64336);
  not i64339(x64339, x64338);
  not i64341(x64341, x64340);
  not i64343(x64343, x64342);
  not i64345(x64345, x64344);
  not i64347(x64347, x64346);
  not i64349(x64349, x64348);
  not i64351(x64351, x64350);
  not i64353(x64353, x64352);
  not i64355(x64355, x64354);
  not i64357(x64357, x64356);
  not i64359(x64359, x64358);
  not i64361(x64361, x64360);
  not i64363(x64363, x64362);
  not i64365(x64365, x64364);
  not i64367(x64367, x64366);
  not i64369(x64369, x64368);
  not i64371(x64371, x64370);
  not i64373(x64373, x64372);
  not i64375(x64375, x64374);
  not i64377(x64377, x64376);
  not i64379(x64379, x64378);
  not i64381(x64381, x64380);
  not i64383(x64383, x64382);
  not i64385(x64385, x64384);
  not i64387(x64387, x64386);
  not i64389(x64389, x64388);
  not i64391(x64391, x64390);
  not i64393(x64393, x64392);
  not i64395(x64395, x64394);
  not i64397(x64397, x64396);
  not i64429(x64429, x64400);
  not i64433(x64433, x64403);
  not i64436(x64436, x64435);
  not i64438(x64438, x64406);
  not i64441(x64441, x64440);
  not i64443(x64443, x64409);
  not i64446(x64446, x64445);
  not i64448(x64448, x64412);
  not i64451(x64451, x64450);
  not i64453(x64453, x64415);
  not i64456(x64456, x64455);
  not i64458(x64458, x64418);
  not i64461(x64461, x64460);
  not i64463(x64463, x64421);
  not i64466(x64466, x64465);
  not i64468(x64468, x64424);
  not i64471(x64471, x64470);
  not i64473(x64473, x64427);
  not i64476(x64476, x64475);
  not i64477(x64477, x64428);
  not i64478(x64478, x64432);
  not i64479(x64479, x64437);
  not i64480(x64480, x64442);
  not i64481(x64481, x64447);
  not i64482(x64482, x64452);
  not i64483(x64483, x64457);
  not i64484(x64484, x64462);
  not i64490(x64490, x64489);
  not i64494(x64494, x64493);
  not i64498(x64498, x64497);
  not i64502(x64502, x64501);
  not i64506(x64506, x64505);
  not i64510(x64510, x64509);
  not i64514(x64514, x64513);
  not i64515(x64515, x64486);
  not i64517(x64517, x64488);
  not i64520(x64520, x64492);
  not i64523(x64523, x64496);
  not i64526(x64526, x64525);
  not i64528(x64528, x64500);
  not i64531(x64531, x64530);
  not i64533(x64533, x64504);
  not i64536(x64536, x64535);
  not i64538(x64538, x64508);
  not i64541(x64541, x64540);
  not i64543(x64543, x64512);
  not i64546(x64546, x64545);
  not i64547(x64547, x64521);
  not i64549(x64549, x64524);
  not i64552(x64552, x64529);
  not i64555(x64555, x64534);
  not i64558(x64558, x64539);
  not i64561(x64561, x64544);
  not i64564(x64564, x64563);
  not i64565(x64565, x64559);
  not i64567(x64567, x64562);
  not i64574(x64574, x64573);
  not i64576(x64576, x64518);
  not i64579(x64579, x64578);
  not i64583(x64583, x64582);
  not i64585(x64585, x64550);
  not i64588(x64588, x64587);
  not i64590(x64590, x64553);
  not i64593(x64593, x64592);
  not i64595(x64595, x64556);
  not i64598(x64598, x64597);
  not i64602(x64602, x64601);
  not i64604(x64604, x64568);
  not i64607(x64607, x64606);
  not i64646(x64646, x64640);
  not i64741(x64741, x64641);
  not i64834(x64834, x64642);
  not i64923(x64923, x64643);
  not i65004(x65004, x64644);
  not i65099(x65099, x65070);
  not i65103(x65103, x65073);
  not i65106(x65106, x65105);
  not i65108(x65108, x65076);
  not i65111(x65111, x65110);
  not i65113(x65113, x65079);
  not i65116(x65116, x65115);
  not i65118(x65118, x65082);
  not i65121(x65121, x65120);
  not i65123(x65123, x65085);
  not i65126(x65126, x65125);
  not i65128(x65128, x65088);
  not i65131(x65131, x65130);
  not i65133(x65133, x65091);
  not i65136(x65136, x65135);
  not i65138(x65138, x65094);
  not i65141(x65141, x65140);
  not i65143(x65143, x65097);
  not i65146(x65146, x65145);
  not i65147(x65147, x65098);
  not i65148(x65148, x65102);
  not i65149(x65149, x65107);
  not i65150(x65150, x65112);
  not i65151(x65151, x65117);
  not i65152(x65152, x65122);
  not i65153(x65153, x65127);
  not i65154(x65154, x65132);
  not i65160(x65160, x65159);
  not i65164(x65164, x65163);
  not i65168(x65168, x65167);
  not i65172(x65172, x65171);
  not i65176(x65176, x65175);
  not i65180(x65180, x65179);
  not i65184(x65184, x65183);
  not i65185(x65185, x65156);
  not i65187(x65187, x65158);
  not i65190(x65190, x65162);
  not i65193(x65193, x65166);
  not i65196(x65196, x65195);
  not i65198(x65198, x65170);
  not i65201(x65201, x65200);
  not i65203(x65203, x65174);
  not i65206(x65206, x65205);
  not i65208(x65208, x65178);
  not i65211(x65211, x65210);
  not i65213(x65213, x65182);
  not i65216(x65216, x65215);
  not i65217(x65217, x65191);
  not i65219(x65219, x65194);
  not i65222(x65222, x65199);
  not i65225(x65225, x65204);
  not i65228(x65228, x65209);
  not i65231(x65231, x65214);
  not i65234(x65234, x65233);
  not i65235(x65235, x65229);
  not i65237(x65237, x65232);
  not i65244(x65244, x65243);
  not i65246(x65246, x65188);
  not i65249(x65249, x65248);
  not i65253(x65253, x65252);
  not i65255(x65255, x65220);
  not i65258(x65258, x65257);
  not i65260(x65260, x65223);
  not i65263(x65263, x65262);
  not i65265(x65265, x65226);
  not i65268(x65268, x65267);
  not i65272(x65272, x65271);
  not i65274(x65274, x65238);
  not i65277(x65277, x65276);
  not i65316(x65316, x65310);
  not i65411(x65411, x65311);
  not i65504(x65504, x65312);
  not i65593(x65593, x65313);
  not i65674(x65674, x65314);
  not i65769(x65769, x65740);
  not i65773(x65773, x65743);
  not i65776(x65776, x65775);
  not i65778(x65778, x65746);
  not i65781(x65781, x65780);
  not i65783(x65783, x65749);
  not i65786(x65786, x65785);
  not i65788(x65788, x65752);
  not i65791(x65791, x65790);
  not i65793(x65793, x65755);
  not i65796(x65796, x65795);
  not i65798(x65798, x65758);
  not i65801(x65801, x65800);
  not i65803(x65803, x65761);
  not i65806(x65806, x65805);
  not i65808(x65808, x65764);
  not i65811(x65811, x65810);
  not i65813(x65813, x65767);
  not i65816(x65816, x65815);
  not i65817(x65817, x65768);
  not i65818(x65818, x65772);
  not i65819(x65819, x65777);
  not i65820(x65820, x65782);
  not i65821(x65821, x65787);
  not i65822(x65822, x65792);
  not i65823(x65823, x65797);
  not i65824(x65824, x65802);
  not i65830(x65830, x65829);
  not i65834(x65834, x65833);
  not i65838(x65838, x65837);
  not i65842(x65842, x65841);
  not i65846(x65846, x65845);
  not i65850(x65850, x65849);
  not i65854(x65854, x65853);
  not i65855(x65855, x65826);
  not i65857(x65857, x65828);
  not i65860(x65860, x65832);
  not i65863(x65863, x65836);
  not i65866(x65866, x65865);
  not i65868(x65868, x65840);
  not i65871(x65871, x65870);
  not i65873(x65873, x65844);
  not i65876(x65876, x65875);
  not i65878(x65878, x65848);
  not i65881(x65881, x65880);
  not i65883(x65883, x65852);
  not i65886(x65886, x65885);
  not i65887(x65887, x65861);
  not i65889(x65889, x65864);
  not i65892(x65892, x65869);
  not i65895(x65895, x65874);
  not i65898(x65898, x65879);
  not i65901(x65901, x65884);
  not i65904(x65904, x65903);
  not i65905(x65905, x65899);
  not i65907(x65907, x65902);
  not i65914(x65914, x65913);
  not i65916(x65916, x65858);
  not i65919(x65919, x65918);
  not i65923(x65923, x65922);
  not i65925(x65925, x65890);
  not i65928(x65928, x65927);
  not i65930(x65930, x65893);
  not i65933(x65933, x65932);
  not i65935(x65935, x65896);
  not i65938(x65938, x65937);
  not i65942(x65942, x65941);
  not i65944(x65944, x65908);
  not i65947(x65947, x65946);
  not i65986(x65986, x65980);
  not i66081(x66081, x65981);
  not i66174(x66174, x65982);
  not i66263(x66263, x65983);
  not i66344(x66344, x65984);
  not i66409(x66409, x66408);
  not i66470(x66470, x68742);
  not i66472(x66472, x66471);
  not i66603(x66603, x78106);
  not i67463(x67463, x68743);
  not i67465(x67465, x67464);
  not i67596(x67596, x79441);
  not i68458(x68458, x68456);
  not i68459(x68459, x68457);
  not i68461(x68461, x68460);
  not i68464(x68464, x68463);
  not i68467(x68467, x68466);
  not i68469(x68469, x68468);
  not i68470(x68470, x68618);
  not i68471(x68471, x68619);
  not i68473(x68473, x68472);
  not i68475(x68475, x68620);
  not i68478(x68478, x68477);
  not i68480(x68480, x68621);
  not i68483(x68483, x68482);
  not i68485(x68485, x68622);
  not i68488(x68488, x68487);
  not i68491(x68491, x68476);
  not i68494(x68494, x68481);
  not i68498(x68498, x68486);
  not i68501(x68501, x68500);
  not i68502(x68502, x68495);
  not i68505(x68505, x68499);
  not i68509(x68509, x68508);
  not i68511(x68511, x68489);
  not i68514(x68514, x68513);
  not i68516(x68516, x68492);
  not i68519(x68519, x68518);
  not i68521(x68521, x68503);
  not i68524(x68524, x68523);
  not i68526(x68526, x68506);
  not i68529(x68529, x68528);
  not i68530(x68530, x68623);
  not i68533(x68533, x68532);
  not i68535(x68535, x68534);
  not i68537(x68537, x68536);
  not i68541(x68541, x68540);
  not i68545(x68545, x68544);
  not i68549(x68549, x68548);
  not i68553(x68553, x68552);
  not i68557(x68557, x68556);
  not i68561(x68561, x68560);
  not i68563(x68563, x71128);
  not i68570(x68570, x83382);
  not i68624(x68624, x60824);
  not i68625(x68625, x61407);
  not i68626(x68626, x62913);
  not i68627(x68627, x66453);
  not i68628(x68628, x67445);
  not i68629(x68629, x68438);
  not i68639(x68639, x68636);
  not i68640(x68640, x68637);
  not i68641(x68641, x68638);
  not i68643(x68643, x68642);
  not i68654(x68654, x68651);
  not i68655(x68655, x68652);
  not i68656(x68656, x68653);
  not i68658(x68658, x68657);
  not i68660(x68660, x68631);
  not i68661(x68661, x68632);
  not i68662(x68662, x68633);
  not i68663(x68663, x68635);
  not i68671(x68671, x68670);
  not i68677(x68677, x68675);
  not i68679(x68679, x68678);
  not i68681(x68681, x68646);
  not i68682(x68682, x68647);
  not i68683(x68683, x68648);
  not i68684(x68684, x68650);
  not i68692(x68692, x68691);
  not i68698(x68698, x68696);
  not i68700(x68700, x68699);
  not i68702(x68702, x68630);
  not i68703(x68703, x68634);
  not i68720(x68720, x68645);
  not i68721(x68721, x68649);
  not i68745(x68745, x68680);
  not i68810(x68810, x68701);
  not i71027(x71027, x14990);
  not i71028(x71028, x70737);
  not i71032(x71032, x15011);
  not i71033(x71033, x70753);
  not i71037(x71037, x15032);
  not i71038(x71038, x70769);
  not i71042(x71042, x15053);
  not i71043(x71043, x70785);
  not i71047(x71047, x15074);
  not i71048(x71048, x70801);
  not i71052(x71052, x15095);
  not i71053(x71053, x70817);
  not i71057(x71057, x71056);
  not i71059(x71059, x71058);
  not i71061(x71061, x71060);
  not i71063(x71063, x71062);
  not i71065(x71065, x71064);
  not i71067(x71067, x71066);
  not i71069(x71069, x71068);
  not i71071(x71071, x71070);
  not i71073(x71073, x71072);
  not i71075(x71075, x71074);
  not i71077(x71077, x2137);
  not i71078(x71078, x70945);
  not i71082(x71082, x2158);
  not i71083(x71083, x70961);
  not i71087(x71087, x2179);
  not i71088(x71088, x70977);
  not i71092(x71092, x2200);
  not i71093(x71093, x70993);
  not i71097(x71097, x2221);
  not i71098(x71098, x71009);
  not i71102(x71102, x2242);
  not i71103(x71103, x71025);
  not i71107(x71107, x71106);
  not i71109(x71109, x71108);
  not i71111(x71111, x71110);
  not i71113(x71113, x71112);
  not i71115(x71115, x71114);
  not i71117(x71117, x71116);
  not i71119(x71119, x71118);
  not i71121(x71121, x71120);
  not i71123(x71123, x71122);
  not i71125(x71125, x71124);
  not i71126(x71126, x68659);
  not i71127(x71127, x68644);
  not i71132(x71132, x71130);
  not i71133(x71133, x71129);
  not i71135(x71135, x68462);
  not i71136(x71136, x71131);
  not i71138(x71138, x71137);
  not i71139(x71139, x71134);
  not i83383(x83383, x9);
  not i83384(x83384, x16);
  not i83385(x83385, x17);
  not i83386(x83386, x20);
  not i83387(x83387, x94);
  not i83388(x83388, x149);
  not i83389(x83389, x150);
  not i83390(x83390, x201);
  not i83391(x83391, x202);
  not i83392(x83392, x203);
  not i83393(x83393, x204);
  not i83394(x83394, x247);
  not i83395(x83395, x248);
  not i83396(x83396, x249);
  not i83397(x83397, x250);
  not i83398(x83398, x251);
  not i83399(x83399, x252);
  not i83400(x83400, x253);
  not i83401(x83401, x254);
  not i83402(x83402, x281);
  not i83403(x83403, x282);
  not i83404(x83404, x283);
  not i83405(x83405, x284);
  not i83406(x83406, x285);
  not i83407(x83407, x286);
  not i83408(x83408, x287);
  not i83409(x83409, x288);
  not i83410(x83410, x289);
  not i83411(x83411, x290);
  not i83412(x83412, x291);
  not i83413(x83413, x292);
  not i83414(x83414, x293);
  not i83415(x83415, x638);
  not i83416(x83416, x641);
  not i83417(x83417, x658);
  not i83418(x83418, x659);
  not i83419(x83419, x660);
  not i83420(x83420, x661);
  not i83421(x83421, x680);
  not i83422(x83422, x294);
  not i83423(x83423, x681);
  not i83424(x83424, x682);
  not i83425(x83425, x686);
  not i83426(x83426, x690);
  not i83427(x83427, x694);
  not i83428(x83428, x695);
  not i83429(x83429, x696);
  not i83430(x83430, x697);
  not i83431(x83431, x700);
  not i83432(x83432, x701);
  not i83433(x83433, x705);
  not i83434(x83434, x706);
  not i83435(x83435, x707);
  not i83436(x83436, x708);
  not i83437(x83437, x709);
  not i83438(x83438, x712);
  not i83439(x83439, x724);
  not i83440(x83440, x725);
  not i83441(x83441, x726);
  not i83442(x83442, x728);
  not i83443(x83443, x297);
  not i83444(x83444, x729);
  not i83445(x83445, x738);
  not i83446(x83446, x739);
  not i83447(x83447, x740);
  not i83448(x83448, x684);
  not i83449(x83449, x719);
  not i83450(x83450, x746);
  not i83451(x83451, x747);
  not i83452(x83452, x748);
  not i83453(x83453, x750);
  not i83454(x83454, x753);
  not i83455(x83455, x754);
  not i83456(x83456, x755);
  not i83457(x83457, x760);
  not i83458(x83458, x761);
  not i83459(x83459, x762);
  not i83460(x83460, x764);
  not i83461(x83461, x756);
  not i83462(x83462, x770);
  not i83463(x83463, x771);
  not i83464(x83464, x772);
  not i83465(x83465, x780);
  not i83466(x83466, x784);
  not i83467(x83467, x785);
  not i83468(x83468, x786);
  not i83469(x83469, x792);
  not i83470(x83470, x793);
  not i83471(x83471, x794);
  not i83472(x83472, x774);
  not i83473(x83473, x810);
  not i83474(x83474, x811);
  not i83475(x83475, x812);
  not i83476(x83476, x815);
  not i83477(x83477, x826);
  not i83478(x83478, x827);
  not i83479(x83479, x828);
  not i83480(x83480, x840);
  not i83481(x83481, x841);
  not i83482(x83482, x842);
  not i83483(x83483, x713);
  not i83484(x83484, x851);
  not i83485(x83485, x858);
  not i83486(x83486, x865);
  not i83487(x83487, x866);
  not i83488(x83488, x882);
  not i83489(x83489, x883);
  not i83490(x83490, x892);
  not i83491(x83491, x893);
  not i83492(x83492, x894);
  not i83493(x83493, x908);
  not i83494(x83494, x909);
  not i83495(x83495, x910);
  not i83496(x83496, x924);
  not i83497(x83497, x925);
  not i83498(x83498, x942);
  not i83499(x83499, x943);
  not i83500(x83500, x956);
  not i83501(x83501, x957);
  not i83502(x83502, x973);
  not i83503(x83503, x974);
  not i83504(x83504, x986);
  not i83505(x83505, x987);
  not i83506(x83506, x988);
  not i83507(x83507, x989);
  not i83508(x83508, x990);
  not i83509(x83509, x991);
  not i83510(x83510, x992);
  not i83511(x83511, x993);
  not i83512(x83512, x994);
  not i83513(x83513, x997);
  not i83514(x83514, x998);
  not i83515(x83515, x999);
  not i83516(x83516, x15984);
  not i83517(x83517, x15987);
  not i83518(x83518, x15991);
  not i83519(x83519, x15995);
  not i83520(x83520, x15999);
  not i83521(x83521, x16002);
  not i83522(x83522, x16006);
  not i83523(x83523, x16010);
  not i83524(x83524, x16014);
  not i83525(x83525, x16018);
  not i83526(x83526, x16022);
  not i83527(x83527, x16026);
  not i83528(x83528, x16030);
  not i83529(x83529, x16033);
  not i83530(x83530, x16037);
  not i83531(x83531, x16041);
  not i83532(x83532, x16045);
  not i83533(x83533, x16049);
  not i83534(x83534, x16053);
  not i83535(x83535, x16057);
  not i83536(x83536, x16061);
  not i83537(x83537, x16065);
  not i83538(x83538, x16069);
  not i83539(x83539, x16073);
  not i83540(x83540, x16077);
  not i83541(x83541, x16081);
  not i83542(x83542, x16085);
  not i83543(x83543, x16089);
  not i83544(x83544, x16093);
  not i83545(x83545, x16094);
  not i83546(x83546, x16149);
  not i83547(x83547, x16150);
  not i83548(x83548, x16201);
  not i83549(x83549, x16202);
  not i83550(x83550, x16203);
  not i83551(x83551, x16204);
  not i83552(x83552, x16247);
  not i83553(x83553, x16248);
  not i83554(x83554, x16249);
  not i83555(x83555, x16250);
  not i83556(x83556, x16251);
  not i83557(x83557, x16252);
  not i83558(x83558, x16253);
  not i83559(x83559, x16254);
  not i83560(x83560, x16281);
  not i83561(x83561, x16282);
  not i83562(x83562, x16283);
  not i83563(x83563, x16284);
  not i83564(x83564, x16285);
  not i83565(x83565, x16286);
  not i83566(x83566, x16287);
  not i83567(x83567, x16288);
  not i83568(x83568, x16289);
  not i83569(x83569, x16290);
  not i83570(x83570, x16291);
  not i83571(x83571, x16292);
  not i83572(x83572, x16293);
  not i83573(x83573, x15234);
  not i83574(x83574, x15976);
  not i83575(x83575, x18976);
  not i83576(x83576, x17956);
  not i83577(x83577, x19031);
  not i83578(x83578, x19029);
  not i83579(x83579, x18009);
  not i83580(x83580, x19112);
  not i83581(x83581, x19218);
  not i83582(x83582, x18169);
  not i83583(x83583, x19354);
  not i83584(x83584, x19352);
  not i83585(x83585, x18276);
  not i83586(x83586, x19516);
  not i83587(x83587, x19703);
  not i83588(x83588, x18544);
  not i83589(x83589, x19920);
  not i83590(x83590, x19918);
  not i83591(x83591, x18705);
  not i83592(x83592, x20163);
  not i83593(x83593, x18884);
  not i83594(x83594, x17921);
  not i83595(x83595, x18978);
  not i83596(x83596, x18993);
  not i83597(x83597, x20441);
  not i83598(x83598, x20449);
  not i83599(x83599, x20462);
  not i83600(x83600, x19110);
  not i83601(x83601, x20579);
  not i83602(x83602, x20576);
  not i83603(x83603, x20604);
  not i83604(x83604, x20600);
  not i83605(x83605, x20614);
  not i83606(x83606, x20632);
  not i83607(x83607, x20628);
  not i83608(x83608, x20642);
  not i83609(x83609, x20676);
  not i83610(x83610, x19514);
  not i83611(x83611, x19523);
  not i83612(x83612, x19585);
  not i83613(x83613, x18401);
  not i83614(x83614, x19647);
  not i83615(x83615, x19705);
  not i83616(x83616, x20909);
  not i83617(x83617, x20906);
  not i83618(x83618, x19712);
  not i83619(x83619, x19774);
  not i83620(x83620, x20955);
  not i83621(x83621, x20951);
  not i83622(x83622, x19782);
  not i83623(x83623, x20976);
  not i83624(x83624, x20974);
  not i83625(x83625, x21005);
  not i83626(x83626, x21001);
  not i83627(x83627, x19853);
  not i83628(x83628, x21026);
  not i83629(x83629, x21024);
  not i83630(x83630, x19927);
  not i83631(x83631, x21082);
  not i83632(x83632, x21080);
  not i83633(x83633, x20007);
  not i83634(x83634, x20087);
  not i83635(x83635, x20161);
  not i83636(x83636, x21245);
  not i83637(x83637, x21313);
  not i83638(x83638, x18949);
  not i83639(x83639, x18958);
  not i83640(x83640, x18966);
  not i83641(x83641, x18974);
  not i83642(x83642, x18985);
  not i83643(x83643, x20430);
  not i83644(x83644, x19001);
  not i83645(x83645, x20434);
  not i83646(x83646, x20439);
  not i83647(x83647, x20446);
  not i83648(x83648, x19018);
  not i83649(x83649, x20442);
  not i83650(x83650, x20447);
  not i83651(x83651, x20458);
  not i83652(x83652, x19038);
  not i83653(x83653, x20460);
  not i83654(x83654, x20472);
  not i83655(x83655, x19064);
  not i83656(x83656, x20492);
  not i83657(x83657, x19090);
  not i83658(x83658, x20512);
  not i83659(x83659, x19119);
  not i83660(x83660, x20532);
  not i83661(x83661, x19154);
  not i83662(x83662, x18080);
  not i83663(x83663, x20553);
  not i83664(x83664, x19189);
  not i83665(x83665, x19220);
  not i83666(x83666, x20574);
  not i83667(x83667, x19227);
  not i83668(x83668, x19262);
  not i83669(x83669, x21484);
  not i83670(x83670, x20598);
  not i83671(x83671, x21486);
  not i83672(x83672, x19270);
  not i83673(x83673, x20616);
  not i83674(x83674, x21497);
  not i83675(x83675, x21494);
  not i83676(x83676, x21499);
  not i83677(x83677, x20626);
  not i83678(x83678, x21503);
  not i83679(x83679, x19314);
  not i83680(x83680, x20644);
  not i83681(x83681, x21514);
  not i83682(x83682, x21511);
  not i83683(x83683, x21516);
  not i83684(x83684, x20654);
  not i83685(x83685, x21520);
  not i83686(x83686, x19361);
  not i83687(x83687, x20678);
  not i83688(x83688, x21532);
  not i83689(x83689, x21528);
  not i83690(x83690, x21534);
  not i83691(x83691, x20688);
  not i83692(x83692, x21538);
  not i83693(x83693, x19414);
  not i83694(x83694, x20717);
  not i83695(x83695, x21550);
  not i83696(x83696, x21546);
  not i83697(x83697, x21552);
  not i83698(x83698, x20728);
  not i83699(x83699, x21557);
  not i83700(x83700, x19467);
  not i83701(x83701, x20757);
  not i83702(x83702, x21569);
  not i83703(x83703, x21565);
  not i83704(x83704, x21571);
  not i83705(x83705, x20768);
  not i83706(x83706, x21576);
  not i83707(x83707, x20797);
  not i83708(x83708, x21593);
  not i83709(x83709, x21589);
  not i83710(x83710, x21595);
  not i83711(x83711, x20808);
  not i83712(x83712, x21600);
  not i83713(x83713, x21615);
  not i83714(x83714, x21613);
  not i83715(x83715, x21620);
  not i83716(x83716, x21616);
  not i83717(x83717, x21622);
  not i83718(x83718, x20850);
  not i83719(x83719, x21627);
  not i83720(x83720, x21642);
  not i83721(x83721, x21640);
  not i83722(x83722, x21647);
  not i83723(x83723, x21643);
  not i83724(x83724, x21649);
  not i83725(x83725, x20892);
  not i83726(x83726, x21654);
  not i83727(x83727, x21669);
  not i83728(x83728, x21667);
  not i83729(x83729, x21682);
  not i83730(x83730, x20937);
  not i83731(x83731, x21687);
  not i83732(x83732, x21702);
  not i83733(x83733, x21700);
  not i83734(x83734, x21715);
  not i83735(x83735, x21740);
  not i83736(x83736, x21738);
  not i83737(x83737, x21753);
  not i83738(x83738, x21778);
  not i83739(x83739, x21776);
  not i83740(x83740, x21792);
  not i83741(x83741, x21817);
  not i83742(x83742, x21815);
  not i83743(x83743, x21831);
  not i83744(x83744, x21857);
  not i83745(x83745, x21855);
  not i83746(x83746, x21871);
  not i83747(x83747, x21897);
  not i83748(x83748, x21895);
  not i83749(x83749, x20433);
  not i83750(x83750, x21414);
  not i83751(x83751, x20438);
  not i83752(x83752, x22012);
  not i83753(x83753, x21418);
  not i83754(x83754, x21422);
  not i83755(x83755, x21426);
  not i83756(x83756, x21431);
  not i83757(x83757, x21437);
  not i83758(x83758, x21443);
  not i83759(x83759, x21447);
  not i83760(x83760, x21453);
  not i83761(x83761, x21457);
  not i83762(x83762, x21463);
  not i83763(x83763, x21467);
  not i83764(x83764, x21473);
  not i83765(x83765, x21477);
  not i83766(x83766, x21481);
  not i83767(x83767, x22128);
  not i83768(x83768, x21490);
  not i83769(x83769, x22132);
  not i83770(x83770, x21507);
  not i83771(x83771, x22154);
  not i83772(x83772, x21524);
  not i83773(x83773, x22176);
  not i83774(x83774, x21542);
  not i83775(x83775, x22198);
  not i83776(x83776, x21561);
  not i83777(x83777, x22220);
  not i83778(x83778, x22243);
  not i83779(x83779, x21406);
  not i83780(x83780, x22001);
  not i83781(x83781, x21410);
  not i83782(x83782, x22005);
  not i83783(x83783, x22011);
  not i83784(x83784, x22009);
  not i83785(x83785, x22557);
  not i83786(x83786, x22018);
  not i83787(x83787, x22561);
  not i83788(x83788, x22016);
  not i83789(x83789, x22564);
  not i83790(x83790, x22030);
  not i83791(x83791, x22569);
  not i83792(x83792, x22028);
  not i83793(x83793, x22572);
  not i83794(x83794, x22042);
  not i83795(x83795, x22577);
  not i83796(x83796, x22040);
  not i83797(x83797, x22580);
  not i83798(x83798, x22054);
  not i83799(x83799, x22585);
  not i83800(x83800, x22052);
  not i83801(x83801, x22588);
  not i83802(x83802, x22066);
  not i83803(x83803, x22593);
  not i83804(x83804, x22064);
  not i83805(x83805, x22596);
  not i83806(x83806, x22076);
  not i83807(x83807, x22610);
  not i83808(x83808, x22089);
  not i83809(x83809, x22624);
  not i83810(x83810, x22102);
  not i83811(x83811, x22638);
  not i83812(x83812, x22115);
  not i83813(x83813, x22652);
  not i83814(x83814, x22000);
  not i83815(x83815, x22550);
  not i83816(x83816, x22548);
  not i83817(x83817, x22553);
  not i83818(x83818, x22551);
  not i83819(x83819, x22556);
  not i83820(x83820, x22554);
  not i83821(x83821, x22563);
  not i83822(x83822, x22571);
  not i83823(x83823, x22579);
  not i83824(x83824, x22587);
  not i83825(x83825, x22595);
  not i83826(x83826, x21995);
  not i83827(x83827, x23330);
  not i83828(x83828, x21998);
  not i83829(x83829, x22972);
  not i83830(x83830, x23333);
  not i83831(x83831, x22975);
  not i83832(x83832, x23336);
  not i83833(x83833, x22979);
  not i83834(x83834, x23340);
  not i83835(x83835, x23345);
  not i83836(x83836, x23350);
  not i83837(x83837, x23355);
  not i83838(x83838, x23360);
  not i83839(x83839, x22974);
  not i83840(x83840, x23561);
  not i83841(x83841, x23335);
  not i83842(x83842, x23565);
  not i83843(x83843, x18951);
  not i83844(x83844, x21997);
  not i83845(x83845, x23332);
  not i83846(x83846, x23559);
  not i83847(x83847, x23814);
  not i83848(x83848, x24576);
  not i83849(x83849, x24633);
  not i83850(x83850, x24634);
  not i83851(x83851, x24635);
  not i83852(x83852, x24684);
  not i83853(x83853, x24685);
  not i83854(x83854, x24686);
  not i83855(x83855, x24687);
  not i83856(x83856, x24688);
  not i83857(x83857, x24689);
  not i83858(x83858, x24690);
  not i83859(x83859, x24691);
  not i83860(x83860, x24722);
  not i83861(x83861, x24723);
  not i83862(x83862, x24724);
  not i83863(x83863, x24725);
  not i83864(x83864, x24726);
  not i83865(x83865, x24727);
  not i83866(x83866, x24728);
  not i83867(x83867, x24729);
  not i83868(x83868, x24730);
  not i83869(x83869, x24731);
  not i83870(x83870, x24732);
  not i83871(x83871, x24733);
  not i83872(x83872, x24734);
  not i83873(x83873, x24735);
  not i83874(x83874, x24736);
  not i83875(x83875, x24989);
  not i83876(x83876, x25052);
  not i83877(x83877, x25053);
  not i83878(x83878, x25144);
  not i83879(x83879, x25145);
  not i83880(x83880, x25146);
  not i83881(x83881, x25147);
  not i83882(x83882, x25232);
  not i83883(x83883, x25233);
  not i83884(x83884, x25234);
  not i83885(x83885, x25235);
  not i83886(x83886, x25236);
  not i83887(x83887, x25237);
  not i83888(x83888, x25238);
  not i83889(x83889, x25239);
  not i83890(x83890, x25312);
  not i83891(x83891, x25313);
  not i83892(x83892, x25314);
  not i83893(x83893, x25315);
  not i83894(x83894, x25316);
  not i83895(x83895, x25317);
  not i83896(x83896, x25318);
  not i83897(x83897, x25319);
  not i83898(x83898, x25320);
  not i83899(x83899, x25321);
  not i83900(x83900, x25322);
  not i83901(x83901, x25323);
  not i83902(x83902, x25324);
  not i83903(x83903, x25325);
  not i83904(x83904, x25326);
  not i83905(x83905, x25327);
  not i83906(x83906, x25050);
  not i83907(x83907, x25497);
  not i83908(x83908, x25498);
  not i83909(x83909, x25583);
  not i83910(x83910, x25584);
  not i83911(x83911, x25585);
  not i83912(x83912, x25586);
  not i83913(x83913, x25659);
  not i83914(x83914, x25660);
  not i83915(x83915, x25661);
  not i83916(x83916, x25662);
  not i83917(x83917, x25663);
  not i83918(x83918, x25664);
  not i83919(x83919, x25665);
  not i83920(x83920, x25666);
  not i83921(x83921, x25715);
  not i83922(x83922, x25716);
  not i83923(x83923, x25717);
  not i83924(x83924, x25718);
  not i83925(x83925, x25719);
  not i83926(x83926, x25720);
  not i83927(x83927, x25721);
  not i83928(x83928, x25722);
  not i83929(x83929, x25723);
  not i83930(x83930, x25724);
  not i83931(x83931, x25725);
  not i83932(x83932, x25726);
  not i83933(x83933, x25727);
  not i83934(x83934, x25728);
  not i83935(x83935, x25729);
  not i83936(x83936, x25730);
  not i83937(x83937, x25731);
  not i83938(x83938, x25732);
  not i83939(x83939, x25736);
  not i83940(x83940, x25737);
  not i83941(x83941, x25748);
  not i83942(x83942, x25750);
  not i83943(x83943, x25751);
  not i83944(x83944, x25770);
  not i83945(x83945, x25781);
  not i83946(x83946, x25783);
  not i83947(x83947, x25791);
  not i83948(x83948, x25799);
  not i83949(x83949, x25800);
  not i83950(x83950, x25804);
  not i83951(x83951, x25805);
  not i83952(x83952, x25816);
  not i83953(x83953, x25817);
  not i83954(x83954, x25818);
  not i83955(x83955, x25837);
  not i83956(x83956, x25847);
  not i83957(x83957, x25848);
  not i83958(x83958, x25855);
  not i83959(x83959, x25862);
  not i83960(x83960, x25863);
  not i83961(x83961, x25867);
  not i83962(x83962, x25868);
  not i83963(x83963, x25879);
  not i83964(x83964, x25880);
  not i83965(x83965, x25881);
  not i83966(x83966, x25900);
  not i83967(x83967, x25910);
  not i83968(x83968, x25911);
  not i83969(x83969, x25918);
  not i83970(x83970, x25925);
  not i83971(x83971, x25926);
  not i83972(x83972, x25930);
  not i83973(x83973, x25931);
  not i83974(x83974, x25942);
  not i83975(x83975, x25943);
  not i83976(x83976, x25944);
  not i83977(x83977, x25963);
  not i83978(x83978, x25973);
  not i83979(x83979, x25974);
  not i83980(x83980, x25981);
  not i83981(x83981, x25988);
  not i83982(x83982, x25989);
  not i83983(x83983, x25993);
  not i83984(x83984, x25994);
  not i83985(x83985, x26005);
  not i83986(x83986, x26006);
  not i83987(x83987, x26007);
  not i83988(x83988, x26026);
  not i83989(x83989, x26036);
  not i83990(x83990, x26037);
  not i83991(x83991, x26044);
  not i83992(x83992, x26051);
  not i83993(x83993, x26052);
  not i83994(x83994, x26056);
  not i83995(x83995, x26057);
  not i83996(x83996, x26068);
  not i83997(x83997, x26069);
  not i83998(x83998, x26070);
  not i83999(x83999, x26089);
  not i84000(x84000, x26099);
  not i84001(x84001, x26100);
  not i84002(x84002, x26107);
  not i84003(x84003, x26114);
  not i84004(x84004, x26115);
  not i84005(x84005, x26119);
  not i84006(x84006, x26120);
  not i84007(x84007, x26131);
  not i84008(x84008, x26132);
  not i84009(x84009, x26133);
  not i84010(x84010, x26152);
  not i84011(x84011, x26162);
  not i84012(x84012, x26163);
  not i84013(x84013, x26170);
  not i84014(x84014, x26177);
  not i84015(x84015, x26178);
  not i84016(x84016, x26182);
  not i84017(x84017, x26183);
  not i84018(x84018, x26194);
  not i84019(x84019, x26195);
  not i84020(x84020, x26196);
  not i84021(x84021, x26215);
  not i84022(x84022, x26225);
  not i84023(x84023, x26226);
  not i84024(x84024, x26233);
  not i84025(x84025, x26240);
  not i84026(x84026, x26241);
  not i84027(x84027, x26245);
  not i84028(x84028, x26246);
  not i84029(x84029, x26257);
  not i84030(x84030, x26258);
  not i84031(x84031, x26259);
  not i84032(x84032, x26278);
  not i84033(x84033, x26288);
  not i84034(x84034, x26289);
  not i84035(x84035, x26296);
  not i84036(x84036, x26303);
  not i84037(x84037, x26304);
  not i84038(x84038, x26308);
  not i84039(x84039, x26309);
  not i84040(x84040, x26320);
  not i84041(x84041, x26321);
  not i84042(x84042, x26322);
  not i84043(x84043, x26341);
  not i84044(x84044, x26351);
  not i84045(x84045, x26352);
  not i84046(x84046, x26359);
  not i84047(x84047, x26366);
  not i84048(x84048, x26367);
  not i84049(x84049, x26371);
  not i84050(x84050, x26372);
  not i84051(x84051, x26383);
  not i84052(x84052, x26384);
  not i84053(x84053, x26385);
  not i84054(x84054, x26404);
  not i84055(x84055, x26414);
  not i84056(x84056, x26415);
  not i84057(x84057, x26422);
  not i84058(x84058, x26429);
  not i84059(x84059, x26430);
  not i84060(x84060, x26434);
  not i84061(x84061, x26435);
  not i84062(x84062, x26446);
  not i84063(x84063, x26447);
  not i84064(x84064, x26448);
  not i84065(x84065, x26467);
  not i84066(x84066, x26477);
  not i84067(x84067, x26478);
  not i84068(x84068, x26485);
  not i84069(x84069, x26492);
  not i84070(x84070, x26493);
  not i84071(x84071, x26497);
  not i84072(x84072, x26498);
  not i84073(x84073, x26509);
  not i84074(x84074, x26510);
  not i84075(x84075, x26511);
  not i84076(x84076, x26530);
  not i84077(x84077, x26540);
  not i84078(x84078, x26541);
  not i84079(x84079, x26548);
  not i84080(x84080, x26555);
  not i84081(x84081, x26556);
  not i84082(x84082, x26560);
  not i84083(x84083, x26561);
  not i84084(x84084, x26572);
  not i84085(x84085, x26573);
  not i84086(x84086, x26574);
  not i84087(x84087, x26593);
  not i84088(x84088, x26603);
  not i84089(x84089, x26604);
  not i84090(x84090, x26611);
  not i84091(x84091, x26618);
  not i84092(x84092, x26619);
  not i84093(x84093, x26623);
  not i84094(x84094, x26624);
  not i84095(x84095, x26635);
  not i84096(x84096, x26636);
  not i84097(x84097, x26637);
  not i84098(x84098, x26656);
  not i84099(x84099, x26666);
  not i84100(x84100, x26667);
  not i84101(x84101, x26674);
  not i84102(x84102, x26681);
  not i84103(x84103, x26682);
  not i84104(x84104, x26686);
  not i84105(x84105, x26687);
  not i84106(x84106, x26698);
  not i84107(x84107, x26699);
  not i84108(x84108, x26700);
  not i84109(x84109, x26719);
  not i84110(x84110, x26729);
  not i84111(x84111, x26730);
  not i84112(x84112, x26737);
  not i84113(x84113, x26744);
  not i84114(x84114, x26745);
  not i84115(x84115, x26749);
  not i84116(x84116, x26750);
  not i84117(x84117, x26761);
  not i84118(x84118, x26762);
  not i84119(x84119, x26763);
  not i84120(x84120, x26782);
  not i84121(x84121, x26792);
  not i84122(x84122, x26793);
  not i84123(x84123, x26800);
  not i84124(x84124, x26807);
  not i84125(x84125, x26808);
  not i84126(x84126, x26812);
  not i84127(x84127, x26813);
  not i84128(x84128, x26824);
  not i84129(x84129, x26825);
  not i84130(x84130, x26826);
  not i84131(x84131, x26845);
  not i84132(x84132, x26855);
  not i84133(x84133, x26856);
  not i84134(x84134, x26863);
  not i84135(x84135, x26870);
  not i84136(x84136, x26871);
  not i84137(x84137, x26875);
  not i84138(x84138, x26876);
  not i84139(x84139, x26887);
  not i84140(x84140, x26888);
  not i84141(x84141, x26889);
  not i84142(x84142, x26908);
  not i84143(x84143, x26918);
  not i84144(x84144, x26919);
  not i84145(x84145, x26926);
  not i84146(x84146, x26933);
  not i84147(x84147, x26934);
  not i84148(x84148, x26938);
  not i84149(x84149, x26939);
  not i84150(x84150, x26950);
  not i84151(x84151, x26951);
  not i84152(x84152, x26952);
  not i84153(x84153, x26971);
  not i84154(x84154, x26981);
  not i84155(x84155, x26982);
  not i84156(x84156, x26989);
  not i84157(x84157, x26996);
  not i84158(x84158, x26997);
  not i84159(x84159, x27001);
  not i84160(x84160, x27002);
  not i84161(x84161, x27013);
  not i84162(x84162, x27014);
  not i84163(x84163, x27015);
  not i84164(x84164, x27034);
  not i84165(x84165, x27044);
  not i84166(x84166, x27045);
  not i84167(x84167, x27052);
  not i84168(x84168, x27059);
  not i84169(x84169, x27060);
  not i84170(x84170, x27064);
  not i84171(x84171, x27065);
  not i84172(x84172, x27076);
  not i84173(x84173, x27077);
  not i84174(x84174, x27078);
  not i84175(x84175, x27097);
  not i84176(x84176, x27107);
  not i84177(x84177, x27108);
  not i84178(x84178, x27115);
  not i84179(x84179, x27122);
  not i84180(x84180, x27123);
  not i84181(x84181, x27127);
  not i84182(x84182, x27128);
  not i84183(x84183, x27139);
  not i84184(x84184, x27140);
  not i84185(x84185, x27141);
  not i84186(x84186, x27160);
  not i84187(x84187, x27170);
  not i84188(x84188, x27171);
  not i84189(x84189, x27178);
  not i84190(x84190, x27185);
  not i84191(x84191, x27186);
  not i84192(x84192, x27190);
  not i84193(x84193, x27191);
  not i84194(x84194, x27202);
  not i84195(x84195, x27203);
  not i84196(x84196, x27204);
  not i84197(x84197, x27223);
  not i84198(x84198, x27233);
  not i84199(x84199, x27234);
  not i84200(x84200, x27241);
  not i84201(x84201, x27248);
  not i84202(x84202, x27249);
  not i84203(x84203, x27253);
  not i84204(x84204, x27254);
  not i84205(x84205, x27265);
  not i84206(x84206, x27266);
  not i84207(x84207, x27267);
  not i84208(x84208, x27286);
  not i84209(x84209, x27296);
  not i84210(x84210, x27297);
  not i84211(x84211, x27304);
  not i84212(x84212, x27311);
  not i84213(x84213, x27312);
  not i84214(x84214, x27316);
  not i84215(x84215, x27317);
  not i84216(x84216, x27328);
  not i84217(x84217, x27329);
  not i84218(x84218, x27330);
  not i84219(x84219, x27349);
  not i84220(x84220, x27359);
  not i84221(x84221, x27360);
  not i84222(x84222, x27367);
  not i84223(x84223, x27374);
  not i84224(x84224, x27375);
  not i84225(x84225, x27379);
  not i84226(x84226, x27380);
  not i84227(x84227, x27391);
  not i84228(x84228, x27392);
  not i84229(x84229, x27393);
  not i84230(x84230, x27412);
  not i84231(x84231, x27422);
  not i84232(x84232, x27423);
  not i84233(x84233, x27430);
  not i84234(x84234, x27437);
  not i84235(x84235, x27438);
  not i84236(x84236, x27442);
  not i84237(x84237, x27443);
  not i84238(x84238, x27454);
  not i84239(x84239, x27455);
  not i84240(x84240, x27456);
  not i84241(x84241, x27475);
  not i84242(x84242, x27485);
  not i84243(x84243, x27486);
  not i84244(x84244, x27493);
  not i84245(x84245, x27500);
  not i84246(x84246, x27501);
  not i84247(x84247, x27505);
  not i84248(x84248, x27506);
  not i84249(x84249, x27517);
  not i84250(x84250, x27518);
  not i84251(x84251, x27519);
  not i84252(x84252, x27538);
  not i84253(x84253, x27548);
  not i84254(x84254, x27549);
  not i84255(x84255, x27556);
  not i84256(x84256, x27563);
  not i84257(x84257, x27564);
  not i84258(x84258, x27568);
  not i84259(x84259, x27569);
  not i84260(x84260, x27580);
  not i84261(x84261, x27581);
  not i84262(x84262, x27582);
  not i84263(x84263, x27601);
  not i84264(x84264, x27611);
  not i84265(x84265, x27612);
  not i84266(x84266, x27619);
  not i84267(x84267, x27626);
  not i84268(x84268, x27627);
  not i84269(x84269, x27631);
  not i84270(x84270, x27632);
  not i84271(x84271, x27643);
  not i84272(x84272, x27644);
  not i84273(x84273, x27645);
  not i84274(x84274, x27664);
  not i84275(x84275, x27674);
  not i84276(x84276, x27675);
  not i84277(x84277, x27682);
  not i84278(x84278, x27689);
  not i84279(x84279, x27690);
  not i84280(x84280, x27694);
  not i84281(x84281, x27695);
  not i84282(x84282, x27706);
  not i84283(x84283, x27707);
  not i84284(x84284, x27708);
  not i84285(x84285, x27727);
  not i84286(x84286, x27737);
  not i84287(x84287, x27738);
  not i84288(x84288, x27745);
  not i84289(x84289, x30076);
  not i84290(x84290, x29056);
  not i84291(x84291, x30131);
  not i84292(x84292, x30129);
  not i84293(x84293, x29109);
  not i84294(x84294, x30212);
  not i84295(x84295, x30318);
  not i84296(x84296, x29269);
  not i84297(x84297, x30454);
  not i84298(x84298, x30452);
  not i84299(x84299, x29376);
  not i84300(x84300, x30616);
  not i84301(x84301, x30803);
  not i84302(x84302, x29644);
  not i84303(x84303, x31020);
  not i84304(x84304, x31018);
  not i84305(x84305, x29805);
  not i84306(x84306, x31263);
  not i84307(x84307, x29984);
  not i84308(x84308, x29021);
  not i84309(x84309, x30078);
  not i84310(x84310, x30093);
  not i84311(x84311, x31541);
  not i84312(x84312, x31549);
  not i84313(x84313, x31562);
  not i84314(x84314, x30210);
  not i84315(x84315, x31679);
  not i84316(x84316, x31676);
  not i84317(x84317, x31704);
  not i84318(x84318, x31700);
  not i84319(x84319, x31714);
  not i84320(x84320, x31732);
  not i84321(x84321, x31728);
  not i84322(x84322, x31742);
  not i84323(x84323, x31776);
  not i84324(x84324, x30614);
  not i84325(x84325, x30623);
  not i84326(x84326, x30685);
  not i84327(x84327, x29501);
  not i84328(x84328, x30747);
  not i84329(x84329, x30805);
  not i84330(x84330, x32009);
  not i84331(x84331, x32006);
  not i84332(x84332, x30812);
  not i84333(x84333, x30874);
  not i84334(x84334, x32055);
  not i84335(x84335, x32051);
  not i84336(x84336, x30882);
  not i84337(x84337, x32076);
  not i84338(x84338, x32074);
  not i84339(x84339, x32105);
  not i84340(x84340, x32101);
  not i84341(x84341, x30953);
  not i84342(x84342, x32126);
  not i84343(x84343, x32124);
  not i84344(x84344, x31027);
  not i84345(x84345, x32182);
  not i84346(x84346, x32180);
  not i84347(x84347, x31107);
  not i84348(x84348, x31187);
  not i84349(x84349, x31261);
  not i84350(x84350, x32345);
  not i84351(x84351, x32413);
  not i84352(x84352, x30049);
  not i84353(x84353, x30058);
  not i84354(x84354, x30066);
  not i84355(x84355, x30074);
  not i84356(x84356, x30085);
  not i84357(x84357, x31530);
  not i84358(x84358, x30101);
  not i84359(x84359, x31534);
  not i84360(x84360, x31539);
  not i84361(x84361, x31546);
  not i84362(x84362, x30118);
  not i84363(x84363, x31542);
  not i84364(x84364, x31547);
  not i84365(x84365, x31558);
  not i84366(x84366, x30138);
  not i84367(x84367, x31560);
  not i84368(x84368, x31572);
  not i84369(x84369, x30164);
  not i84370(x84370, x31592);
  not i84371(x84371, x30190);
  not i84372(x84372, x31612);
  not i84373(x84373, x30219);
  not i84374(x84374, x31632);
  not i84375(x84375, x30254);
  not i84376(x84376, x29180);
  not i84377(x84377, x31653);
  not i84378(x84378, x30289);
  not i84379(x84379, x30320);
  not i84380(x84380, x31674);
  not i84381(x84381, x30327);
  not i84382(x84382, x30362);
  not i84383(x84383, x32584);
  not i84384(x84384, x31698);
  not i84385(x84385, x32586);
  not i84386(x84386, x30370);
  not i84387(x84387, x31716);
  not i84388(x84388, x32597);
  not i84389(x84389, x32594);
  not i84390(x84390, x32599);
  not i84391(x84391, x31726);
  not i84392(x84392, x32603);
  not i84393(x84393, x30414);
  not i84394(x84394, x31744);
  not i84395(x84395, x32614);
  not i84396(x84396, x32611);
  not i84397(x84397, x32616);
  not i84398(x84398, x31754);
  not i84399(x84399, x32620);
  not i84400(x84400, x30461);
  not i84401(x84401, x31778);
  not i84402(x84402, x32632);
  not i84403(x84403, x32628);
  not i84404(x84404, x32634);
  not i84405(x84405, x31788);
  not i84406(x84406, x32638);
  not i84407(x84407, x30514);
  not i84408(x84408, x31817);
  not i84409(x84409, x32650);
  not i84410(x84410, x32646);
  not i84411(x84411, x32652);
  not i84412(x84412, x31828);
  not i84413(x84413, x32657);
  not i84414(x84414, x30567);
  not i84415(x84415, x31857);
  not i84416(x84416, x32669);
  not i84417(x84417, x32665);
  not i84418(x84418, x32671);
  not i84419(x84419, x31868);
  not i84420(x84420, x32676);
  not i84421(x84421, x31897);
  not i84422(x84422, x32693);
  not i84423(x84423, x32689);
  not i84424(x84424, x32695);
  not i84425(x84425, x31908);
  not i84426(x84426, x32700);
  not i84427(x84427, x32715);
  not i84428(x84428, x32713);
  not i84429(x84429, x32720);
  not i84430(x84430, x32716);
  not i84431(x84431, x32722);
  not i84432(x84432, x31950);
  not i84433(x84433, x32727);
  not i84434(x84434, x32742);
  not i84435(x84435, x32740);
  not i84436(x84436, x32747);
  not i84437(x84437, x32743);
  not i84438(x84438, x32749);
  not i84439(x84439, x31992);
  not i84440(x84440, x32754);
  not i84441(x84441, x32769);
  not i84442(x84442, x32767);
  not i84443(x84443, x32782);
  not i84444(x84444, x32037);
  not i84445(x84445, x32787);
  not i84446(x84446, x32802);
  not i84447(x84447, x32800);
  not i84448(x84448, x32815);
  not i84449(x84449, x32840);
  not i84450(x84450, x32838);
  not i84451(x84451, x32853);
  not i84452(x84452, x32878);
  not i84453(x84453, x32876);
  not i84454(x84454, x32892);
  not i84455(x84455, x32917);
  not i84456(x84456, x32915);
  not i84457(x84457, x32931);
  not i84458(x84458, x32957);
  not i84459(x84459, x32955);
  not i84460(x84460, x32971);
  not i84461(x84461, x32997);
  not i84462(x84462, x32995);
  not i84463(x84463, x31533);
  not i84464(x84464, x32514);
  not i84465(x84465, x31538);
  not i84466(x84466, x33112);
  not i84467(x84467, x32518);
  not i84468(x84468, x32522);
  not i84469(x84469, x32526);
  not i84470(x84470, x32531);
  not i84471(x84471, x32537);
  not i84472(x84472, x32543);
  not i84473(x84473, x32547);
  not i84474(x84474, x32553);
  not i84475(x84475, x32557);
  not i84476(x84476, x32563);
  not i84477(x84477, x32567);
  not i84478(x84478, x32573);
  not i84479(x84479, x32577);
  not i84480(x84480, x32581);
  not i84481(x84481, x33228);
  not i84482(x84482, x32590);
  not i84483(x84483, x33232);
  not i84484(x84484, x32607);
  not i84485(x84485, x33254);
  not i84486(x84486, x32624);
  not i84487(x84487, x33276);
  not i84488(x84488, x32642);
  not i84489(x84489, x33298);
  not i84490(x84490, x32661);
  not i84491(x84491, x33320);
  not i84492(x84492, x33343);
  not i84493(x84493, x32506);
  not i84494(x84494, x33101);
  not i84495(x84495, x32510);
  not i84496(x84496, x33105);
  not i84497(x84497, x33111);
  not i84498(x84498, x33109);
  not i84499(x84499, x33657);
  not i84500(x84500, x33118);
  not i84501(x84501, x33661);
  not i84502(x84502, x33116);
  not i84503(x84503, x33664);
  not i84504(x84504, x33130);
  not i84505(x84505, x33669);
  not i84506(x84506, x33128);
  not i84507(x84507, x33672);
  not i84508(x84508, x33142);
  not i84509(x84509, x33677);
  not i84510(x84510, x33140);
  not i84511(x84511, x33680);
  not i84512(x84512, x33154);
  not i84513(x84513, x33685);
  not i84514(x84514, x33152);
  not i84515(x84515, x33688);
  not i84516(x84516, x33166);
  not i84517(x84517, x33693);
  not i84518(x84518, x33164);
  not i84519(x84519, x33696);
  not i84520(x84520, x33176);
  not i84521(x84521, x33710);
  not i84522(x84522, x33189);
  not i84523(x84523, x33724);
  not i84524(x84524, x33202);
  not i84525(x84525, x33738);
  not i84526(x84526, x33215);
  not i84527(x84527, x33752);
  not i84528(x84528, x33100);
  not i84529(x84529, x33650);
  not i84530(x84530, x33648);
  not i84531(x84531, x33653);
  not i84532(x84532, x33651);
  not i84533(x84533, x33656);
  not i84534(x84534, x33654);
  not i84535(x84535, x33663);
  not i84536(x84536, x33671);
  not i84537(x84537, x33679);
  not i84538(x84538, x33687);
  not i84539(x84539, x33695);
  not i84540(x84540, x33095);
  not i84541(x84541, x34430);
  not i84542(x84542, x33098);
  not i84543(x84543, x34072);
  not i84544(x84544, x34433);
  not i84545(x84545, x34075);
  not i84546(x84546, x34436);
  not i84547(x84547, x34079);
  not i84548(x84548, x34440);
  not i84549(x84549, x34445);
  not i84550(x84550, x34450);
  not i84551(x84551, x34455);
  not i84552(x84552, x34460);
  not i84553(x84553, x34074);
  not i84554(x84554, x34661);
  not i84555(x84555, x34435);
  not i84556(x84556, x34665);
  not i84557(x84557, x30051);
  not i84558(x84558, x33097);
  not i84559(x84559, x34432);
  not i84560(x84560, x34659);
  not i84561(x84561, x34914);
  not i84562(x84562, x35676);
  not i84563(x84563, x35733);
  not i84564(x84564, x35734);
  not i84565(x84565, x35735);
  not i84566(x84566, x35784);
  not i84567(x84567, x35785);
  not i84568(x84568, x35786);
  not i84569(x84569, x35787);
  not i84570(x84570, x35788);
  not i84571(x84571, x35789);
  not i84572(x84572, x35790);
  not i84573(x84573, x35791);
  not i84574(x84574, x35822);
  not i84575(x84575, x35823);
  not i84576(x84576, x35824);
  not i84577(x84577, x35825);
  not i84578(x84578, x35826);
  not i84579(x84579, x35827);
  not i84580(x84580, x35828);
  not i84581(x84581, x35829);
  not i84582(x84582, x35830);
  not i84583(x84583, x35831);
  not i84584(x84584, x35832);
  not i84585(x84585, x35833);
  not i84586(x84586, x35834);
  not i84587(x84587, x35835);
  not i84588(x84588, x35836);
  not i84589(x84589, x36089);
  not i84590(x84590, x36152);
  not i84591(x84591, x36153);
  not i84592(x84592, x36244);
  not i84593(x84593, x36245);
  not i84594(x84594, x36246);
  not i84595(x84595, x36247);
  not i84596(x84596, x36332);
  not i84597(x84597, x36333);
  not i84598(x84598, x36334);
  not i84599(x84599, x36335);
  not i84600(x84600, x36336);
  not i84601(x84601, x36337);
  not i84602(x84602, x36338);
  not i84603(x84603, x36339);
  not i84604(x84604, x36412);
  not i84605(x84605, x36413);
  not i84606(x84606, x36414);
  not i84607(x84607, x36415);
  not i84608(x84608, x36416);
  not i84609(x84609, x36417);
  not i84610(x84610, x36418);
  not i84611(x84611, x36419);
  not i84612(x84612, x36420);
  not i84613(x84613, x36421);
  not i84614(x84614, x36422);
  not i84615(x84615, x36423);
  not i84616(x84616, x36424);
  not i84617(x84617, x36425);
  not i84618(x84618, x36426);
  not i84619(x84619, x36427);
  not i84620(x84620, x36150);
  not i84621(x84621, x36597);
  not i84622(x84622, x36598);
  not i84623(x84623, x36683);
  not i84624(x84624, x36684);
  not i84625(x84625, x36685);
  not i84626(x84626, x36686);
  not i84627(x84627, x36759);
  not i84628(x84628, x36760);
  not i84629(x84629, x36761);
  not i84630(x84630, x36762);
  not i84631(x84631, x36763);
  not i84632(x84632, x36764);
  not i84633(x84633, x36765);
  not i84634(x84634, x36766);
  not i84635(x84635, x36815);
  not i84636(x84636, x36816);
  not i84637(x84637, x36817);
  not i84638(x84638, x36818);
  not i84639(x84639, x36819);
  not i84640(x84640, x36820);
  not i84641(x84641, x36821);
  not i84642(x84642, x36822);
  not i84643(x84643, x36823);
  not i84644(x84644, x36824);
  not i84645(x84645, x36825);
  not i84646(x84646, x36826);
  not i84647(x84647, x36827);
  not i84648(x84648, x36828);
  not i84649(x84649, x36829);
  not i84650(x84650, x36830);
  not i84651(x84651, x36831);
  not i84652(x84652, x36834);
  not i84653(x84653, x36835);
  not i84654(x84654, x36846);
  not i84655(x84655, x36847);
  not i84656(x84656, x36866);
  not i84657(x84657, x36875);
  not i84658(x84658, x36876);
  not i84659(x84659, x36883);
  not i84660(x84660, x36890);
  not i84661(x84661, x36893);
  not i84662(x84662, x36894);
  not i84663(x84663, x36905);
  not i84664(x84664, x36906);
  not i84665(x84665, x36925);
  not i84666(x84666, x36934);
  not i84667(x84667, x36935);
  not i84668(x84668, x36942);
  not i84669(x84669, x36949);
  not i84670(x84670, x36952);
  not i84671(x84671, x36953);
  not i84672(x84672, x36964);
  not i84673(x84673, x36965);
  not i84674(x84674, x36984);
  not i84675(x84675, x36993);
  not i84676(x84676, x36994);
  not i84677(x84677, x37001);
  not i84678(x84678, x37008);
  not i84679(x84679, x37011);
  not i84680(x84680, x37012);
  not i84681(x84681, x37023);
  not i84682(x84682, x37024);
  not i84683(x84683, x37043);
  not i84684(x84684, x37052);
  not i84685(x84685, x37053);
  not i84686(x84686, x37060);
  not i84687(x84687, x37067);
  not i84688(x84688, x37070);
  not i84689(x84689, x37071);
  not i84690(x84690, x37082);
  not i84691(x84691, x37083);
  not i84692(x84692, x37102);
  not i84693(x84693, x37111);
  not i84694(x84694, x37112);
  not i84695(x84695, x37119);
  not i84696(x84696, x37126);
  not i84697(x84697, x37129);
  not i84698(x84698, x37130);
  not i84699(x84699, x37141);
  not i84700(x84700, x37142);
  not i84701(x84701, x37161);
  not i84702(x84702, x37170);
  not i84703(x84703, x37171);
  not i84704(x84704, x37178);
  not i84705(x84705, x37185);
  not i84706(x84706, x37188);
  not i84707(x84707, x37189);
  not i84708(x84708, x37200);
  not i84709(x84709, x37201);
  not i84710(x84710, x37220);
  not i84711(x84711, x37229);
  not i84712(x84712, x37230);
  not i84713(x84713, x37237);
  not i84714(x84714, x37244);
  not i84715(x84715, x37247);
  not i84716(x84716, x37248);
  not i84717(x84717, x37259);
  not i84718(x84718, x37260);
  not i84719(x84719, x37279);
  not i84720(x84720, x37288);
  not i84721(x84721, x37289);
  not i84722(x84722, x37296);
  not i84723(x84723, x37303);
  not i84724(x84724, x37306);
  not i84725(x84725, x37307);
  not i84726(x84726, x37318);
  not i84727(x84727, x37319);
  not i84728(x84728, x37338);
  not i84729(x84729, x37347);
  not i84730(x84730, x37348);
  not i84731(x84731, x37355);
  not i84732(x84732, x37362);
  not i84733(x84733, x37365);
  not i84734(x84734, x37366);
  not i84735(x84735, x37377);
  not i84736(x84736, x37378);
  not i84737(x84737, x37397);
  not i84738(x84738, x37406);
  not i84739(x84739, x37407);
  not i84740(x84740, x37414);
  not i84741(x84741, x37421);
  not i84742(x84742, x37424);
  not i84743(x84743, x37425);
  not i84744(x84744, x37436);
  not i84745(x84745, x37437);
  not i84746(x84746, x37456);
  not i84747(x84747, x37465);
  not i84748(x84748, x37466);
  not i84749(x84749, x37473);
  not i84750(x84750, x37480);
  not i84751(x84751, x37483);
  not i84752(x84752, x37484);
  not i84753(x84753, x37495);
  not i84754(x84754, x37496);
  not i84755(x84755, x37515);
  not i84756(x84756, x37524);
  not i84757(x84757, x37525);
  not i84758(x84758, x37532);
  not i84759(x84759, x37539);
  not i84760(x84760, x37542);
  not i84761(x84761, x37543);
  not i84762(x84762, x37554);
  not i84763(x84763, x37555);
  not i84764(x84764, x37574);
  not i84765(x84765, x37583);
  not i84766(x84766, x37584);
  not i84767(x84767, x37591);
  not i84768(x84768, x37598);
  not i84769(x84769, x37601);
  not i84770(x84770, x37602);
  not i84771(x84771, x37613);
  not i84772(x84772, x37614);
  not i84773(x84773, x37633);
  not i84774(x84774, x37642);
  not i84775(x84775, x37643);
  not i84776(x84776, x37650);
  not i84777(x84777, x37657);
  not i84778(x84778, x37660);
  not i84779(x84779, x37661);
  not i84780(x84780, x37672);
  not i84781(x84781, x37673);
  not i84782(x84782, x37692);
  not i84783(x84783, x37701);
  not i84784(x84784, x37702);
  not i84785(x84785, x37709);
  not i84786(x84786, x37716);
  not i84787(x84787, x37719);
  not i84788(x84788, x37720);
  not i84789(x84789, x37731);
  not i84790(x84790, x37732);
  not i84791(x84791, x37751);
  not i84792(x84792, x37760);
  not i84793(x84793, x37761);
  not i84794(x84794, x37768);
  not i84795(x84795, x37775);
  not i84796(x84796, x37778);
  not i84797(x84797, x37779);
  not i84798(x84798, x37790);
  not i84799(x84799, x37791);
  not i84800(x84800, x37810);
  not i84801(x84801, x37819);
  not i84802(x84802, x37820);
  not i84803(x84803, x37827);
  not i84804(x84804, x37834);
  not i84805(x84805, x37837);
  not i84806(x84806, x37838);
  not i84807(x84807, x37849);
  not i84808(x84808, x37850);
  not i84809(x84809, x37869);
  not i84810(x84810, x37878);
  not i84811(x84811, x37879);
  not i84812(x84812, x37886);
  not i84813(x84813, x37893);
  not i84814(x84814, x37896);
  not i84815(x84815, x37897);
  not i84816(x84816, x37908);
  not i84817(x84817, x37909);
  not i84818(x84818, x37928);
  not i84819(x84819, x37937);
  not i84820(x84820, x37938);
  not i84821(x84821, x37945);
  not i84822(x84822, x37952);
  not i84823(x84823, x37955);
  not i84824(x84824, x37956);
  not i84825(x84825, x37967);
  not i84826(x84826, x37968);
  not i84827(x84827, x37987);
  not i84828(x84828, x37996);
  not i84829(x84829, x37997);
  not i84830(x84830, x38004);
  not i84831(x84831, x38011);
  not i84832(x84832, x38014);
  not i84833(x84833, x38015);
  not i84834(x84834, x38026);
  not i84835(x84835, x38027);
  not i84836(x84836, x38046);
  not i84837(x84837, x38055);
  not i84838(x84838, x38056);
  not i84839(x84839, x38063);
  not i84840(x84840, x38070);
  not i84841(x84841, x38073);
  not i84842(x84842, x38074);
  not i84843(x84843, x38085);
  not i84844(x84844, x38086);
  not i84845(x84845, x38105);
  not i84846(x84846, x38114);
  not i84847(x84847, x38115);
  not i84848(x84848, x38122);
  not i84849(x84849, x38129);
  not i84850(x84850, x38132);
  not i84851(x84851, x38133);
  not i84852(x84852, x38144);
  not i84853(x84853, x38145);
  not i84854(x84854, x38164);
  not i84855(x84855, x38173);
  not i84856(x84856, x38174);
  not i84857(x84857, x38181);
  not i84858(x84858, x38188);
  not i84859(x84859, x38191);
  not i84860(x84860, x38192);
  not i84861(x84861, x38203);
  not i84862(x84862, x38204);
  not i84863(x84863, x38223);
  not i84864(x84864, x38232);
  not i84865(x84865, x38233);
  not i84866(x84866, x38240);
  not i84867(x84867, x38247);
  not i84868(x84868, x38250);
  not i84869(x84869, x38251);
  not i84870(x84870, x38262);
  not i84871(x84871, x38263);
  not i84872(x84872, x38282);
  not i84873(x84873, x38291);
  not i84874(x84874, x38292);
  not i84875(x84875, x38299);
  not i84876(x84876, x38306);
  not i84877(x84877, x38309);
  not i84878(x84878, x38310);
  not i84879(x84879, x38321);
  not i84880(x84880, x38322);
  not i84881(x84881, x38341);
  not i84882(x84882, x38350);
  not i84883(x84883, x38351);
  not i84884(x84884, x38358);
  not i84885(x84885, x38365);
  not i84886(x84886, x38368);
  not i84887(x84887, x38369);
  not i84888(x84888, x38380);
  not i84889(x84889, x38381);
  not i84890(x84890, x38400);
  not i84891(x84891, x38409);
  not i84892(x84892, x38410);
  not i84893(x84893, x38417);
  not i84894(x84894, x38424);
  not i84895(x84895, x38427);
  not i84896(x84896, x38428);
  not i84897(x84897, x38439);
  not i84898(x84898, x38440);
  not i84899(x84899, x38459);
  not i84900(x84900, x38468);
  not i84901(x84901, x38469);
  not i84902(x84902, x38476);
  not i84903(x84903, x38483);
  not i84904(x84904, x38486);
  not i84905(x84905, x38487);
  not i84906(x84906, x38498);
  not i84907(x84907, x38499);
  not i84908(x84908, x38518);
  not i84909(x84909, x38527);
  not i84910(x84910, x38528);
  not i84911(x84911, x38535);
  not i84912(x84912, x38542);
  not i84913(x84913, x38545);
  not i84914(x84914, x38546);
  not i84915(x84915, x38557);
  not i84916(x84916, x38558);
  not i84917(x84917, x38577);
  not i84918(x84918, x38586);
  not i84919(x84919, x38587);
  not i84920(x84920, x38594);
  not i84921(x84921, x38601);
  not i84922(x84922, x38604);
  not i84923(x84923, x38605);
  not i84924(x84924, x38616);
  not i84925(x84925, x38617);
  not i84926(x84926, x38636);
  not i84927(x84927, x38645);
  not i84928(x84928, x38646);
  not i84929(x84929, x38653);
  not i84930(x84930, x38660);
  not i84931(x84931, x38663);
  not i84932(x84932, x38664);
  not i84933(x84933, x38675);
  not i84934(x84934, x38676);
  not i84935(x84935, x38695);
  not i84936(x84936, x38704);
  not i84937(x84937, x38705);
  not i84938(x84938, x38712);
  not i84939(x84939, x41043);
  not i84940(x84940, x40023);
  not i84941(x84941, x41098);
  not i84942(x84942, x41096);
  not i84943(x84943, x40076);
  not i84944(x84944, x41179);
  not i84945(x84945, x41285);
  not i84946(x84946, x40236);
  not i84947(x84947, x41421);
  not i84948(x84948, x41419);
  not i84949(x84949, x40343);
  not i84950(x84950, x41583);
  not i84951(x84951, x41770);
  not i84952(x84952, x40611);
  not i84953(x84953, x41987);
  not i84954(x84954, x41985);
  not i84955(x84955, x40772);
  not i84956(x84956, x42230);
  not i84957(x84957, x40951);
  not i84958(x84958, x39988);
  not i84959(x84959, x41045);
  not i84960(x84960, x41060);
  not i84961(x84961, x42508);
  not i84962(x84962, x42516);
  not i84963(x84963, x42529);
  not i84964(x84964, x41177);
  not i84965(x84965, x42646);
  not i84966(x84966, x42643);
  not i84967(x84967, x42671);
  not i84968(x84968, x42667);
  not i84969(x84969, x42681);
  not i84970(x84970, x42699);
  not i84971(x84971, x42695);
  not i84972(x84972, x42709);
  not i84973(x84973, x42743);
  not i84974(x84974, x41581);
  not i84975(x84975, x41590);
  not i84976(x84976, x41652);
  not i84977(x84977, x40468);
  not i84978(x84978, x41714);
  not i84979(x84979, x41772);
  not i84980(x84980, x42976);
  not i84981(x84981, x42973);
  not i84982(x84982, x41779);
  not i84983(x84983, x41841);
  not i84984(x84984, x43022);
  not i84985(x84985, x43018);
  not i84986(x84986, x41849);
  not i84987(x84987, x43043);
  not i84988(x84988, x43041);
  not i84989(x84989, x43072);
  not i84990(x84990, x43068);
  not i84991(x84991, x41920);
  not i84992(x84992, x43093);
  not i84993(x84993, x43091);
  not i84994(x84994, x41994);
  not i84995(x84995, x43149);
  not i84996(x84996, x43147);
  not i84997(x84997, x42074);
  not i84998(x84998, x42154);
  not i84999(x84999, x42228);
  not i85000(x85000, x43312);
  not i85001(x85001, x43380);
  not i85002(x85002, x41016);
  not i85003(x85003, x41025);
  not i85004(x85004, x41033);
  not i85005(x85005, x41041);
  not i85006(x85006, x41052);
  not i85007(x85007, x42497);
  not i85008(x85008, x41068);
  not i85009(x85009, x42501);
  not i85010(x85010, x42506);
  not i85011(x85011, x42513);
  not i85012(x85012, x41085);
  not i85013(x85013, x42509);
  not i85014(x85014, x42514);
  not i85015(x85015, x42525);
  not i85016(x85016, x41105);
  not i85017(x85017, x42527);
  not i85018(x85018, x42539);
  not i85019(x85019, x41131);
  not i85020(x85020, x42559);
  not i85021(x85021, x41157);
  not i85022(x85022, x42579);
  not i85023(x85023, x41186);
  not i85024(x85024, x42599);
  not i85025(x85025, x41221);
  not i85026(x85026, x40147);
  not i85027(x85027, x42620);
  not i85028(x85028, x41256);
  not i85029(x85029, x41287);
  not i85030(x85030, x42641);
  not i85031(x85031, x41294);
  not i85032(x85032, x41329);
  not i85033(x85033, x43551);
  not i85034(x85034, x42665);
  not i85035(x85035, x43553);
  not i85036(x85036, x41337);
  not i85037(x85037, x42683);
  not i85038(x85038, x43564);
  not i85039(x85039, x43561);
  not i85040(x85040, x43566);
  not i85041(x85041, x42693);
  not i85042(x85042, x43570);
  not i85043(x85043, x41381);
  not i85044(x85044, x42711);
  not i85045(x85045, x43581);
  not i85046(x85046, x43578);
  not i85047(x85047, x43583);
  not i85048(x85048, x42721);
  not i85049(x85049, x43587);
  not i85050(x85050, x41428);
  not i85051(x85051, x42745);
  not i85052(x85052, x43599);
  not i85053(x85053, x43595);
  not i85054(x85054, x43601);
  not i85055(x85055, x42755);
  not i85056(x85056, x43605);
  not i85057(x85057, x41481);
  not i85058(x85058, x42784);
  not i85059(x85059, x43617);
  not i85060(x85060, x43613);
  not i85061(x85061, x43619);
  not i85062(x85062, x42795);
  not i85063(x85063, x43624);
  not i85064(x85064, x41534);
  not i85065(x85065, x42824);
  not i85066(x85066, x43636);
  not i85067(x85067, x43632);
  not i85068(x85068, x43638);
  not i85069(x85069, x42835);
  not i85070(x85070, x43643);
  not i85071(x85071, x42864);
  not i85072(x85072, x43660);
  not i85073(x85073, x43656);
  not i85074(x85074, x43662);
  not i85075(x85075, x42875);
  not i85076(x85076, x43667);
  not i85077(x85077, x43682);
  not i85078(x85078, x43680);
  not i85079(x85079, x43687);
  not i85080(x85080, x43683);
  not i85081(x85081, x43689);
  not i85082(x85082, x42917);
  not i85083(x85083, x43694);
  not i85084(x85084, x43709);
  not i85085(x85085, x43707);
  not i85086(x85086, x43714);
  not i85087(x85087, x43710);
  not i85088(x85088, x43716);
  not i85089(x85089, x42959);
  not i85090(x85090, x43721);
  not i85091(x85091, x43736);
  not i85092(x85092, x43734);
  not i85093(x85093, x43749);
  not i85094(x85094, x43004);
  not i85095(x85095, x43754);
  not i85096(x85096, x43769);
  not i85097(x85097, x43767);
  not i85098(x85098, x43782);
  not i85099(x85099, x43807);
  not i85100(x85100, x43805);
  not i85101(x85101, x43820);
  not i85102(x85102, x43845);
  not i85103(x85103, x43843);
  not i85104(x85104, x43859);
  not i85105(x85105, x43884);
  not i85106(x85106, x43882);
  not i85107(x85107, x43898);
  not i85108(x85108, x43924);
  not i85109(x85109, x43922);
  not i85110(x85110, x43938);
  not i85111(x85111, x43964);
  not i85112(x85112, x43962);
  not i85113(x85113, x42500);
  not i85114(x85114, x43481);
  not i85115(x85115, x42505);
  not i85116(x85116, x44079);
  not i85117(x85117, x43485);
  not i85118(x85118, x43489);
  not i85119(x85119, x43493);
  not i85120(x85120, x43498);
  not i85121(x85121, x43504);
  not i85122(x85122, x43510);
  not i85123(x85123, x43514);
  not i85124(x85124, x43520);
  not i85125(x85125, x43524);
  not i85126(x85126, x43530);
  not i85127(x85127, x43534);
  not i85128(x85128, x43540);
  not i85129(x85129, x43544);
  not i85130(x85130, x43548);
  not i85131(x85131, x44195);
  not i85132(x85132, x43557);
  not i85133(x85133, x44199);
  not i85134(x85134, x43574);
  not i85135(x85135, x44221);
  not i85136(x85136, x43591);
  not i85137(x85137, x44243);
  not i85138(x85138, x43609);
  not i85139(x85139, x44265);
  not i85140(x85140, x43628);
  not i85141(x85141, x44287);
  not i85142(x85142, x44310);
  not i85143(x85143, x43473);
  not i85144(x85144, x44068);
  not i85145(x85145, x43477);
  not i85146(x85146, x44072);
  not i85147(x85147, x44078);
  not i85148(x85148, x44076);
  not i85149(x85149, x44624);
  not i85150(x85150, x44085);
  not i85151(x85151, x44628);
  not i85152(x85152, x44083);
  not i85153(x85153, x44631);
  not i85154(x85154, x44097);
  not i85155(x85155, x44636);
  not i85156(x85156, x44095);
  not i85157(x85157, x44639);
  not i85158(x85158, x44109);
  not i85159(x85159, x44644);
  not i85160(x85160, x44107);
  not i85161(x85161, x44647);
  not i85162(x85162, x44121);
  not i85163(x85163, x44652);
  not i85164(x85164, x44119);
  not i85165(x85165, x44655);
  not i85166(x85166, x44133);
  not i85167(x85167, x44660);
  not i85168(x85168, x44131);
  not i85169(x85169, x44663);
  not i85170(x85170, x44143);
  not i85171(x85171, x44677);
  not i85172(x85172, x44156);
  not i85173(x85173, x44691);
  not i85174(x85174, x44169);
  not i85175(x85175, x44705);
  not i85176(x85176, x44182);
  not i85177(x85177, x44719);
  not i85178(x85178, x44067);
  not i85179(x85179, x44617);
  not i85180(x85180, x44615);
  not i85181(x85181, x44620);
  not i85182(x85182, x44618);
  not i85183(x85183, x44623);
  not i85184(x85184, x44621);
  not i85185(x85185, x44630);
  not i85186(x85186, x44638);
  not i85187(x85187, x44646);
  not i85188(x85188, x44654);
  not i85189(x85189, x44662);
  not i85190(x85190, x44062);
  not i85191(x85191, x45397);
  not i85192(x85192, x44065);
  not i85193(x85193, x45039);
  not i85194(x85194, x45400);
  not i85195(x85195, x45042);
  not i85196(x85196, x45403);
  not i85197(x85197, x45046);
  not i85198(x85198, x45407);
  not i85199(x85199, x45412);
  not i85200(x85200, x45417);
  not i85201(x85201, x45422);
  not i85202(x85202, x45427);
  not i85203(x85203, x45041);
  not i85204(x85204, x45628);
  not i85205(x85205, x45402);
  not i85206(x85206, x45632);
  not i85207(x85207, x41018);
  not i85208(x85208, x44064);
  not i85209(x85209, x45399);
  not i85210(x85210, x45626);
  not i85211(x85211, x45881);
  not i85212(x85212, x46643);
  not i85213(x85213, x46700);
  not i85214(x85214, x46701);
  not i85215(x85215, x46702);
  not i85216(x85216, x46751);
  not i85217(x85217, x46752);
  not i85218(x85218, x46753);
  not i85219(x85219, x46754);
  not i85220(x85220, x46755);
  not i85221(x85221, x46756);
  not i85222(x85222, x46757);
  not i85223(x85223, x46758);
  not i85224(x85224, x46789);
  not i85225(x85225, x46790);
  not i85226(x85226, x46791);
  not i85227(x85227, x46792);
  not i85228(x85228, x46793);
  not i85229(x85229, x46794);
  not i85230(x85230, x46795);
  not i85231(x85231, x46796);
  not i85232(x85232, x46797);
  not i85233(x85233, x46798);
  not i85234(x85234, x46799);
  not i85235(x85235, x46800);
  not i85236(x85236, x46801);
  not i85237(x85237, x46802);
  not i85238(x85238, x46803);
  not i85239(x85239, x47056);
  not i85240(x85240, x47119);
  not i85241(x85241, x47120);
  not i85242(x85242, x47211);
  not i85243(x85243, x47212);
  not i85244(x85244, x47213);
  not i85245(x85245, x47214);
  not i85246(x85246, x47299);
  not i85247(x85247, x47300);
  not i85248(x85248, x47301);
  not i85249(x85249, x47302);
  not i85250(x85250, x47303);
  not i85251(x85251, x47304);
  not i85252(x85252, x47305);
  not i85253(x85253, x47306);
  not i85254(x85254, x47379);
  not i85255(x85255, x47380);
  not i85256(x85256, x47381);
  not i85257(x85257, x47382);
  not i85258(x85258, x47383);
  not i85259(x85259, x47384);
  not i85260(x85260, x47385);
  not i85261(x85261, x47386);
  not i85262(x85262, x47387);
  not i85263(x85263, x47388);
  not i85264(x85264, x47389);
  not i85265(x85265, x47390);
  not i85266(x85266, x47391);
  not i85267(x85267, x47392);
  not i85268(x85268, x47393);
  not i85269(x85269, x47394);
  not i85270(x85270, x47117);
  not i85271(x85271, x47564);
  not i85272(x85272, x47565);
  not i85273(x85273, x47650);
  not i85274(x85274, x47651);
  not i85275(x85275, x47652);
  not i85276(x85276, x47653);
  not i85277(x85277, x47726);
  not i85278(x85278, x47727);
  not i85279(x85279, x47728);
  not i85280(x85280, x47729);
  not i85281(x85281, x47730);
  not i85282(x85282, x47731);
  not i85283(x85283, x47732);
  not i85284(x85284, x47733);
  not i85285(x85285, x47782);
  not i85286(x85286, x47783);
  not i85287(x85287, x47784);
  not i85288(x85288, x47785);
  not i85289(x85289, x47786);
  not i85290(x85290, x47787);
  not i85291(x85291, x47788);
  not i85292(x85292, x47789);
  not i85293(x85293, x47790);
  not i85294(x85294, x47791);
  not i85295(x85295, x47792);
  not i85296(x85296, x47793);
  not i85297(x85297, x47794);
  not i85298(x85298, x47795);
  not i85299(x85299, x47796);
  not i85300(x85300, x47797);
  not i85301(x85301, x47798);
  not i85302(x85302, x47801);
  not i85303(x85303, x47802);
  not i85304(x85304, x47813);
  not i85305(x85305, x47814);
  not i85306(x85306, x47833);
  not i85307(x85307, x47842);
  not i85308(x85308, x47843);
  not i85309(x85309, x47850);
  not i85310(x85310, x47857);
  not i85311(x85311, x47860);
  not i85312(x85312, x47861);
  not i85313(x85313, x47872);
  not i85314(x85314, x47873);
  not i85315(x85315, x47892);
  not i85316(x85316, x47901);
  not i85317(x85317, x47902);
  not i85318(x85318, x47909);
  not i85319(x85319, x47916);
  not i85320(x85320, x47919);
  not i85321(x85321, x47920);
  not i85322(x85322, x47931);
  not i85323(x85323, x47932);
  not i85324(x85324, x47951);
  not i85325(x85325, x47960);
  not i85326(x85326, x47961);
  not i85327(x85327, x47968);
  not i85328(x85328, x47975);
  not i85329(x85329, x47978);
  not i85330(x85330, x47979);
  not i85331(x85331, x47990);
  not i85332(x85332, x47991);
  not i85333(x85333, x48010);
  not i85334(x85334, x48019);
  not i85335(x85335, x48020);
  not i85336(x85336, x48027);
  not i85337(x85337, x48034);
  not i85338(x85338, x48037);
  not i85339(x85339, x48038);
  not i85340(x85340, x48049);
  not i85341(x85341, x48050);
  not i85342(x85342, x48069);
  not i85343(x85343, x48078);
  not i85344(x85344, x48079);
  not i85345(x85345, x48086);
  not i85346(x85346, x48093);
  not i85347(x85347, x48096);
  not i85348(x85348, x48097);
  not i85349(x85349, x48108);
  not i85350(x85350, x48109);
  not i85351(x85351, x48128);
  not i85352(x85352, x48137);
  not i85353(x85353, x48138);
  not i85354(x85354, x48145);
  not i85355(x85355, x48152);
  not i85356(x85356, x48155);
  not i85357(x85357, x48156);
  not i85358(x85358, x48167);
  not i85359(x85359, x48168);
  not i85360(x85360, x48187);
  not i85361(x85361, x48196);
  not i85362(x85362, x48197);
  not i85363(x85363, x48204);
  not i85364(x85364, x48211);
  not i85365(x85365, x48214);
  not i85366(x85366, x48215);
  not i85367(x85367, x48226);
  not i85368(x85368, x48227);
  not i85369(x85369, x48246);
  not i85370(x85370, x48255);
  not i85371(x85371, x48256);
  not i85372(x85372, x48263);
  not i85373(x85373, x48270);
  not i85374(x85374, x48273);
  not i85375(x85375, x48274);
  not i85376(x85376, x48285);
  not i85377(x85377, x48286);
  not i85378(x85378, x48305);
  not i85379(x85379, x48314);
  not i85380(x85380, x48315);
  not i85381(x85381, x48322);
  not i85382(x85382, x48329);
  not i85383(x85383, x48332);
  not i85384(x85384, x48333);
  not i85385(x85385, x48344);
  not i85386(x85386, x48345);
  not i85387(x85387, x48364);
  not i85388(x85388, x48373);
  not i85389(x85389, x48374);
  not i85390(x85390, x48381);
  not i85391(x85391, x48388);
  not i85392(x85392, x48391);
  not i85393(x85393, x48392);
  not i85394(x85394, x48403);
  not i85395(x85395, x48404);
  not i85396(x85396, x48423);
  not i85397(x85397, x48432);
  not i85398(x85398, x48433);
  not i85399(x85399, x48440);
  not i85400(x85400, x48447);
  not i85401(x85401, x48450);
  not i85402(x85402, x48451);
  not i85403(x85403, x48462);
  not i85404(x85404, x48463);
  not i85405(x85405, x48482);
  not i85406(x85406, x48491);
  not i85407(x85407, x48492);
  not i85408(x85408, x48499);
  not i85409(x85409, x48506);
  not i85410(x85410, x48509);
  not i85411(x85411, x48510);
  not i85412(x85412, x48521);
  not i85413(x85413, x48522);
  not i85414(x85414, x48541);
  not i85415(x85415, x48550);
  not i85416(x85416, x48551);
  not i85417(x85417, x48558);
  not i85418(x85418, x48565);
  not i85419(x85419, x48568);
  not i85420(x85420, x48569);
  not i85421(x85421, x48580);
  not i85422(x85422, x48581);
  not i85423(x85423, x48600);
  not i85424(x85424, x48609);
  not i85425(x85425, x48610);
  not i85426(x85426, x48617);
  not i85427(x85427, x48624);
  not i85428(x85428, x48627);
  not i85429(x85429, x48628);
  not i85430(x85430, x48639);
  not i85431(x85431, x48640);
  not i85432(x85432, x48659);
  not i85433(x85433, x48668);
  not i85434(x85434, x48669);
  not i85435(x85435, x48676);
  not i85436(x85436, x48683);
  not i85437(x85437, x48686);
  not i85438(x85438, x48687);
  not i85439(x85439, x48698);
  not i85440(x85440, x48699);
  not i85441(x85441, x48718);
  not i85442(x85442, x48727);
  not i85443(x85443, x48728);
  not i85444(x85444, x48735);
  not i85445(x85445, x48742);
  not i85446(x85446, x48745);
  not i85447(x85447, x48746);
  not i85448(x85448, x48757);
  not i85449(x85449, x48758);
  not i85450(x85450, x48777);
  not i85451(x85451, x48786);
  not i85452(x85452, x48787);
  not i85453(x85453, x48794);
  not i85454(x85454, x48801);
  not i85455(x85455, x48804);
  not i85456(x85456, x48805);
  not i85457(x85457, x48816);
  not i85458(x85458, x48817);
  not i85459(x85459, x48836);
  not i85460(x85460, x48845);
  not i85461(x85461, x48846);
  not i85462(x85462, x48853);
  not i85463(x85463, x48860);
  not i85464(x85464, x48863);
  not i85465(x85465, x48864);
  not i85466(x85466, x48875);
  not i85467(x85467, x48876);
  not i85468(x85468, x48895);
  not i85469(x85469, x48904);
  not i85470(x85470, x48905);
  not i85471(x85471, x48912);
  not i85472(x85472, x48919);
  not i85473(x85473, x48922);
  not i85474(x85474, x48923);
  not i85475(x85475, x48934);
  not i85476(x85476, x48935);
  not i85477(x85477, x48954);
  not i85478(x85478, x48963);
  not i85479(x85479, x48964);
  not i85480(x85480, x48971);
  not i85481(x85481, x48978);
  not i85482(x85482, x48981);
  not i85483(x85483, x48982);
  not i85484(x85484, x48993);
  not i85485(x85485, x48994);
  not i85486(x85486, x49013);
  not i85487(x85487, x49022);
  not i85488(x85488, x49023);
  not i85489(x85489, x49030);
  not i85490(x85490, x49037);
  not i85491(x85491, x49040);
  not i85492(x85492, x49041);
  not i85493(x85493, x49052);
  not i85494(x85494, x49053);
  not i85495(x85495, x49072);
  not i85496(x85496, x49081);
  not i85497(x85497, x49082);
  not i85498(x85498, x49089);
  not i85499(x85499, x49096);
  not i85500(x85500, x49099);
  not i85501(x85501, x49100);
  not i85502(x85502, x49111);
  not i85503(x85503, x49112);
  not i85504(x85504, x49131);
  not i85505(x85505, x49140);
  not i85506(x85506, x49141);
  not i85507(x85507, x49148);
  not i85508(x85508, x49155);
  not i85509(x85509, x49158);
  not i85510(x85510, x49159);
  not i85511(x85511, x49170);
  not i85512(x85512, x49171);
  not i85513(x85513, x49190);
  not i85514(x85514, x49199);
  not i85515(x85515, x49200);
  not i85516(x85516, x49207);
  not i85517(x85517, x49214);
  not i85518(x85518, x49217);
  not i85519(x85519, x49218);
  not i85520(x85520, x49229);
  not i85521(x85521, x49230);
  not i85522(x85522, x49249);
  not i85523(x85523, x49258);
  not i85524(x85524, x49259);
  not i85525(x85525, x49266);
  not i85526(x85526, x49273);
  not i85527(x85527, x49276);
  not i85528(x85528, x49277);
  not i85529(x85529, x49288);
  not i85530(x85530, x49289);
  not i85531(x85531, x49308);
  not i85532(x85532, x49317);
  not i85533(x85533, x49318);
  not i85534(x85534, x49325);
  not i85535(x85535, x49332);
  not i85536(x85536, x49335);
  not i85537(x85537, x49336);
  not i85538(x85538, x49347);
  not i85539(x85539, x49348);
  not i85540(x85540, x49367);
  not i85541(x85541, x49376);
  not i85542(x85542, x49377);
  not i85543(x85543, x49384);
  not i85544(x85544, x49391);
  not i85545(x85545, x49394);
  not i85546(x85546, x49395);
  not i85547(x85547, x49406);
  not i85548(x85548, x49407);
  not i85549(x85549, x49426);
  not i85550(x85550, x49435);
  not i85551(x85551, x49436);
  not i85552(x85552, x49443);
  not i85553(x85553, x49450);
  not i85554(x85554, x49453);
  not i85555(x85555, x49454);
  not i85556(x85556, x49465);
  not i85557(x85557, x49466);
  not i85558(x85558, x49485);
  not i85559(x85559, x49494);
  not i85560(x85560, x49495);
  not i85561(x85561, x49502);
  not i85562(x85562, x49509);
  not i85563(x85563, x49512);
  not i85564(x85564, x49513);
  not i85565(x85565, x49524);
  not i85566(x85566, x49525);
  not i85567(x85567, x49544);
  not i85568(x85568, x49553);
  not i85569(x85569, x49554);
  not i85570(x85570, x49561);
  not i85571(x85571, x49568);
  not i85572(x85572, x49571);
  not i85573(x85573, x49572);
  not i85574(x85574, x49583);
  not i85575(x85575, x49584);
  not i85576(x85576, x49603);
  not i85577(x85577, x49612);
  not i85578(x85578, x49613);
  not i85579(x85579, x49620);
  not i85580(x85580, x49627);
  not i85581(x85581, x49630);
  not i85582(x85582, x49631);
  not i85583(x85583, x49642);
  not i85584(x85584, x49643);
  not i85585(x85585, x49662);
  not i85586(x85586, x49671);
  not i85587(x85587, x49672);
  not i85588(x85588, x49679);
  not i85589(x85589, x52010);
  not i85590(x85590, x50990);
  not i85591(x85591, x52065);
  not i85592(x85592, x52063);
  not i85593(x85593, x51043);
  not i85594(x85594, x52146);
  not i85595(x85595, x52252);
  not i85596(x85596, x51203);
  not i85597(x85597, x52388);
  not i85598(x85598, x52386);
  not i85599(x85599, x51310);
  not i85600(x85600, x52550);
  not i85601(x85601, x52737);
  not i85602(x85602, x51578);
  not i85603(x85603, x52954);
  not i85604(x85604, x52952);
  not i85605(x85605, x51739);
  not i85606(x85606, x53197);
  not i85607(x85607, x51918);
  not i85608(x85608, x50955);
  not i85609(x85609, x52012);
  not i85610(x85610, x52027);
  not i85611(x85611, x53475);
  not i85612(x85612, x53483);
  not i85613(x85613, x53496);
  not i85614(x85614, x52144);
  not i85615(x85615, x53613);
  not i85616(x85616, x53610);
  not i85617(x85617, x53638);
  not i85618(x85618, x53634);
  not i85619(x85619, x53648);
  not i85620(x85620, x53666);
  not i85621(x85621, x53662);
  not i85622(x85622, x53676);
  not i85623(x85623, x53710);
  not i85624(x85624, x52548);
  not i85625(x85625, x52557);
  not i85626(x85626, x52619);
  not i85627(x85627, x51435);
  not i85628(x85628, x52681);
  not i85629(x85629, x52739);
  not i85630(x85630, x53943);
  not i85631(x85631, x53940);
  not i85632(x85632, x52746);
  not i85633(x85633, x52808);
  not i85634(x85634, x53989);
  not i85635(x85635, x53985);
  not i85636(x85636, x52816);
  not i85637(x85637, x54010);
  not i85638(x85638, x54008);
  not i85639(x85639, x54039);
  not i85640(x85640, x54035);
  not i85641(x85641, x52887);
  not i85642(x85642, x54060);
  not i85643(x85643, x54058);
  not i85644(x85644, x52961);
  not i85645(x85645, x54116);
  not i85646(x85646, x54114);
  not i85647(x85647, x53041);
  not i85648(x85648, x53121);
  not i85649(x85649, x53195);
  not i85650(x85650, x54279);
  not i85651(x85651, x54347);
  not i85652(x85652, x51983);
  not i85653(x85653, x51992);
  not i85654(x85654, x52000);
  not i85655(x85655, x52008);
  not i85656(x85656, x52019);
  not i85657(x85657, x53464);
  not i85658(x85658, x52035);
  not i85659(x85659, x53468);
  not i85660(x85660, x53473);
  not i85661(x85661, x53480);
  not i85662(x85662, x52052);
  not i85663(x85663, x53476);
  not i85664(x85664, x53481);
  not i85665(x85665, x53492);
  not i85666(x85666, x52072);
  not i85667(x85667, x53494);
  not i85668(x85668, x53506);
  not i85669(x85669, x52098);
  not i85670(x85670, x53526);
  not i85671(x85671, x52124);
  not i85672(x85672, x53546);
  not i85673(x85673, x52153);
  not i85674(x85674, x53566);
  not i85675(x85675, x52188);
  not i85676(x85676, x51114);
  not i85677(x85677, x53587);
  not i85678(x85678, x52223);
  not i85679(x85679, x52254);
  not i85680(x85680, x53608);
  not i85681(x85681, x52261);
  not i85682(x85682, x52296);
  not i85683(x85683, x54518);
  not i85684(x85684, x53632);
  not i85685(x85685, x54520);
  not i85686(x85686, x52304);
  not i85687(x85687, x53650);
  not i85688(x85688, x54531);
  not i85689(x85689, x54528);
  not i85690(x85690, x54533);
  not i85691(x85691, x53660);
  not i85692(x85692, x54537);
  not i85693(x85693, x52348);
  not i85694(x85694, x53678);
  not i85695(x85695, x54548);
  not i85696(x85696, x54545);
  not i85697(x85697, x54550);
  not i85698(x85698, x53688);
  not i85699(x85699, x54554);
  not i85700(x85700, x52395);
  not i85701(x85701, x53712);
  not i85702(x85702, x54566);
  not i85703(x85703, x54562);
  not i85704(x85704, x54568);
  not i85705(x85705, x53722);
  not i85706(x85706, x54572);
  not i85707(x85707, x52448);
  not i85708(x85708, x53751);
  not i85709(x85709, x54584);
  not i85710(x85710, x54580);
  not i85711(x85711, x54586);
  not i85712(x85712, x53762);
  not i85713(x85713, x54591);
  not i85714(x85714, x52501);
  not i85715(x85715, x53791);
  not i85716(x85716, x54603);
  not i85717(x85717, x54599);
  not i85718(x85718, x54605);
  not i85719(x85719, x53802);
  not i85720(x85720, x54610);
  not i85721(x85721, x53831);
  not i85722(x85722, x54627);
  not i85723(x85723, x54623);
  not i85724(x85724, x54629);
  not i85725(x85725, x53842);
  not i85726(x85726, x54634);
  not i85727(x85727, x54649);
  not i85728(x85728, x54647);
  not i85729(x85729, x54654);
  not i85730(x85730, x54650);
  not i85731(x85731, x54656);
  not i85732(x85732, x53884);
  not i85733(x85733, x54661);
  not i85734(x85734, x54676);
  not i85735(x85735, x54674);
  not i85736(x85736, x54681);
  not i85737(x85737, x54677);
  not i85738(x85738, x54683);
  not i85739(x85739, x53926);
  not i85740(x85740, x54688);
  not i85741(x85741, x54703);
  not i85742(x85742, x54701);
  not i85743(x85743, x54716);
  not i85744(x85744, x53971);
  not i85745(x85745, x54721);
  not i85746(x85746, x54736);
  not i85747(x85747, x54734);
  not i85748(x85748, x54749);
  not i85749(x85749, x54774);
  not i85750(x85750, x54772);
  not i85751(x85751, x54787);
  not i85752(x85752, x54812);
  not i85753(x85753, x54810);
  not i85754(x85754, x54826);
  not i85755(x85755, x54851);
  not i85756(x85756, x54849);
  not i85757(x85757, x54865);
  not i85758(x85758, x54891);
  not i85759(x85759, x54889);
  not i85760(x85760, x54905);
  not i85761(x85761, x54931);
  not i85762(x85762, x54929);
  not i85763(x85763, x53467);
  not i85764(x85764, x54448);
  not i85765(x85765, x53472);
  not i85766(x85766, x55046);
  not i85767(x85767, x54452);
  not i85768(x85768, x54456);
  not i85769(x85769, x54460);
  not i85770(x85770, x54465);
  not i85771(x85771, x54471);
  not i85772(x85772, x54477);
  not i85773(x85773, x54481);
  not i85774(x85774, x54487);
  not i85775(x85775, x54491);
  not i85776(x85776, x54497);
  not i85777(x85777, x54501);
  not i85778(x85778, x54507);
  not i85779(x85779, x54511);
  not i85780(x85780, x54515);
  not i85781(x85781, x55162);
  not i85782(x85782, x54524);
  not i85783(x85783, x55166);
  not i85784(x85784, x54541);
  not i85785(x85785, x55188);
  not i85786(x85786, x54558);
  not i85787(x85787, x55210);
  not i85788(x85788, x54576);
  not i85789(x85789, x55232);
  not i85790(x85790, x54595);
  not i85791(x85791, x55254);
  not i85792(x85792, x55277);
  not i85793(x85793, x54440);
  not i85794(x85794, x55035);
  not i85795(x85795, x54444);
  not i85796(x85796, x55039);
  not i85797(x85797, x55045);
  not i85798(x85798, x55043);
  not i85799(x85799, x55591);
  not i85800(x85800, x55052);
  not i85801(x85801, x55595);
  not i85802(x85802, x55050);
  not i85803(x85803, x55598);
  not i85804(x85804, x55064);
  not i85805(x85805, x55603);
  not i85806(x85806, x55062);
  not i85807(x85807, x55606);
  not i85808(x85808, x55076);
  not i85809(x85809, x55611);
  not i85810(x85810, x55074);
  not i85811(x85811, x55614);
  not i85812(x85812, x55088);
  not i85813(x85813, x55619);
  not i85814(x85814, x55086);
  not i85815(x85815, x55622);
  not i85816(x85816, x55100);
  not i85817(x85817, x55627);
  not i85818(x85818, x55098);
  not i85819(x85819, x55630);
  not i85820(x85820, x55110);
  not i85821(x85821, x55644);
  not i85822(x85822, x55123);
  not i85823(x85823, x55658);
  not i85824(x85824, x55136);
  not i85825(x85825, x55672);
  not i85826(x85826, x55149);
  not i85827(x85827, x55686);
  not i85828(x85828, x55034);
  not i85829(x85829, x55584);
  not i85830(x85830, x55582);
  not i85831(x85831, x55587);
  not i85832(x85832, x55585);
  not i85833(x85833, x55590);
  not i85834(x85834, x55588);
  not i85835(x85835, x55597);
  not i85836(x85836, x55605);
  not i85837(x85837, x55613);
  not i85838(x85838, x55621);
  not i85839(x85839, x55629);
  not i85840(x85840, x55029);
  not i85841(x85841, x56364);
  not i85842(x85842, x55032);
  not i85843(x85843, x56006);
  not i85844(x85844, x56367);
  not i85845(x85845, x56009);
  not i85846(x85846, x56370);
  not i85847(x85847, x56013);
  not i85848(x85848, x56374);
  not i85849(x85849, x56379);
  not i85850(x85850, x56384);
  not i85851(x85851, x56389);
  not i85852(x85852, x56394);
  not i85853(x85853, x56008);
  not i85854(x85854, x56595);
  not i85855(x85855, x56369);
  not i85856(x85856, x56599);
  not i85857(x85857, x51985);
  not i85858(x85858, x55031);
  not i85859(x85859, x56366);
  not i85860(x85860, x56593);
  not i85861(x85861, x56848);
  not i85862(x85862, x57610);
  not i85863(x85863, x57667);
  not i85864(x85864, x57668);
  not i85865(x85865, x57669);
  not i85866(x85866, x57718);
  not i85867(x85867, x57719);
  not i85868(x85868, x57720);
  not i85869(x85869, x57721);
  not i85870(x85870, x57722);
  not i85871(x85871, x57723);
  not i85872(x85872, x57724);
  not i85873(x85873, x57725);
  not i85874(x85874, x57756);
  not i85875(x85875, x57757);
  not i85876(x85876, x57758);
  not i85877(x85877, x57759);
  not i85878(x85878, x57760);
  not i85879(x85879, x57761);
  not i85880(x85880, x57762);
  not i85881(x85881, x57763);
  not i85882(x85882, x57764);
  not i85883(x85883, x57765);
  not i85884(x85884, x57766);
  not i85885(x85885, x57767);
  not i85886(x85886, x57768);
  not i85887(x85887, x57769);
  not i85888(x85888, x57770);
  not i85889(x85889, x58023);
  not i85890(x85890, x58086);
  not i85891(x85891, x58087);
  not i85892(x85892, x58178);
  not i85893(x85893, x58179);
  not i85894(x85894, x58180);
  not i85895(x85895, x58181);
  not i85896(x85896, x58266);
  not i85897(x85897, x58267);
  not i85898(x85898, x58268);
  not i85899(x85899, x58269);
  not i85900(x85900, x58270);
  not i85901(x85901, x58271);
  not i85902(x85902, x58272);
  not i85903(x85903, x58273);
  not i85904(x85904, x58346);
  not i85905(x85905, x58347);
  not i85906(x85906, x58348);
  not i85907(x85907, x58349);
  not i85908(x85908, x58350);
  not i85909(x85909, x58351);
  not i85910(x85910, x58352);
  not i85911(x85911, x58353);
  not i85912(x85912, x58354);
  not i85913(x85913, x58355);
  not i85914(x85914, x58356);
  not i85915(x85915, x58357);
  not i85916(x85916, x58358);
  not i85917(x85917, x58359);
  not i85918(x85918, x58360);
  not i85919(x85919, x58361);
  not i85920(x85920, x58084);
  not i85921(x85921, x58531);
  not i85922(x85922, x58532);
  not i85923(x85923, x58617);
  not i85924(x85924, x58618);
  not i85925(x85925, x58619);
  not i85926(x85926, x58620);
  not i85927(x85927, x58693);
  not i85928(x85928, x58694);
  not i85929(x85929, x58695);
  not i85930(x85930, x58696);
  not i85931(x85931, x58697);
  not i85932(x85932, x58698);
  not i85933(x85933, x58699);
  not i85934(x85934, x58700);
  not i85935(x85935, x58749);
  not i85936(x85936, x58750);
  not i85937(x85937, x58751);
  not i85938(x85938, x58752);
  not i85939(x85939, x58753);
  not i85940(x85940, x58754);
  not i85941(x85941, x58755);
  not i85942(x85942, x58756);
  not i85943(x85943, x58757);
  not i85944(x85944, x58758);
  not i85945(x85945, x58759);
  not i85946(x85946, x58760);
  not i85947(x85947, x58761);
  not i85948(x85948, x58762);
  not i85949(x85949, x58763);
  not i85950(x85950, x58764);
  not i85951(x85951, x58765);
  not i85952(x85952, x58768);
  not i85953(x85953, x58769);
  not i85954(x85954, x58780);
  not i85955(x85955, x58781);
  not i85956(x85956, x58800);
  not i85957(x85957, x58809);
  not i85958(x85958, x58810);
  not i85959(x85959, x58817);
  not i85960(x85960, x58824);
  not i85961(x85961, x58827);
  not i85962(x85962, x58828);
  not i85963(x85963, x58839);
  not i85964(x85964, x58840);
  not i85965(x85965, x58859);
  not i85966(x85966, x58868);
  not i85967(x85967, x58869);
  not i85968(x85968, x58876);
  not i85969(x85969, x58883);
  not i85970(x85970, x58886);
  not i85971(x85971, x58887);
  not i85972(x85972, x58898);
  not i85973(x85973, x58899);
  not i85974(x85974, x58918);
  not i85975(x85975, x58927);
  not i85976(x85976, x58928);
  not i85977(x85977, x58935);
  not i85978(x85978, x58942);
  not i85979(x85979, x58945);
  not i85980(x85980, x58946);
  not i85981(x85981, x58957);
  not i85982(x85982, x58958);
  not i85983(x85983, x58977);
  not i85984(x85984, x58986);
  not i85985(x85985, x58987);
  not i85986(x85986, x58994);
  not i85987(x85987, x59001);
  not i85988(x85988, x59004);
  not i85989(x85989, x59005);
  not i85990(x85990, x59016);
  not i85991(x85991, x59017);
  not i85992(x85992, x59036);
  not i85993(x85993, x59045);
  not i85994(x85994, x59046);
  not i85995(x85995, x59053);
  not i85996(x85996, x59060);
  not i85997(x85997, x59063);
  not i85998(x85998, x59064);
  not i85999(x85999, x59075);
  not i86000(x86000, x59076);
  not i86001(x86001, x59095);
  not i86002(x86002, x59104);
  not i86003(x86003, x59105);
  not i86004(x86004, x59112);
  not i86005(x86005, x59119);
  not i86006(x86006, x59122);
  not i86007(x86007, x59123);
  not i86008(x86008, x59134);
  not i86009(x86009, x59135);
  not i86010(x86010, x59154);
  not i86011(x86011, x59163);
  not i86012(x86012, x59164);
  not i86013(x86013, x59171);
  not i86014(x86014, x59178);
  not i86015(x86015, x59181);
  not i86016(x86016, x59182);
  not i86017(x86017, x59193);
  not i86018(x86018, x59194);
  not i86019(x86019, x59213);
  not i86020(x86020, x59222);
  not i86021(x86021, x59223);
  not i86022(x86022, x59230);
  not i86023(x86023, x59237);
  not i86024(x86024, x59240);
  not i86025(x86025, x59241);
  not i86026(x86026, x59252);
  not i86027(x86027, x59253);
  not i86028(x86028, x59272);
  not i86029(x86029, x59281);
  not i86030(x86030, x59282);
  not i86031(x86031, x59289);
  not i86032(x86032, x59296);
  not i86033(x86033, x59299);
  not i86034(x86034, x59300);
  not i86035(x86035, x59311);
  not i86036(x86036, x59312);
  not i86037(x86037, x59331);
  not i86038(x86038, x59340);
  not i86039(x86039, x59341);
  not i86040(x86040, x59348);
  not i86041(x86041, x59355);
  not i86042(x86042, x59358);
  not i86043(x86043, x59359);
  not i86044(x86044, x59370);
  not i86045(x86045, x59371);
  not i86046(x86046, x59390);
  not i86047(x86047, x59399);
  not i86048(x86048, x59400);
  not i86049(x86049, x59407);
  not i86050(x86050, x59414);
  not i86051(x86051, x59417);
  not i86052(x86052, x59418);
  not i86053(x86053, x59429);
  not i86054(x86054, x59430);
  not i86055(x86055, x59449);
  not i86056(x86056, x59458);
  not i86057(x86057, x59459);
  not i86058(x86058, x59466);
  not i86059(x86059, x59473);
  not i86060(x86060, x59476);
  not i86061(x86061, x59477);
  not i86062(x86062, x59488);
  not i86063(x86063, x59489);
  not i86064(x86064, x59508);
  not i86065(x86065, x59517);
  not i86066(x86066, x59518);
  not i86067(x86067, x59525);
  not i86068(x86068, x59532);
  not i86069(x86069, x59535);
  not i86070(x86070, x59536);
  not i86071(x86071, x59547);
  not i86072(x86072, x59548);
  not i86073(x86073, x59567);
  not i86074(x86074, x59576);
  not i86075(x86075, x59577);
  not i86076(x86076, x59584);
  not i86077(x86077, x59591);
  not i86078(x86078, x59594);
  not i86079(x86079, x59595);
  not i86080(x86080, x59606);
  not i86081(x86081, x59607);
  not i86082(x86082, x59626);
  not i86083(x86083, x59635);
  not i86084(x86084, x59636);
  not i86085(x86085, x59643);
  not i86086(x86086, x59650);
  not i86087(x86087, x59653);
  not i86088(x86088, x59654);
  not i86089(x86089, x59665);
  not i86090(x86090, x59666);
  not i86091(x86091, x59685);
  not i86092(x86092, x59694);
  not i86093(x86093, x59695);
  not i86094(x86094, x59702);
  not i86095(x86095, x59709);
  not i86096(x86096, x59712);
  not i86097(x86097, x59713);
  not i86098(x86098, x59724);
  not i86099(x86099, x59725);
  not i86100(x86100, x59744);
  not i86101(x86101, x59753);
  not i86102(x86102, x59754);
  not i86103(x86103, x59761);
  not i86104(x86104, x59768);
  not i86105(x86105, x59771);
  not i86106(x86106, x59772);
  not i86107(x86107, x59783);
  not i86108(x86108, x59784);
  not i86109(x86109, x59803);
  not i86110(x86110, x59812);
  not i86111(x86111, x59813);
  not i86112(x86112, x59820);
  not i86113(x86113, x59827);
  not i86114(x86114, x59830);
  not i86115(x86115, x59831);
  not i86116(x86116, x59842);
  not i86117(x86117, x59843);
  not i86118(x86118, x59862);
  not i86119(x86119, x59871);
  not i86120(x86120, x59872);
  not i86121(x86121, x59879);
  not i86122(x86122, x59886);
  not i86123(x86123, x59889);
  not i86124(x86124, x59890);
  not i86125(x86125, x59901);
  not i86126(x86126, x59902);
  not i86127(x86127, x59921);
  not i86128(x86128, x59930);
  not i86129(x86129, x59931);
  not i86130(x86130, x59938);
  not i86131(x86131, x59945);
  not i86132(x86132, x59948);
  not i86133(x86133, x59949);
  not i86134(x86134, x59960);
  not i86135(x86135, x59961);
  not i86136(x86136, x59980);
  not i86137(x86137, x59989);
  not i86138(x86138, x59990);
  not i86139(x86139, x59997);
  not i86140(x86140, x60004);
  not i86141(x86141, x60007);
  not i86142(x86142, x60008);
  not i86143(x86143, x60019);
  not i86144(x86144, x60020);
  not i86145(x86145, x60039);
  not i86146(x86146, x60048);
  not i86147(x86147, x60049);
  not i86148(x86148, x60056);
  not i86149(x86149, x60063);
  not i86150(x86150, x60066);
  not i86151(x86151, x60067);
  not i86152(x86152, x60078);
  not i86153(x86153, x60079);
  not i86154(x86154, x60098);
  not i86155(x86155, x60107);
  not i86156(x86156, x60108);
  not i86157(x86157, x60115);
  not i86158(x86158, x60122);
  not i86159(x86159, x60125);
  not i86160(x86160, x60126);
  not i86161(x86161, x60137);
  not i86162(x86162, x60138);
  not i86163(x86163, x60157);
  not i86164(x86164, x60166);
  not i86165(x86165, x60167);
  not i86166(x86166, x60174);
  not i86167(x86167, x60181);
  not i86168(x86168, x60184);
  not i86169(x86169, x60185);
  not i86170(x86170, x60196);
  not i86171(x86171, x60197);
  not i86172(x86172, x60216);
  not i86173(x86173, x60225);
  not i86174(x86174, x60226);
  not i86175(x86175, x60233);
  not i86176(x86176, x60240);
  not i86177(x86177, x60243);
  not i86178(x86178, x60244);
  not i86179(x86179, x60255);
  not i86180(x86180, x60256);
  not i86181(x86181, x60275);
  not i86182(x86182, x60284);
  not i86183(x86183, x60285);
  not i86184(x86184, x60292);
  not i86185(x86185, x60299);
  not i86186(x86186, x60302);
  not i86187(x86187, x60303);
  not i86188(x86188, x60314);
  not i86189(x86189, x60315);
  not i86190(x86190, x60334);
  not i86191(x86191, x60343);
  not i86192(x86192, x60344);
  not i86193(x86193, x60351);
  not i86194(x86194, x60358);
  not i86195(x86195, x60361);
  not i86196(x86196, x60362);
  not i86197(x86197, x60373);
  not i86198(x86198, x60374);
  not i86199(x86199, x60393);
  not i86200(x86200, x60402);
  not i86201(x86201, x60403);
  not i86202(x86202, x60410);
  not i86203(x86203, x60417);
  not i86204(x86204, x60420);
  not i86205(x86205, x60421);
  not i86206(x86206, x60432);
  not i86207(x86207, x60433);
  not i86208(x86208, x60452);
  not i86209(x86209, x60461);
  not i86210(x86210, x60462);
  not i86211(x86211, x60469);
  not i86212(x86212, x60476);
  not i86213(x86213, x60479);
  not i86214(x86214, x60480);
  not i86215(x86215, x60491);
  not i86216(x86216, x60492);
  not i86217(x86217, x60511);
  not i86218(x86218, x60520);
  not i86219(x86219, x60521);
  not i86220(x86220, x60528);
  not i86221(x86221, x60535);
  not i86222(x86222, x60538);
  not i86223(x86223, x60539);
  not i86224(x86224, x60550);
  not i86225(x86225, x60551);
  not i86226(x86226, x60570);
  not i86227(x86227, x60579);
  not i86228(x86228, x60580);
  not i86229(x86229, x60587);
  not i86230(x86230, x60594);
  not i86231(x86231, x60597);
  not i86232(x86232, x60598);
  not i86233(x86233, x60609);
  not i86234(x86234, x60610);
  not i86235(x86235, x60629);
  not i86236(x86236, x60638);
  not i86237(x86237, x60639);
  not i86238(x86238, x60646);
  not i86239(x86239, x60945);
  not i86240(x86240, x60956);
  not i86241(x86241, x60960);
  not i86242(x86242, x60965);
  not i86243(x86243, x60971);
  not i86244(x86244, x60972);
  not i86245(x86245, x61078);
  not i86246(x86246, x61088);
  not i86247(x86247, x61092);
  not i86248(x86248, x61096);
  not i86249(x86249, x61100);
  not i86250(x86250, x61101);
  not i86251(x86251, x61207);
  not i86252(x86252, x61217);
  not i86253(x86253, x61221);
  not i86254(x86254, x61225);
  not i86255(x86255, x61229);
  not i86256(x86256, x61230);
  not i86257(x86257, x61336);
  not i86258(x86258, x61346);
  not i86259(x86259, x61350);
  not i86260(x86260, x61354);
  not i86261(x86261, x61358);
  not i86262(x86262, x61359);
  not i86263(x86263, x62872);
  not i86264(x86264, x63030);
  not i86265(x86265, x63753);
  not i86266(x86266, x64007);
  not i86267(x86267, x64099);
  not i86268(x86268, x64100);
  not i86269(x86269, x64186);
  not i86270(x86270, x64187);
  not i86271(x86271, x64188);
  not i86272(x86272, x64189);
  not i86273(x86273, x64263);
  not i86274(x86274, x64264);
  not i86275(x86275, x64265);
  not i86276(x86276, x64266);
  not i86277(x86277, x64267);
  not i86278(x86278, x64268);
  not i86279(x86279, x64269);
  not i86280(x86280, x64270);
  not i86281(x86281, x64320);
  not i86282(x86282, x64321);
  not i86283(x86283, x64322);
  not i86284(x86284, x64323);
  not i86285(x86285, x64324);
  not i86286(x86286, x64325);
  not i86287(x86287, x64326);
  not i86288(x86288, x64327);
  not i86289(x86289, x64328);
  not i86290(x86290, x64329);
  not i86291(x86291, x64330);
  not i86292(x86292, x64331);
  not i86293(x86293, x64332);
  not i86294(x86294, x64333);
  not i86295(x86295, x64334);
  not i86296(x86296, x64335);
  not i86297(x86297, x64431);
  not i86298(x86298, x64570);
  not i86299(x86299, x64739);
  not i86300(x86300, x64831);
  not i86301(x86301, x64832);
  not i86302(x86302, x64918);
  not i86303(x86303, x64919);
  not i86304(x86304, x64920);
  not i86305(x86305, x64921);
  not i86306(x86306, x64995);
  not i86307(x86307, x64996);
  not i86308(x86308, x64997);
  not i86309(x86309, x64998);
  not i86310(x86310, x64999);
  not i86311(x86311, x65000);
  not i86312(x86312, x65001);
  not i86313(x86313, x65002);
  not i86314(x86314, x65052);
  not i86315(x86315, x65053);
  not i86316(x86316, x65054);
  not i86317(x86317, x65055);
  not i86318(x86318, x65056);
  not i86319(x86319, x65057);
  not i86320(x86320, x65058);
  not i86321(x86321, x65059);
  not i86322(x86322, x65060);
  not i86323(x86323, x65061);
  not i86324(x86324, x65062);
  not i86325(x86325, x65063);
  not i86326(x86326, x65064);
  not i86327(x86327, x65065);
  not i86328(x86328, x65066);
  not i86329(x86329, x65067);
  not i86330(x86330, x65101);
  not i86331(x86331, x65240);
  not i86332(x86332, x65409);
  not i86333(x86333, x65501);
  not i86334(x86334, x65502);
  not i86335(x86335, x65588);
  not i86336(x86336, x65589);
  not i86337(x86337, x65590);
  not i86338(x86338, x65591);
  not i86339(x86339, x65665);
  not i86340(x86340, x65666);
  not i86341(x86341, x65667);
  not i86342(x86342, x65668);
  not i86343(x86343, x65669);
  not i86344(x86344, x65670);
  not i86345(x86345, x65671);
  not i86346(x86346, x65672);
  not i86347(x86347, x65722);
  not i86348(x86348, x65723);
  not i86349(x86349, x65724);
  not i86350(x86350, x65725);
  not i86351(x86351, x65726);
  not i86352(x86352, x65727);
  not i86353(x86353, x65728);
  not i86354(x86354, x65729);
  not i86355(x86355, x65730);
  not i86356(x86356, x65731);
  not i86357(x86357, x65732);
  not i86358(x86358, x65733);
  not i86359(x86359, x65734);
  not i86360(x86360, x65735);
  not i86361(x86361, x65736);
  not i86362(x86362, x65737);
  not i86363(x86363, x65771);
  not i86364(x86364, x65910);
  not i86365(x86365, x66079);
  not i86366(x86366, x66171);
  not i86367(x86367, x66172);
  not i86368(x86368, x66258);
  not i86369(x86369, x66259);
  not i86370(x86370, x66260);
  not i86371(x86371, x66261);
  not i86372(x86372, x66335);
  not i86373(x86373, x66336);
  not i86374(x86374, x66337);
  not i86375(x86375, x66338);
  not i86376(x86376, x66339);
  not i86377(x86377, x66340);
  not i86378(x86378, x66341);
  not i86379(x86379, x66342);
  not i86380(x86380, x66392);
  not i86381(x86381, x66393);
  not i86382(x86382, x66394);
  not i86383(x86383, x66395);
  not i86384(x86384, x66396);
  not i86385(x86385, x66397);
  not i86386(x86386, x66398);
  not i86387(x86387, x66399);
  not i86388(x86388, x66400);
  not i86389(x86389, x66401);
  not i86390(x86390, x66402);
  not i86391(x86391, x66403);
  not i86392(x86392, x66404);
  not i86393(x86393, x66405);
  not i86394(x86394, x66406);
  not i86395(x86395, x66407);
  not i86396(x86396, x67404);
  not i86397(x86397, x68397);
  not i86398(x86398, x68531);
  not i86399(x86399, x68538);
  not i86400(x86400, x68539);
  not i86401(x86401, x68542);
  not i86402(x86402, x68664);
  not i86403(x86403, x68666);
  not i86404(x86404, x68685);
  not i86405(x86405, x68687);
  not i86406(x86406, x68704);
  not i86407(x86407, x68705);
  not i86408(x86408, x68706);
  not i86409(x86409, x68707);
  not i86410(x86410, x68722);
  not i86411(x86411, x68723);
  not i86412(x86412, x68724);
  not i86413(x86413, x68725);
  not i86414(x86414, x68754);
  not i86415(x86415, x68770);
  not i86416(x86416, x68786);
  not i86417(x86417, x68802);
  not i86418(x86418, x68819);
  not i86419(x86419, x68835);
  not i86420(x86420, x68851);
  not i86421(x86421, x68867);
  not i86422(x86422, x68883);
  not i86423(x86423, x68896);
  not i86424(x86424, x68897);
  not i86425(x86425, x68910);
  not i86426(x86426, x68911);
  not i86427(x86427, x68924);
  not i86428(x86428, x68925);
  not i86429(x86429, x68938);
  not i86430(x86430, x68939);
  not i86431(x86431, x68952);
  not i86432(x86432, x68953);
  not i86433(x86433, x68966);
  not i86434(x86434, x68967);
  not i86435(x86435, x68980);
  not i86436(x86436, x68981);
  not i86437(x86437, x68994);
  not i86438(x86438, x68995);
  not i86439(x86439, x69008);
  not i86440(x86440, x69009);
  not i86441(x86441, x69022);
  not i86442(x86442, x69023);
  not i86443(x86443, x69036);
  not i86444(x86444, x69037);
  not i86445(x86445, x69050);
  not i86446(x86446, x69051);
  not i86447(x86447, x69064);
  not i86448(x86448, x69065);
  not i86449(x86449, x69078);
  not i86450(x86450, x69079);
  not i86451(x86451, x69092);
  not i86452(x86452, x69093);
  not i86453(x86453, x69106);
  not i86454(x86454, x69107);
  not i86455(x86455, x69120);
  not i86456(x86456, x69121);
  not i86457(x86457, x69134);
  not i86458(x86458, x69135);
  not i86459(x86459, x69148);
  not i86460(x86460, x69149);
  not i86461(x86461, x69162);
  not i86462(x86462, x69163);
  not i86463(x86463, x69176);
  not i86464(x86464, x69177);
  not i86465(x86465, x69190);
  not i86466(x86466, x69191);
  not i86467(x86467, x69204);
  not i86468(x86468, x69205);
  not i86469(x86469, x69218);
  not i86470(x86470, x69219);
  not i86471(x86471, x69232);
  not i86472(x86472, x69233);
  not i86473(x86473, x69246);
  not i86474(x86474, x69247);
  not i86475(x86475, x69260);
  not i86476(x86476, x69261);
  not i86477(x86477, x69274);
  not i86478(x86478, x69275);
  not i86479(x86479, x69288);
  not i86480(x86480, x69289);
  not i86481(x86481, x69302);
  not i86482(x86482, x69303);
  not i86483(x86483, x69316);
  not i86484(x86484, x69317);
  not i86485(x86485, x69333);
  not i86486(x86486, x69346);
  not i86487(x86487, x69347);
  not i86488(x86488, x69360);
  not i86489(x86489, x69361);
  not i86490(x86490, x69374);
  not i86491(x86491, x69375);
  not i86492(x86492, x69388);
  not i86493(x86493, x69389);
  not i86494(x86494, x69402);
  not i86495(x86495, x69403);
  not i86496(x86496, x69416);
  not i86497(x86497, x69417);
  not i86498(x86498, x69430);
  not i86499(x86499, x69431);
  not i86500(x86500, x69444);
  not i86501(x86501, x69445);
  not i86502(x86502, x69458);
  not i86503(x86503, x69459);
  not i86504(x86504, x69472);
  not i86505(x86505, x69473);
  not i86506(x86506, x69486);
  not i86507(x86507, x69487);
  not i86508(x86508, x69500);
  not i86509(x86509, x69501);
  not i86510(x86510, x69514);
  not i86511(x86511, x69515);
  not i86512(x86512, x69528);
  not i86513(x86513, x69529);
  not i86514(x86514, x69542);
  not i86515(x86515, x69543);
  not i86516(x86516, x69556);
  not i86517(x86517, x69557);
  not i86518(x86518, x69570);
  not i86519(x86519, x69571);
  not i86520(x86520, x69584);
  not i86521(x86521, x69585);
  not i86522(x86522, x69598);
  not i86523(x86523, x69599);
  not i86524(x86524, x69612);
  not i86525(x86525, x69613);
  not i86526(x86526, x69626);
  not i86527(x86527, x69627);
  not i86528(x86528, x69640);
  not i86529(x86529, x69641);
  not i86530(x86530, x69654);
  not i86531(x86531, x69655);
  not i86532(x86532, x69668);
  not i86533(x86533, x69669);
  not i86534(x86534, x69682);
  not i86535(x86535, x69683);
  not i86536(x86536, x69696);
  not i86537(x86537, x69697);
  not i86538(x86538, x69710);
  not i86539(x86539, x69711);
  not i86540(x86540, x69724);
  not i86541(x86541, x69725);
  not i86542(x86542, x69738);
  not i86543(x86543, x69739);
  not i86544(x86544, x69752);
  not i86545(x86545, x69753);
  not i86546(x86546, x69766);
  not i86547(x86547, x69767);
  not i86548(x86548, x69783);
  not i86549(x86549, x69796);
  not i86550(x86550, x69797);
  not i86551(x86551, x69810);
  not i86552(x86552, x69811);
  not i86553(x86553, x69824);
  not i86554(x86554, x69825);
  not i86555(x86555, x69838);
  not i86556(x86556, x69839);
  not i86557(x86557, x69852);
  not i86558(x86558, x69853);
  not i86559(x86559, x69866);
  not i86560(x86560, x69867);
  not i86561(x86561, x69880);
  not i86562(x86562, x69881);
  not i86563(x86563, x69894);
  not i86564(x86564, x69895);
  not i86565(x86565, x69908);
  not i86566(x86566, x69909);
  not i86567(x86567, x69922);
  not i86568(x86568, x69923);
  not i86569(x86569, x69936);
  not i86570(x86570, x69937);
  not i86571(x86571, x69950);
  not i86572(x86572, x69951);
  not i86573(x86573, x69964);
  not i86574(x86574, x69965);
  not i86575(x86575, x69978);
  not i86576(x86576, x69979);
  not i86577(x86577, x69992);
  not i86578(x86578, x69993);
  not i86579(x86579, x70006);
  not i86580(x86580, x70007);
  not i86581(x86581, x70020);
  not i86582(x86582, x70021);
  not i86583(x86583, x70034);
  not i86584(x86584, x70035);
  not i86585(x86585, x70048);
  not i86586(x86586, x70049);
  not i86587(x86587, x70062);
  not i86588(x86588, x70063);
  not i86589(x86589, x70076);
  not i86590(x86590, x70077);
  not i86591(x86591, x70090);
  not i86592(x86592, x70091);
  not i86593(x86593, x70104);
  not i86594(x86594, x70105);
  not i86595(x86595, x70118);
  not i86596(x86596, x70119);
  not i86597(x86597, x70132);
  not i86598(x86598, x70133);
  not i86599(x86599, x70146);
  not i86600(x86600, x70147);
  not i86601(x86601, x70160);
  not i86602(x86602, x70161);
  not i86603(x86603, x70174);
  not i86604(x86604, x70175);
  not i86605(x86605, x70188);
  not i86606(x86606, x70189);
  not i86607(x86607, x70202);
  not i86608(x86608, x70203);
  not i86609(x86609, x70216);
  not i86610(x86610, x70217);
  not i86611(x86611, x70233);
  not i86612(x86612, x70246);
  not i86613(x86613, x70247);
  not i86614(x86614, x70260);
  not i86615(x86615, x70261);
  not i86616(x86616, x70274);
  not i86617(x86617, x70275);
  not i86618(x86618, x70288);
  not i86619(x86619, x70289);
  not i86620(x86620, x70302);
  not i86621(x86621, x70303);
  not i86622(x86622, x70316);
  not i86623(x86623, x70317);
  not i86624(x86624, x70330);
  not i86625(x86625, x70331);
  not i86626(x86626, x70344);
  not i86627(x86627, x70345);
  not i86628(x86628, x70358);
  not i86629(x86629, x70359);
  not i86630(x86630, x70372);
  not i86631(x86631, x70373);
  not i86632(x86632, x70386);
  not i86633(x86633, x70387);
  not i86634(x86634, x70400);
  not i86635(x86635, x70401);
  not i86636(x86636, x70414);
  not i86637(x86637, x70415);
  not i86638(x86638, x70428);
  not i86639(x86639, x70429);
  not i86640(x86640, x70442);
  not i86641(x86641, x70443);
  not i86642(x86642, x70456);
  not i86643(x86643, x70457);
  not i86644(x86644, x70470);
  not i86645(x86645, x70471);
  not i86646(x86646, x70484);
  not i86647(x86647, x70485);
  not i86648(x86648, x70498);
  not i86649(x86649, x70499);
  not i86650(x86650, x70512);
  not i86651(x86651, x70513);
  not i86652(x86652, x70526);
  not i86653(x86653, x70527);
  not i86654(x86654, x70540);
  not i86655(x86655, x70541);
  not i86656(x86656, x70554);
  not i86657(x86657, x70555);
  not i86658(x86658, x70568);
  not i86659(x86659, x70569);
  not i86660(x86660, x70582);
  not i86661(x86661, x70583);
  not i86662(x86662, x70596);
  not i86663(x86663, x70597);
  not i86664(x86664, x70610);
  not i86665(x86665, x70611);
  not i86666(x86666, x70624);
  not i86667(x86667, x70625);
  not i86668(x86668, x70638);
  not i86669(x86669, x70639);
  not i86670(x86670, x70652);
  not i86671(x86671, x70653);
  not i86672(x86672, x70666);
  not i86673(x86673, x70667);
  not i86674(x86674, x70683);
  not i86675(x86675, x70699);
  not i86676(x86676, x70715);
  not i86677(x86677, x70731);
  not i86678(x86678, x70747);
  not i86679(x86679, x70763);
  not i86680(x86680, x70779);
  not i86681(x86681, x70795);
  not i86682(x86682, x70811);
  not i86683(x86683, x70827);
  not i86684(x86684, x70843);
  not i86685(x86685, x70859);
  not i86686(x86686, x70875);
  not i86687(x86687, x70891);
  not i86688(x86688, x70907);
  not i86689(x86689, x70923);
  not i86690(x86690, x70939);
  not i86691(x86691, x70955);
  not i86692(x86692, x70971);
  not i86693(x86693, x70987);
  not i86694(x86694, x71003);
  not i86695(x86695, x71019);
  not i86696(x86696, x71143);
  not i86697(x86697, x71148);
  not i86698(x86698, x71153);
  not i86699(x86699, x71158);
  not i86700(x86700, x71163);
  not i86701(x86701, x71168);
  not i86702(x86702, x71173);
  not i86703(x86703, x71178);
  not i86704(x86704, x71198);
  not i86705(x86705, x71206);
  not i86706(x86706, x71211);
  not i86707(x86707, x71216);
  not i86708(x86708, x71221);
  not i86709(x86709, x71226);
  not i86710(x86710, x71231);
  not i86711(x86711, x71236);
  not i86712(x86712, x71241);
  not i86713(x86713, x71246);
  not i86714(x86714, x71251);
  not i86715(x86715, x71256);
  not i86716(x86716, x71261);
  not i86717(x86717, x71266);
  not i86718(x86718, x71271);
  not i86719(x86719, x71276);
  not i86720(x86720, x71278);
  not i86721(x86721, x71280);
  not i86722(x86722, x71285);
  not i86723(x86723, x71290);
  not i86724(x86724, x71295);
  not i86725(x86725, x71300);
  not i86726(x86726, x71305);
  not i86727(x86727, x71310);
  not i86728(x86728, x71315);
  not i86729(x86729, x71320);
  not i86730(x86730, x71325);
  not i86731(x86731, x71330);
  not i86732(x86732, x71335);
  not i86733(x86733, x71340);
  not i86734(x86734, x71345);
  not i86735(x86735, x71350);
  not i86736(x86736, x71355);
  not i86737(x86737, x71360);
  not i86738(x86738, x71365);
  not i86739(x86739, x71370);
  not i86740(x86740, x71375);
  not i86741(x86741, x71380);
  not i86742(x86742, x71385);
  not i86743(x86743, x71390);
  not i86744(x86744, x71395);
  not i86745(x86745, x71400);
  not i86746(x86746, x71405);
  not i86747(x86747, x71410);
  not i86748(x86748, x71415);
  not i86749(x86749, x71420);
  not i86750(x86750, x71425);
  not i86751(x86751, x71430);
  not i86752(x86752, x71435);
  not i86753(x86753, x71440);
  not i86754(x86754, x71445);
  not i86755(x86755, x71450);
  not i86756(x86756, x71455);
  not i86757(x86757, x71460);
  not i86758(x86758, x71465);
  not i86759(x86759, x71470);
  not i86760(x86760, x71475);
  not i86761(x86761, x71486);
  not i86762(x86762, x71491);
  not i86763(x86763, x71496);
  not i86764(x86764, x71501);
  not i86765(x86765, x71506);
  not i86766(x86766, x71511);
  not i86767(x86767, x71516);
  not i86768(x86768, x71521);
  not i86769(x86769, x71526);
  not i86770(x86770, x71531);
  not i86771(x86771, x71536);
  not i86772(x86772, x71541);
  not i86773(x86773, x71546);
  not i86774(x86774, x71551);
  not i86775(x86775, x71556);
  not i86776(x86776, x71561);
  not i86777(x86777, x71566);
  not i86778(x86778, x71571);
  not i86779(x86779, x71576);
  not i86780(x86780, x71581);
  not i86781(x86781, x71586);
  not i86782(x86782, x71591);
  not i86783(x86783, x71596);
  not i86784(x86784, x71601);
  not i86785(x86785, x71606);
  not i86786(x86786, x71611);
  not i86787(x86787, x71616);
  not i86788(x86788, x71621);
  not i86789(x86789, x71626);
  not i86790(x86790, x71631);
  not i86791(x86791, x71638);
  not i86792(x86792, x71643);
  not i86793(x86793, x71648);
  not i86794(x86794, x71653);
  not i86795(x86795, x71658);
  not i86796(x86796, x71663);
  not i86797(x86797, x71668);
  not i86798(x86798, x71673);
  not i86799(x86799, x71678);
  not i86800(x86800, x71683);
  not i86801(x86801, x71688);
  not i86802(x86802, x71693);
  not i86803(x86803, x71698);
  not i86804(x86804, x71703);
  not i86805(x86805, x71708);
  not i86806(x86806, x71713);
  not i86807(x86807, x71718);
  not i86808(x86808, x71723);
  not i86809(x86809, x71728);
  not i86810(x86810, x71733);
  not i86811(x86811, x71738);
  not i86812(x86812, x71743);
  not i86813(x86813, x71748);
  not i86814(x86814, x71753);
  not i86815(x86815, x71758);
  not i86816(x86816, x71763);
  not i86817(x86817, x71768);
  not i86818(x86818, x71773);
  not i86819(x86819, x71778);
  not i86820(x86820, x71783);
  not i86821(x86821, x71788);
  not i86822(x86822, x71793);
  not i86823(x86823, x71798);
  not i86824(x86824, x71803);
  not i86825(x86825, x71808);
  not i86826(x86826, x71813);
  not i86827(x86827, x71818);
  not i86828(x86828, x71823);
  not i86829(x86829, x71828);
  not i86830(x86830, x71833);
  not i86831(x86831, x71838);
  not i86832(x86832, x71843);
  not i86833(x86833, x71848);
  not i86834(x86834, x71853);
  not i86835(x86835, x71858);
  not i86836(x86836, x71863);
  not i86837(x86837, x71868);
  not i86838(x86838, x71873);
  not i86839(x86839, x71878);
  not i86840(x86840, x71883);
  not i86841(x86841, x71888);
  not i86842(x86842, x71893);
  not i86843(x86843, x71898);
  not i86844(x86844, x71903);
  not i86845(x86845, x71938);
  not i86846(x86846, x71943);
  not i86847(x86847, x71948);
  not i86848(x86848, x71953);
  not i86849(x86849, x71958);
  not i86850(x86850, x71963);
  not i86851(x86851, x71968);
  not i86852(x86852, x71973);
  not i86853(x86853, x71978);
  not i86854(x86854, x71983);
  not i86855(x86855, x71988);
  not i86856(x86856, x71993);
  not i86857(x86857, x71998);
  not i86858(x86858, x72003);
  not i86859(x86859, x72008);
  not i86860(x86860, x72013);
  not i86861(x86861, x72018);
  not i86862(x86862, x72023);
  not i86863(x86863, x72028);
  not i86864(x86864, x72033);
  not i86865(x86865, x72038);
  not i86866(x86866, x72043);
  not i86867(x86867, x72048);
  not i86868(x86868, x72053);
  not i86869(x86869, x72058);
  not i86870(x86870, x72063);
  not i86871(x86871, x72068);
  not i86872(x86872, x72073);
  not i86873(x86873, x72078);
  not i86874(x86874, x72083);
  not i86875(x86875, x72088);
  not i86876(x86876, x72093);
  not i86877(x86877, x72098);
  not i86878(x86878, x72103);
  not i86879(x86879, x72108);
  not i86880(x86880, x72113);
  not i86881(x86881, x72118);
  not i86882(x86882, x72123);
  not i86883(x86883, x72128);
  not i86884(x86884, x72133);
  not i86885(x86885, x72138);
  not i86886(x86886, x72143);
  not i86887(x86887, x72148);
  not i86888(x86888, x72153);
  not i86889(x86889, x72158);
  not i86890(x86890, x72163);
  not i86891(x86891, x72168);
  not i86892(x86892, x72173);
  not i86893(x86893, x72178);
  not i86894(x86894, x72183);
  not i86895(x86895, x72188);
  not i86896(x86896, x72193);
  not i86897(x86897, x72198);
  not i86898(x86898, x72203);
  not i86899(x86899, x72208);
  not i86900(x86900, x72213);
  not i86901(x86901, x72218);
  not i86902(x86902, x72223);
  not i86903(x86903, x72228);
  not i86904(x86904, x72233);
  not i86905(x86905, x72238);
  not i86906(x86906, x72243);
  not i86907(x86907, x72248);
  not i86908(x86908, x72253);
  not i86909(x86909, x72258);
  not i86910(x86910, x72263);
  not i86911(x86911, x72268);
  not i86912(x86912, x72273);
  not i86913(x86913, x72278);
  not i86914(x86914, x72283);
  not i86915(x86915, x72288);
  not i86916(x86916, x72293);
  not i86917(x86917, x72298);
  not i86918(x86918, x72303);
  not i86919(x86919, x72308);
  not i86920(x86920, x72313);
  not i86921(x86921, x72318);
  not i86922(x86922, x72323);
  not i86923(x86923, x72328);
  not i86924(x86924, x72333);
  not i86925(x86925, x72338);
  not i86926(x86926, x72343);
  not i86927(x86927, x72348);
  not i86928(x86928, x72353);
  not i86929(x86929, x72358);
  not i86930(x86930, x72363);
  not i86931(x86931, x72368);
  not i86932(x86932, x72373);
  not i86933(x86933, x72378);
  not i86934(x86934, x72383);
  not i86935(x86935, x72388);
  not i86936(x86936, x72393);
  not i86937(x86937, x72398);
  not i86938(x86938, x72403);
  not i86939(x86939, x72408);
  not i86940(x86940, x72413);
  not i86941(x86941, x72418);
  not i86942(x86942, x72423);
  not i86943(x86943, x72428);
  not i86944(x86944, x72433);
  not i86945(x86945, x72438);
  not i86946(x86946, x72443);
  not i86947(x86947, x72448);
  not i86948(x86948, x72453);
  not i86949(x86949, x72458);
  not i86950(x86950, x72463);
  not i86951(x86951, x72468);
  not i86952(x86952, x72473);
  not i86953(x86953, x72478);
  not i86954(x86954, x72483);
  not i86955(x86955, x72488);
  not i86956(x86956, x72493);
  not i86957(x86957, x72498);
  not i86958(x86958, x72503);
  not i86959(x86959, x72508);
  not i86960(x86960, x72513);
  not i86961(x86961, x72518);
  not i86962(x86962, x72523);
  not i86963(x86963, x72528);
  not i86964(x86964, x72533);
  not i86965(x86965, x72538);
  not i86966(x86966, x72543);
  not i86967(x86967, x72548);
  not i86968(x86968, x72553);
  not i86969(x86969, x72558);
  not i86970(x86970, x72563);
  not i86971(x86971, x72568);
  not i86972(x86972, x72573);
  not i86973(x86973, x72578);
  not i86974(x86974, x72583);
  not i86975(x86975, x72588);
  not i86976(x86976, x72593);
  not i86977(x86977, x72598);
  not i86978(x86978, x72603);
  not i86979(x86979, x72608);
  not i86980(x86980, x72613);
  not i86981(x86981, x72618);
  not i86982(x86982, x72623);
  not i86983(x86983, x72628);
  not i86984(x86984, x72633);
  not i86985(x86985, x72638);
  not i86986(x86986, x72643);
  not i86987(x86987, x72648);
  not i86988(x86988, x72653);
  not i86989(x86989, x72658);
  not i86990(x86990, x72663);
  not i86991(x86991, x72668);
  not i86992(x86992, x72673);
  not i86993(x86993, x72678);
  not i86994(x86994, x72683);
  not i86995(x86995, x72688);
  not i86996(x86996, x72693);
  not i86997(x86997, x72698);
  not i86998(x86998, x72703);
  not i86999(x86999, x72708);
  not i87000(x87000, x72713);
  not i87001(x87001, x72718);
  not i87002(x87002, x72723);
  not i87003(x87003, x72728);
  not i87004(x87004, x72733);
  not i87005(x87005, x72738);
  not i87006(x87006, x72743);
  not i87007(x87007, x72748);
  not i87008(x87008, x72753);
  not i87009(x87009, x72758);
  not i87010(x87010, x72763);
  not i87011(x87011, x72768);
  not i87012(x87012, x72773);
  not i87013(x87013, x72778);
  not i87014(x87014, x72783);
  not i87015(x87015, x72788);
  not i87016(x87016, x72793);
  not i87017(x87017, x72798);
  not i87018(x87018, x72803);
  not i87019(x87019, x72808);
  not i87020(x87020, x72813);
  not i87021(x87021, x72818);
  not i87022(x87022, x72823);
  not i87023(x87023, x72828);
  not i87024(x87024, x72833);
  not i87025(x87025, x72838);
  not i87026(x87026, x72843);
  not i87027(x87027, x72848);
  not i87028(x87028, x72853);
  not i87029(x87029, x72858);
  not i87030(x87030, x72863);
  not i87031(x87031, x72868);
  not i87032(x87032, x72873);
  not i87033(x87033, x72878);
  not i87034(x87034, x72883);
  not i87035(x87035, x72888);
  not i87036(x87036, x72893);
  not i87037(x87037, x72898);
  not i87038(x87038, x72903);
  not i87039(x87039, x72908);
  not i87040(x87040, x72913);
  not i87041(x87041, x72918);
  not i87042(x87042, x72923);
  not i87043(x87043, x72928);
  not i87044(x87044, x72933);
  not i87045(x87045, x72938);
  not i87046(x87046, x72943);
  not i87047(x87047, x72948);
  not i87048(x87048, x72953);
  not i87049(x87049, x72958);
  not i87050(x87050, x72963);
  not i87051(x87051, x72968);
  not i87052(x87052, x72973);
  not i87053(x87053, x72978);
  not i87054(x87054, x72983);
  not i87055(x87055, x72988);
  not i87056(x87056, x72993);
  not i87057(x87057, x72998);
  not i87058(x87058, x73003);
  not i87059(x87059, x73008);
  not i87060(x87060, x73013);
  not i87061(x87061, x73018);
  not i87062(x87062, x73023);
  not i87063(x87063, x73028);
  not i87064(x87064, x73033);
  not i87065(x87065, x73038);
  not i87066(x87066, x73043);
  not i87067(x87067, x73048);
  not i87068(x87068, x73053);
  not i87069(x87069, x73058);
  not i87070(x87070, x73063);
  not i87071(x87071, x73068);
  not i87072(x87072, x73073);
  not i87073(x87073, x73078);
  not i87074(x87074, x73083);
  not i87075(x87075, x73088);
  not i87076(x87076, x73093);
  not i87077(x87077, x73098);
  not i87078(x87078, x73103);
  not i87079(x87079, x73108);
  not i87080(x87080, x73113);
  not i87081(x87081, x73118);
  not i87082(x87082, x73123);
  not i87083(x87083, x73128);
  not i87084(x87084, x73133);
  not i87085(x87085, x73138);
  not i87086(x87086, x73143);
  not i87087(x87087, x73148);
  not i87088(x87088, x73153);
  not i87089(x87089, x73158);
  not i87090(x87090, x73163);
  not i87091(x87091, x73168);
  not i87092(x87092, x73173);
  not i87093(x87093, x73178);
  not i87094(x87094, x73183);
  not i87095(x87095, x73188);
  not i87096(x87096, x73193);
  not i87097(x87097, x73198);
  not i87098(x87098, x73203);
  not i87099(x87099, x73208);
  not i87100(x87100, x73213);
  not i87101(x87101, x73218);
  not i87102(x87102, x73223);
  not i87103(x87103, x73228);
  not i87104(x87104, x73233);
  not i87105(x87105, x73238);
  not i87106(x87106, x73243);
  not i87107(x87107, x73248);
  not i87108(x87108, x73253);
  not i87109(x87109, x73258);
  not i87110(x87110, x73263);
  not i87111(x87111, x73268);
  not i87112(x87112, x73273);
  not i87113(x87113, x73278);
  not i87114(x87114, x73283);
  not i87115(x87115, x73288);
  not i87116(x87116, x73293);
  not i87117(x87117, x73298);
  not i87118(x87118, x73303);
  not i87119(x87119, x73308);
  not i87120(x87120, x73313);
  not i87121(x87121, x73318);
  not i87122(x87122, x73323);
  not i87123(x87123, x73328);
  not i87124(x87124, x73333);
  not i87125(x87125, x73338);
  not i87126(x87126, x73343);
  not i87127(x87127, x73348);
  not i87128(x87128, x73353);
  not i87129(x87129, x73358);
  not i87130(x87130, x73363);
  not i87131(x87131, x73368);
  not i87132(x87132, x73373);
  not i87133(x87133, x73378);
  not i87134(x87134, x73383);
  not i87135(x87135, x73388);
  not i87136(x87136, x73393);
  not i87137(x87137, x73398);
  not i87138(x87138, x73403);
  not i87139(x87139, x73408);
  not i87140(x87140, x73413);
  not i87141(x87141, x73418);
  not i87142(x87142, x73423);
  not i87143(x87143, x73428);
  not i87144(x87144, x73433);
  not i87145(x87145, x73438);
  not i87146(x87146, x73443);
  not i87147(x87147, x73448);
  not i87148(x87148, x73453);
  not i87149(x87149, x73458);
  not i87150(x87150, x73463);
  not i87151(x87151, x73468);
  not i87152(x87152, x73473);
  not i87153(x87153, x73478);
  not i87154(x87154, x73483);
  not i87155(x87155, x73488);
  not i87156(x87156, x73493);
  not i87157(x87157, x73498);
  not i87158(x87158, x73503);
  not i87159(x87159, x73508);
  not i87160(x87160, x73513);
  not i87161(x87161, x73518);
  not i87162(x87162, x73523);
  not i87163(x87163, x73528);
  not i87164(x87164, x73533);
  not i87165(x87165, x73538);
  not i87166(x87166, x73543);
  not i87167(x87167, x73548);
  not i87168(x87168, x73553);
  not i87169(x87169, x73558);
  not i87170(x87170, x73563);
  not i87171(x87171, x73568);
  not i87172(x87172, x73573);
  not i87173(x87173, x73578);
  not i87174(x87174, x73583);
  not i87175(x87175, x73588);
  not i87176(x87176, x73593);
  not i87177(x87177, x73598);
  not i87178(x87178, x73603);
  not i87179(x87179, x73608);
  not i87180(x87180, x73613);
  not i87181(x87181, x73618);
  not i87182(x87182, x73623);
  not i87183(x87183, x73628);
  not i87184(x87184, x73633);
  not i87185(x87185, x73638);
  not i87186(x87186, x73643);
  not i87187(x87187, x73648);
  not i87188(x87188, x73653);
  not i87189(x87189, x73658);
  not i87190(x87190, x73663);
  not i87191(x87191, x73668);
  not i87192(x87192, x73673);
  not i87193(x87193, x73678);
  not i87194(x87194, x73683);
  not i87195(x87195, x73688);
  not i87196(x87196, x73693);
  not i87197(x87197, x73698);
  not i87198(x87198, x73703);
  not i87199(x87199, x73708);
  not i87200(x87200, x73713);
  not i87201(x87201, x73718);
  not i87202(x87202, x73723);
  not i87203(x87203, x73728);
  not i87204(x87204, x73733);
  not i87205(x87205, x73738);
  not i87206(x87206, x73743);
  not i87207(x87207, x73748);
  not i87208(x87208, x73753);
  not i87209(x87209, x73758);
  not i87210(x87210, x73763);
  not i87211(x87211, x73768);
  not i87212(x87212, x73773);
  not i87213(x87213, x73778);
  not i87214(x87214, x73783);
  not i87215(x87215, x73788);
  not i87216(x87216, x73793);
  not i87217(x87217, x73798);
  not i87218(x87218, x73803);
  not i87219(x87219, x73808);
  not i87220(x87220, x73813);
  not i87221(x87221, x73818);
  not i87222(x87222, x73823);
  not i87223(x87223, x73828);
  not i87224(x87224, x73833);
  not i87225(x87225, x73838);
  not i87226(x87226, x73843);
  not i87227(x87227, x73848);
  not i87228(x87228, x73853);
  not i87229(x87229, x73858);
  not i87230(x87230, x73863);
  not i87231(x87231, x73868);
  not i87232(x87232, x73873);
  not i87233(x87233, x73878);
  not i87234(x87234, x73883);
  not i87235(x87235, x73888);
  not i87236(x87236, x73893);
  not i87237(x87237, x73898);
  not i87238(x87238, x73903);
  not i87239(x87239, x73908);
  not i87240(x87240, x73913);
  not i87241(x87241, x73918);
  not i87242(x87242, x73923);
  not i87243(x87243, x73928);
  not i87244(x87244, x73933);
  not i87245(x87245, x73938);
  not i87246(x87246, x73943);
  not i87247(x87247, x73948);
  not i87248(x87248, x73953);
  not i87249(x87249, x73958);
  not i87250(x87250, x73963);
  not i87251(x87251, x73968);
  not i87252(x87252, x73973);
  not i87253(x87253, x73978);
  not i87254(x87254, x73983);
  not i87255(x87255, x73988);
  not i87256(x87256, x73993);
  not i87257(x87257, x73998);
  not i87258(x87258, x83348);
  not i87259(x87259, x83353);
  not i87260(x87260, x83358);
  not i87261(x87261, x83363);
  not i87262(x87262, x83368);
  not i87263(x87263, x83373);
  not i87264(x87264, x83378);

  assign x61684 = AluDivFinish;
  assign x61428 = AluDivQ[0];
  assign x61429 = AluDivQ[1];
  assign x61430 = AluDivQ[2];
  assign x61431 = AluDivQ[3];
  assign x61432 = AluDivQ[4];
  assign x61433 = AluDivQ[5];
  assign x61434 = AluDivQ[6];
  assign x61435 = AluDivQ[7];
  assign x61436 = AluDivQ[8];
  assign x61437 = AluDivQ[9];
  assign x61438 = AluDivQ[10];
  assign x61439 = AluDivQ[11];
  assign x61440 = AluDivQ[12];
  assign x61441 = AluDivQ[13];
  assign x61442 = AluDivQ[14];
  assign x61443 = AluDivQ[15];
  assign x61444 = AluDivQ[16];
  assign x61445 = AluDivQ[17];
  assign x61446 = AluDivQ[18];
  assign x61447 = AluDivQ[19];
  assign x61448 = AluDivQ[20];
  assign x61449 = AluDivQ[21];
  assign x61450 = AluDivQ[22];
  assign x61451 = AluDivQ[23];
  assign x61452 = AluDivQ[24];
  assign x61453 = AluDivQ[25];
  assign x61454 = AluDivQ[26];
  assign x61455 = AluDivQ[27];
  assign x61456 = AluDivQ[28];
  assign x61457 = AluDivQ[29];
  assign x61458 = AluDivQ[30];
  assign x61459 = AluDivQ[31];
  assign x61460 = AluDivQ[32];
  assign x61461 = AluDivQ[33];
  assign x61462 = AluDivQ[34];
  assign x61463 = AluDivQ[35];
  assign x61464 = AluDivQ[36];
  assign x61465 = AluDivQ[37];
  assign x61466 = AluDivQ[38];
  assign x61467 = AluDivQ[39];
  assign x61468 = AluDivQ[40];
  assign x61469 = AluDivQ[41];
  assign x61470 = AluDivQ[42];
  assign x61471 = AluDivQ[43];
  assign x61472 = AluDivQ[44];
  assign x61473 = AluDivQ[45];
  assign x61474 = AluDivQ[46];
  assign x61475 = AluDivQ[47];
  assign x61476 = AluDivQ[48];
  assign x61477 = AluDivQ[49];
  assign x61478 = AluDivQ[50];
  assign x61479 = AluDivQ[51];
  assign x61480 = AluDivQ[52];
  assign x61481 = AluDivQ[53];
  assign x61482 = AluDivQ[54];
  assign x61483 = AluDivQ[55];
  assign x61484 = AluDivQ[56];
  assign x61485 = AluDivQ[57];
  assign x61486 = AluDivQ[58];
  assign x61487 = AluDivQ[59];
  assign x61488 = AluDivQ[60];
  assign x61489 = AluDivQ[61];
  assign x61490 = AluDivQ[62];
  assign x61491 = AluDivQ[63];
  assign x61492 = AluDivQ[64];
  assign x61493 = AluDivQ[65];
  assign x61494 = AluDivQ[66];
  assign x61495 = AluDivQ[67];
  assign x61496 = AluDivQ[68];
  assign x61497 = AluDivQ[69];
  assign x61498 = AluDivQ[70];
  assign x61499 = AluDivQ[71];
  assign x61500 = AluDivQ[72];
  assign x61501 = AluDivQ[73];
  assign x61502 = AluDivQ[74];
  assign x61503 = AluDivQ[75];
  assign x61504 = AluDivQ[76];
  assign x61505 = AluDivQ[77];
  assign x61506 = AluDivQ[78];
  assign x61507 = AluDivQ[79];
  assign x61508 = AluDivQ[80];
  assign x61509 = AluDivQ[81];
  assign x61510 = AluDivQ[82];
  assign x61511 = AluDivQ[83];
  assign x61512 = AluDivQ[84];
  assign x61513 = AluDivQ[85];
  assign x61514 = AluDivQ[86];
  assign x61515 = AluDivQ[87];
  assign x61516 = AluDivQ[88];
  assign x61517 = AluDivQ[89];
  assign x61518 = AluDivQ[90];
  assign x61519 = AluDivQ[91];
  assign x61520 = AluDivQ[92];
  assign x61521 = AluDivQ[93];
  assign x61522 = AluDivQ[94];
  assign x61523 = AluDivQ[95];
  assign x61524 = AluDivQ[96];
  assign x61525 = AluDivQ[97];
  assign x61526 = AluDivQ[98];
  assign x61527 = AluDivQ[99];
  assign x61528 = AluDivQ[100];
  assign x61529 = AluDivQ[101];
  assign x61530 = AluDivQ[102];
  assign x61531 = AluDivQ[103];
  assign x61532 = AluDivQ[104];
  assign x61533 = AluDivQ[105];
  assign x61534 = AluDivQ[106];
  assign x61535 = AluDivQ[107];
  assign x61536 = AluDivQ[108];
  assign x61537 = AluDivQ[109];
  assign x61538 = AluDivQ[110];
  assign x61539 = AluDivQ[111];
  assign x61540 = AluDivQ[112];
  assign x61541 = AluDivQ[113];
  assign x61542 = AluDivQ[114];
  assign x61543 = AluDivQ[115];
  assign x61544 = AluDivQ[116];
  assign x61545 = AluDivQ[117];
  assign x61546 = AluDivQ[118];
  assign x61547 = AluDivQ[119];
  assign x61548 = AluDivQ[120];
  assign x61549 = AluDivQ[121];
  assign x61550 = AluDivQ[122];
  assign x61551 = AluDivQ[123];
  assign x61552 = AluDivQ[124];
  assign x61553 = AluDivQ[125];
  assign x61554 = AluDivQ[126];
  assign x61555 = AluDivQ[127];
  assign x61556 = AluDivR[0];
  assign x61557 = AluDivR[1];
  assign x61558 = AluDivR[2];
  assign x61559 = AluDivR[3];
  assign x61560 = AluDivR[4];
  assign x61561 = AluDivR[5];
  assign x61562 = AluDivR[6];
  assign x61563 = AluDivR[7];
  assign x61564 = AluDivR[8];
  assign x61565 = AluDivR[9];
  assign x61566 = AluDivR[10];
  assign x61567 = AluDivR[11];
  assign x61568 = AluDivR[12];
  assign x61569 = AluDivR[13];
  assign x61570 = AluDivR[14];
  assign x61571 = AluDivR[15];
  assign x61572 = AluDivR[16];
  assign x61573 = AluDivR[17];
  assign x61574 = AluDivR[18];
  assign x61575 = AluDivR[19];
  assign x61576 = AluDivR[20];
  assign x61577 = AluDivR[21];
  assign x61578 = AluDivR[22];
  assign x61579 = AluDivR[23];
  assign x61580 = AluDivR[24];
  assign x61581 = AluDivR[25];
  assign x61582 = AluDivR[26];
  assign x61583 = AluDivR[27];
  assign x61584 = AluDivR[28];
  assign x61585 = AluDivR[29];
  assign x61586 = AluDivR[30];
  assign x61587 = AluDivR[31];
  assign x61588 = AluDivR[32];
  assign x61589 = AluDivR[33];
  assign x61590 = AluDivR[34];
  assign x61591 = AluDivR[35];
  assign x61592 = AluDivR[36];
  assign x61593 = AluDivR[37];
  assign x61594 = AluDivR[38];
  assign x61595 = AluDivR[39];
  assign x61596 = AluDivR[40];
  assign x61597 = AluDivR[41];
  assign x61598 = AluDivR[42];
  assign x61599 = AluDivR[43];
  assign x61600 = AluDivR[44];
  assign x61601 = AluDivR[45];
  assign x61602 = AluDivR[46];
  assign x61603 = AluDivR[47];
  assign x61604 = AluDivR[48];
  assign x61605 = AluDivR[49];
  assign x61606 = AluDivR[50];
  assign x61607 = AluDivR[51];
  assign x61608 = AluDivR[52];
  assign x61609 = AluDivR[53];
  assign x61610 = AluDivR[54];
  assign x61611 = AluDivR[55];
  assign x61612 = AluDivR[56];
  assign x61613 = AluDivR[57];
  assign x61614 = AluDivR[58];
  assign x61615 = AluDivR[59];
  assign x61616 = AluDivR[60];
  assign x61617 = AluDivR[61];
  assign x61618 = AluDivR[62];
  assign x61619 = AluDivR[63];
  assign x61620 = AluDivR[64];
  assign x61621 = AluDivR[65];
  assign x61622 = AluDivR[66];
  assign x61623 = AluDivR[67];
  assign x61624 = AluDivR[68];
  assign x61625 = AluDivR[69];
  assign x61626 = AluDivR[70];
  assign x61627 = AluDivR[71];
  assign x61628 = AluDivR[72];
  assign x61629 = AluDivR[73];
  assign x61630 = AluDivR[74];
  assign x61631 = AluDivR[75];
  assign x61632 = AluDivR[76];
  assign x61633 = AluDivR[77];
  assign x61634 = AluDivR[78];
  assign x61635 = AluDivR[79];
  assign x61636 = AluDivR[80];
  assign x61637 = AluDivR[81];
  assign x61638 = AluDivR[82];
  assign x61639 = AluDivR[83];
  assign x61640 = AluDivR[84];
  assign x61641 = AluDivR[85];
  assign x61642 = AluDivR[86];
  assign x61643 = AluDivR[87];
  assign x61644 = AluDivR[88];
  assign x61645 = AluDivR[89];
  assign x61646 = AluDivR[90];
  assign x61647 = AluDivR[91];
  assign x61648 = AluDivR[92];
  assign x61649 = AluDivR[93];
  assign x61650 = AluDivR[94];
  assign x61651 = AluDivR[95];
  assign x61652 = AluDivR[96];
  assign x61653 = AluDivR[97];
  assign x61654 = AluDivR[98];
  assign x61655 = AluDivR[99];
  assign x61656 = AluDivR[100];
  assign x61657 = AluDivR[101];
  assign x61658 = AluDivR[102];
  assign x61659 = AluDivR[103];
  assign x61660 = AluDivR[104];
  assign x61661 = AluDivR[105];
  assign x61662 = AluDivR[106];
  assign x61663 = AluDivR[107];
  assign x61664 = AluDivR[108];
  assign x61665 = AluDivR[109];
  assign x61666 = AluDivR[110];
  assign x61667 = AluDivR[111];
  assign x61668 = AluDivR[112];
  assign x61669 = AluDivR[113];
  assign x61670 = AluDivR[114];
  assign x61671 = AluDivR[115];
  assign x61672 = AluDivR[116];
  assign x61673 = AluDivR[117];
  assign x61674 = AluDivR[118];
  assign x61675 = AluDivR[119];
  assign x61676 = AluDivR[120];
  assign x61677 = AluDivR[121];
  assign x61678 = AluDivR[122];
  assign x61679 = AluDivR[123];
  assign x61680 = AluDivR[124];
  assign x61681 = AluDivR[125];
  assign x61682 = AluDivR[126];
  assign x61683 = AluDivR[127];
  assign x66601 = FpuBasicFinish;
  assign x66473 = FpuBasicRes[0];
  assign x66474 = FpuBasicRes[1];
  assign x66475 = FpuBasicRes[2];
  assign x66476 = FpuBasicRes[3];
  assign x66477 = FpuBasicRes[4];
  assign x66478 = FpuBasicRes[5];
  assign x66479 = FpuBasicRes[6];
  assign x66480 = FpuBasicRes[7];
  assign x66481 = FpuBasicRes[8];
  assign x66482 = FpuBasicRes[9];
  assign x66483 = FpuBasicRes[10];
  assign x66484 = FpuBasicRes[11];
  assign x66485 = FpuBasicRes[12];
  assign x66486 = FpuBasicRes[13];
  assign x66487 = FpuBasicRes[14];
  assign x66488 = FpuBasicRes[15];
  assign x66489 = FpuBasicRes[16];
  assign x66490 = FpuBasicRes[17];
  assign x66491 = FpuBasicRes[18];
  assign x66492 = FpuBasicRes[19];
  assign x66493 = FpuBasicRes[20];
  assign x66494 = FpuBasicRes[21];
  assign x66495 = FpuBasicRes[22];
  assign x66496 = FpuBasicRes[23];
  assign x66497 = FpuBasicRes[24];
  assign x66498 = FpuBasicRes[25];
  assign x66499 = FpuBasicRes[26];
  assign x66500 = FpuBasicRes[27];
  assign x66501 = FpuBasicRes[28];
  assign x66502 = FpuBasicRes[29];
  assign x66503 = FpuBasicRes[30];
  assign x66504 = FpuBasicRes[31];
  assign x66505 = FpuBasicRes[32];
  assign x66506 = FpuBasicRes[33];
  assign x66507 = FpuBasicRes[34];
  assign x66508 = FpuBasicRes[35];
  assign x66509 = FpuBasicRes[36];
  assign x66510 = FpuBasicRes[37];
  assign x66511 = FpuBasicRes[38];
  assign x66512 = FpuBasicRes[39];
  assign x66513 = FpuBasicRes[40];
  assign x66514 = FpuBasicRes[41];
  assign x66515 = FpuBasicRes[42];
  assign x66516 = FpuBasicRes[43];
  assign x66517 = FpuBasicRes[44];
  assign x66518 = FpuBasicRes[45];
  assign x66519 = FpuBasicRes[46];
  assign x66520 = FpuBasicRes[47];
  assign x66521 = FpuBasicRes[48];
  assign x66522 = FpuBasicRes[49];
  assign x66523 = FpuBasicRes[50];
  assign x66524 = FpuBasicRes[51];
  assign x66525 = FpuBasicRes[52];
  assign x66526 = FpuBasicRes[53];
  assign x66527 = FpuBasicRes[54];
  assign x66528 = FpuBasicRes[55];
  assign x66529 = FpuBasicRes[56];
  assign x66530 = FpuBasicRes[57];
  assign x66531 = FpuBasicRes[58];
  assign x66532 = FpuBasicRes[59];
  assign x66533 = FpuBasicRes[60];
  assign x66534 = FpuBasicRes[61];
  assign x66535 = FpuBasicRes[62];
  assign x66536 = FpuBasicRes[63];
  assign x66537 = FpuBasicRes[64];
  assign x66538 = FpuBasicRes[65];
  assign x66539 = FpuBasicRes[66];
  assign x66540 = FpuBasicRes[67];
  assign x66541 = FpuBasicRes[68];
  assign x66542 = FpuBasicRes[69];
  assign x66543 = FpuBasicRes[70];
  assign x66544 = FpuBasicRes[71];
  assign x66545 = FpuBasicRes[72];
  assign x66546 = FpuBasicRes[73];
  assign x66547 = FpuBasicRes[74];
  assign x66548 = FpuBasicRes[75];
  assign x66549 = FpuBasicRes[76];
  assign x66550 = FpuBasicRes[77];
  assign x66551 = FpuBasicRes[78];
  assign x66552 = FpuBasicRes[79];
  assign x66553 = FpuBasicRes[80];
  assign x66554 = FpuBasicRes[81];
  assign x66555 = FpuBasicRes[82];
  assign x66556 = FpuBasicRes[83];
  assign x66557 = FpuBasicRes[84];
  assign x66558 = FpuBasicRes[85];
  assign x66559 = FpuBasicRes[86];
  assign x66560 = FpuBasicRes[87];
  assign x66561 = FpuBasicRes[88];
  assign x66562 = FpuBasicRes[89];
  assign x66563 = FpuBasicRes[90];
  assign x66564 = FpuBasicRes[91];
  assign x66565 = FpuBasicRes[92];
  assign x66566 = FpuBasicRes[93];
  assign x66567 = FpuBasicRes[94];
  assign x66568 = FpuBasicRes[95];
  assign x66569 = FpuBasicRes[96];
  assign x66570 = FpuBasicRes[97];
  assign x66571 = FpuBasicRes[98];
  assign x66572 = FpuBasicRes[99];
  assign x66573 = FpuBasicRes[100];
  assign x66574 = FpuBasicRes[101];
  assign x66575 = FpuBasicRes[102];
  assign x66576 = FpuBasicRes[103];
  assign x66577 = FpuBasicRes[104];
  assign x66578 = FpuBasicRes[105];
  assign x66579 = FpuBasicRes[106];
  assign x66580 = FpuBasicRes[107];
  assign x66581 = FpuBasicRes[108];
  assign x66582 = FpuBasicRes[109];
  assign x66583 = FpuBasicRes[110];
  assign x66584 = FpuBasicRes[111];
  assign x66585 = FpuBasicRes[112];
  assign x66586 = FpuBasicRes[113];
  assign x66587 = FpuBasicRes[114];
  assign x66588 = FpuBasicRes[115];
  assign x66589 = FpuBasicRes[116];
  assign x66590 = FpuBasicRes[117];
  assign x66591 = FpuBasicRes[118];
  assign x66592 = FpuBasicRes[119];
  assign x66593 = FpuBasicRes[120];
  assign x66594 = FpuBasicRes[121];
  assign x66595 = FpuBasicRes[122];
  assign x66596 = FpuBasicRes[123];
  assign x66597 = FpuBasicRes[124];
  assign x66598 = FpuBasicRes[125];
  assign x66599 = FpuBasicRes[126];
  assign x66600 = FpuBasicRes[127];
  assign x67594 = FpuMultFinish;
  assign x67466 = FpuMultRes[0];
  assign x67467 = FpuMultRes[1];
  assign x67468 = FpuMultRes[2];
  assign x67469 = FpuMultRes[3];
  assign x67470 = FpuMultRes[4];
  assign x67471 = FpuMultRes[5];
  assign x67472 = FpuMultRes[6];
  assign x67473 = FpuMultRes[7];
  assign x67474 = FpuMultRes[8];
  assign x67475 = FpuMultRes[9];
  assign x67476 = FpuMultRes[10];
  assign x67477 = FpuMultRes[11];
  assign x67478 = FpuMultRes[12];
  assign x67479 = FpuMultRes[13];
  assign x67480 = FpuMultRes[14];
  assign x67481 = FpuMultRes[15];
  assign x67482 = FpuMultRes[16];
  assign x67483 = FpuMultRes[17];
  assign x67484 = FpuMultRes[18];
  assign x67485 = FpuMultRes[19];
  assign x67486 = FpuMultRes[20];
  assign x67487 = FpuMultRes[21];
  assign x67488 = FpuMultRes[22];
  assign x67489 = FpuMultRes[23];
  assign x67490 = FpuMultRes[24];
  assign x67491 = FpuMultRes[25];
  assign x67492 = FpuMultRes[26];
  assign x67493 = FpuMultRes[27];
  assign x67494 = FpuMultRes[28];
  assign x67495 = FpuMultRes[29];
  assign x67496 = FpuMultRes[30];
  assign x67497 = FpuMultRes[31];
  assign x67498 = FpuMultRes[32];
  assign x67499 = FpuMultRes[33];
  assign x67500 = FpuMultRes[34];
  assign x67501 = FpuMultRes[35];
  assign x67502 = FpuMultRes[36];
  assign x67503 = FpuMultRes[37];
  assign x67504 = FpuMultRes[38];
  assign x67505 = FpuMultRes[39];
  assign x67506 = FpuMultRes[40];
  assign x67507 = FpuMultRes[41];
  assign x67508 = FpuMultRes[42];
  assign x67509 = FpuMultRes[43];
  assign x67510 = FpuMultRes[44];
  assign x67511 = FpuMultRes[45];
  assign x67512 = FpuMultRes[46];
  assign x67513 = FpuMultRes[47];
  assign x67514 = FpuMultRes[48];
  assign x67515 = FpuMultRes[49];
  assign x67516 = FpuMultRes[50];
  assign x67517 = FpuMultRes[51];
  assign x67518 = FpuMultRes[52];
  assign x67519 = FpuMultRes[53];
  assign x67520 = FpuMultRes[54];
  assign x67521 = FpuMultRes[55];
  assign x67522 = FpuMultRes[56];
  assign x67523 = FpuMultRes[57];
  assign x67524 = FpuMultRes[58];
  assign x67525 = FpuMultRes[59];
  assign x67526 = FpuMultRes[60];
  assign x67527 = FpuMultRes[61];
  assign x67528 = FpuMultRes[62];
  assign x67529 = FpuMultRes[63];
  assign x67530 = FpuMultRes[64];
  assign x67531 = FpuMultRes[65];
  assign x67532 = FpuMultRes[66];
  assign x67533 = FpuMultRes[67];
  assign x67534 = FpuMultRes[68];
  assign x67535 = FpuMultRes[69];
  assign x67536 = FpuMultRes[70];
  assign x67537 = FpuMultRes[71];
  assign x67538 = FpuMultRes[72];
  assign x67539 = FpuMultRes[73];
  assign x67540 = FpuMultRes[74];
  assign x67541 = FpuMultRes[75];
  assign x67542 = FpuMultRes[76];
  assign x67543 = FpuMultRes[77];
  assign x67544 = FpuMultRes[78];
  assign x67545 = FpuMultRes[79];
  assign x67546 = FpuMultRes[80];
  assign x67547 = FpuMultRes[81];
  assign x67548 = FpuMultRes[82];
  assign x67549 = FpuMultRes[83];
  assign x67550 = FpuMultRes[84];
  assign x67551 = FpuMultRes[85];
  assign x67552 = FpuMultRes[86];
  assign x67553 = FpuMultRes[87];
  assign x67554 = FpuMultRes[88];
  assign x67555 = FpuMultRes[89];
  assign x67556 = FpuMultRes[90];
  assign x67557 = FpuMultRes[91];
  assign x67558 = FpuMultRes[92];
  assign x67559 = FpuMultRes[93];
  assign x67560 = FpuMultRes[94];
  assign x67561 = FpuMultRes[95];
  assign x67562 = FpuMultRes[96];
  assign x67563 = FpuMultRes[97];
  assign x67564 = FpuMultRes[98];
  assign x67565 = FpuMultRes[99];
  assign x67566 = FpuMultRes[100];
  assign x67567 = FpuMultRes[101];
  assign x67568 = FpuMultRes[102];
  assign x67569 = FpuMultRes[103];
  assign x67570 = FpuMultRes[104];
  assign x67571 = FpuMultRes[105];
  assign x67572 = FpuMultRes[106];
  assign x67573 = FpuMultRes[107];
  assign x67574 = FpuMultRes[108];
  assign x67575 = FpuMultRes[109];
  assign x67576 = FpuMultRes[110];
  assign x67577 = FpuMultRes[111];
  assign x67578 = FpuMultRes[112];
  assign x67579 = FpuMultRes[113];
  assign x67580 = FpuMultRes[114];
  assign x67581 = FpuMultRes[115];
  assign x67582 = FpuMultRes[116];
  assign x67583 = FpuMultRes[117];
  assign x67584 = FpuMultRes[118];
  assign x67585 = FpuMultRes[119];
  assign x67586 = FpuMultRes[120];
  assign x67587 = FpuMultRes[121];
  assign x67588 = FpuMultRes[122];
  assign x67589 = FpuMultRes[123];
  assign x67590 = FpuMultRes[124];
  assign x67591 = FpuMultRes[125];
  assign x67592 = FpuMultRes[126];
  assign x67593 = FpuMultRes[127];

  assign AluDivA[0] = x75499;
  assign AluDivA[1] = x75502;
  assign AluDivA[2] = x75505;
  assign AluDivA[3] = x75508;
  assign AluDivA[4] = x75511;
  assign AluDivA[5] = x75514;
  assign AluDivA[6] = x75517;
  assign AluDivA[7] = x75520;
  assign AluDivA[8] = x75523;
  assign AluDivA[9] = x75526;
  assign AluDivA[10] = x75529;
  assign AluDivA[11] = x75532;
  assign AluDivA[12] = x75535;
  assign AluDivA[13] = x75538;
  assign AluDivA[14] = x75541;
  assign AluDivA[15] = x75544;
  assign AluDivA[16] = x75547;
  assign AluDivA[17] = x75550;
  assign AluDivA[18] = x75553;
  assign AluDivA[19] = x75556;
  assign AluDivA[20] = x75559;
  assign AluDivA[21] = x75562;
  assign AluDivA[22] = x75565;
  assign AluDivA[23] = x75568;
  assign AluDivA[24] = x75571;
  assign AluDivA[25] = x75574;
  assign AluDivA[26] = x75577;
  assign AluDivA[27] = x75580;
  assign AluDivA[28] = x75583;
  assign AluDivA[29] = x75586;
  assign AluDivA[30] = x75589;
  assign AluDivA[31] = x75592;
  assign AluDivA[32] = x75793;
  assign AluDivA[33] = x75796;
  assign AluDivA[34] = x75799;
  assign AluDivA[35] = x75802;
  assign AluDivA[36] = x75805;
  assign AluDivA[37] = x75808;
  assign AluDivA[38] = x75811;
  assign AluDivA[39] = x75814;
  assign AluDivA[40] = x75817;
  assign AluDivA[41] = x75820;
  assign AluDivA[42] = x75823;
  assign AluDivA[43] = x75826;
  assign AluDivA[44] = x75829;
  assign AluDivA[45] = x75832;
  assign AluDivA[46] = x75835;
  assign AluDivA[47] = x75838;
  assign AluDivA[48] = x75841;
  assign AluDivA[49] = x75844;
  assign AluDivA[50] = x75847;
  assign AluDivA[51] = x75850;
  assign AluDivA[52] = x75853;
  assign AluDivA[53] = x75856;
  assign AluDivA[54] = x75859;
  assign AluDivA[55] = x75862;
  assign AluDivA[56] = x75865;
  assign AluDivA[57] = x75868;
  assign AluDivA[58] = x75871;
  assign AluDivA[59] = x75874;
  assign AluDivA[60] = x75877;
  assign AluDivA[61] = x75880;
  assign AluDivA[62] = x75883;
  assign AluDivA[63] = x75886;
  assign AluDivA[64] = x76087;
  assign AluDivA[65] = x76090;
  assign AluDivA[66] = x76093;
  assign AluDivA[67] = x76096;
  assign AluDivA[68] = x76099;
  assign AluDivA[69] = x76102;
  assign AluDivA[70] = x76105;
  assign AluDivA[71] = x76108;
  assign AluDivA[72] = x76111;
  assign AluDivA[73] = x76114;
  assign AluDivA[74] = x76117;
  assign AluDivA[75] = x76120;
  assign AluDivA[76] = x76123;
  assign AluDivA[77] = x76126;
  assign AluDivA[78] = x76129;
  assign AluDivA[79] = x76132;
  assign AluDivA[80] = x76135;
  assign AluDivA[81] = x76138;
  assign AluDivA[82] = x76141;
  assign AluDivA[83] = x76144;
  assign AluDivA[84] = x76147;
  assign AluDivA[85] = x76150;
  assign AluDivA[86] = x76153;
  assign AluDivA[87] = x76156;
  assign AluDivA[88] = x76159;
  assign AluDivA[89] = x76162;
  assign AluDivA[90] = x76165;
  assign AluDivA[91] = x76168;
  assign AluDivA[92] = x76171;
  assign AluDivA[93] = x76174;
  assign AluDivA[94] = x76177;
  assign AluDivA[95] = x76180;
  assign AluDivA[96] = x76381;
  assign AluDivA[97] = x76384;
  assign AluDivA[98] = x76387;
  assign AluDivA[99] = x76390;
  assign AluDivA[100] = x76393;
  assign AluDivA[101] = x76396;
  assign AluDivA[102] = x76399;
  assign AluDivA[103] = x76402;
  assign AluDivA[104] = x76405;
  assign AluDivA[105] = x76408;
  assign AluDivA[106] = x76411;
  assign AluDivA[107] = x76414;
  assign AluDivA[108] = x76417;
  assign AluDivA[109] = x76420;
  assign AluDivA[110] = x76423;
  assign AluDivA[111] = x76426;
  assign AluDivA[112] = x76429;
  assign AluDivA[113] = x76432;
  assign AluDivA[114] = x76435;
  assign AluDivA[115] = x76438;
  assign AluDivA[116] = x76441;
  assign AluDivA[117] = x76444;
  assign AluDivA[118] = x76447;
  assign AluDivA[119] = x76450;
  assign AluDivA[120] = x76453;
  assign AluDivA[121] = x76456;
  assign AluDivA[122] = x76459;
  assign AluDivA[123] = x76462;
  assign AluDivA[124] = x76465;
  assign AluDivA[125] = x76468;
  assign AluDivA[126] = x76471;
  assign AluDivA[127] = x76474;
  assign AluDivB[0] = x61688;
  assign AluDivB[1] = x61691;
  assign AluDivB[2] = x61694;
  assign AluDivB[3] = x61697;
  assign AluDivB[4] = x61700;
  assign AluDivB[5] = x61703;
  assign AluDivB[6] = x61706;
  assign AluDivB[7] = x61709;
  assign AluDivB[8] = x61712;
  assign AluDivB[9] = x61715;
  assign AluDivB[10] = x61718;
  assign AluDivB[11] = x61721;
  assign AluDivB[12] = x61724;
  assign AluDivB[13] = x61727;
  assign AluDivB[14] = x61730;
  assign AluDivB[15] = x61733;
  assign AluDivB[16] = x61736;
  assign AluDivB[17] = x61739;
  assign AluDivB[18] = x61742;
  assign AluDivB[19] = x61745;
  assign AluDivB[20] = x61748;
  assign AluDivB[21] = x61751;
  assign AluDivB[22] = x61754;
  assign AluDivB[23] = x61757;
  assign AluDivB[24] = x61760;
  assign AluDivB[25] = x61763;
  assign AluDivB[26] = x61766;
  assign AluDivB[27] = x61769;
  assign AluDivB[28] = x61772;
  assign AluDivB[29] = x61775;
  assign AluDivB[30] = x61778;
  assign AluDivB[31] = x61781;
  assign AluDivB[32] = x61783;
  assign AluDivB[33] = x61785;
  assign AluDivB[34] = x61787;
  assign AluDivB[35] = x61789;
  assign AluDivB[36] = x61791;
  assign AluDivB[37] = x61793;
  assign AluDivB[38] = x61795;
  assign AluDivB[39] = x61797;
  assign AluDivB[40] = x61799;
  assign AluDivB[41] = x61801;
  assign AluDivB[42] = x61803;
  assign AluDivB[43] = x61805;
  assign AluDivB[44] = x61807;
  assign AluDivB[45] = x61809;
  assign AluDivB[46] = x61811;
  assign AluDivB[47] = x61813;
  assign AluDivB[48] = x61815;
  assign AluDivB[49] = x61817;
  assign AluDivB[50] = x61819;
  assign AluDivB[51] = x61821;
  assign AluDivB[52] = x61823;
  assign AluDivB[53] = x61825;
  assign AluDivB[54] = x61827;
  assign AluDivB[55] = x61829;
  assign AluDivB[56] = x61831;
  assign AluDivB[57] = x61833;
  assign AluDivB[58] = x61835;
  assign AluDivB[59] = x61837;
  assign AluDivB[60] = x61839;
  assign AluDivB[61] = x61841;
  assign AluDivB[62] = x61843;
  assign AluDivB[63] = x61845;
  assign AluDivB[64] = x61847;
  assign AluDivB[65] = x61849;
  assign AluDivB[66] = x61851;
  assign AluDivB[67] = x61853;
  assign AluDivB[68] = x61855;
  assign AluDivB[69] = x61857;
  assign AluDivB[70] = x61859;
  assign AluDivB[71] = x61861;
  assign AluDivB[72] = x61863;
  assign AluDivB[73] = x61865;
  assign AluDivB[74] = x61867;
  assign AluDivB[75] = x61869;
  assign AluDivB[76] = x61871;
  assign AluDivB[77] = x61873;
  assign AluDivB[78] = x61875;
  assign AluDivB[79] = x61877;
  assign AluDivB[80] = x61879;
  assign AluDivB[81] = x61881;
  assign AluDivB[82] = x61883;
  assign AluDivB[83] = x61885;
  assign AluDivB[84] = x61887;
  assign AluDivB[85] = x61889;
  assign AluDivB[86] = x61891;
  assign AluDivB[87] = x61893;
  assign AluDivB[88] = x61895;
  assign AluDivB[89] = x61897;
  assign AluDivB[90] = x61899;
  assign AluDivB[91] = x61901;
  assign AluDivB[92] = x61903;
  assign AluDivB[93] = x61905;
  assign AluDivB[94] = x61907;
  assign AluDivB[95] = x61909;
  assign AluDivB[96] = x61911;
  assign AluDivB[97] = x61913;
  assign AluDivB[98] = x61915;
  assign AluDivB[99] = x61917;
  assign AluDivB[100] = x61919;
  assign AluDivB[101] = x61921;
  assign AluDivB[102] = x61923;
  assign AluDivB[103] = x61925;
  assign AluDivB[104] = x61927;
  assign AluDivB[105] = x61929;
  assign AluDivB[106] = x61931;
  assign AluDivB[107] = x61933;
  assign AluDivB[108] = x61935;
  assign AluDivB[109] = x61937;
  assign AluDivB[110] = x61939;
  assign AluDivB[111] = x61941;
  assign AluDivB[112] = x61943;
  assign AluDivB[113] = x61945;
  assign AluDivB[114] = x61947;
  assign AluDivB[115] = x61949;
  assign AluDivB[116] = x61951;
  assign AluDivB[117] = x61953;
  assign AluDivB[118] = x61955;
  assign AluDivB[119] = x61957;
  assign AluDivB[120] = x61959;
  assign AluDivB[121] = x61961;
  assign AluDivB[122] = x61963;
  assign AluDivB[123] = x61965;
  assign AluDivB[124] = x61967;
  assign AluDivB[125] = x61969;
  assign AluDivB[126] = x61971;
  assign AluDivB[127] = x61973;
  assign AluDivStall = x68740;
  assign AluDivValid = x83362;
  assign FpuBasicA[0] = x78169;
  assign FpuBasicA[1] = x78172;
  assign FpuBasicA[2] = x78175;
  assign FpuBasicA[3] = x78178;
  assign FpuBasicA[4] = x78181;
  assign FpuBasicA[5] = x78184;
  assign FpuBasicA[6] = x78187;
  assign FpuBasicA[7] = x78190;
  assign FpuBasicA[8] = x78193;
  assign FpuBasicA[9] = x78196;
  assign FpuBasicA[10] = x78199;
  assign FpuBasicA[11] = x78202;
  assign FpuBasicA[12] = x78205;
  assign FpuBasicA[13] = x78208;
  assign FpuBasicA[14] = x78211;
  assign FpuBasicA[15] = x78214;
  assign FpuBasicA[16] = x78217;
  assign FpuBasicA[17] = x78220;
  assign FpuBasicA[18] = x78223;
  assign FpuBasicA[19] = x78226;
  assign FpuBasicA[20] = x78229;
  assign FpuBasicA[21] = x78232;
  assign FpuBasicA[22] = x78235;
  assign FpuBasicA[23] = x78238;
  assign FpuBasicA[24] = x78241;
  assign FpuBasicA[25] = x78244;
  assign FpuBasicA[26] = x78247;
  assign FpuBasicA[27] = x78250;
  assign FpuBasicA[28] = x78253;
  assign FpuBasicA[29] = x78256;
  assign FpuBasicA[30] = x78259;
  assign FpuBasicA[31] = x78262;
  assign FpuBasicA[32] = x78463;
  assign FpuBasicA[33] = x78466;
  assign FpuBasicA[34] = x78469;
  assign FpuBasicA[35] = x78472;
  assign FpuBasicA[36] = x78475;
  assign FpuBasicA[37] = x78478;
  assign FpuBasicA[38] = x78481;
  assign FpuBasicA[39] = x78484;
  assign FpuBasicA[40] = x78487;
  assign FpuBasicA[41] = x78490;
  assign FpuBasicA[42] = x78493;
  assign FpuBasicA[43] = x78496;
  assign FpuBasicA[44] = x78499;
  assign FpuBasicA[45] = x78502;
  assign FpuBasicA[46] = x78505;
  assign FpuBasicA[47] = x78508;
  assign FpuBasicA[48] = x78511;
  assign FpuBasicA[49] = x78514;
  assign FpuBasicA[50] = x78517;
  assign FpuBasicA[51] = x78520;
  assign FpuBasicA[52] = x78523;
  assign FpuBasicA[53] = x78526;
  assign FpuBasicA[54] = x78529;
  assign FpuBasicA[55] = x78532;
  assign FpuBasicA[56] = x78535;
  assign FpuBasicA[57] = x78538;
  assign FpuBasicA[58] = x78541;
  assign FpuBasicA[59] = x78544;
  assign FpuBasicA[60] = x78547;
  assign FpuBasicA[61] = x78550;
  assign FpuBasicA[62] = x78553;
  assign FpuBasicA[63] = x78556;
  assign FpuBasicA[64] = x78757;
  assign FpuBasicA[65] = x78760;
  assign FpuBasicA[66] = x78763;
  assign FpuBasicA[67] = x78766;
  assign FpuBasicA[68] = x78769;
  assign FpuBasicA[69] = x78772;
  assign FpuBasicA[70] = x78775;
  assign FpuBasicA[71] = x78778;
  assign FpuBasicA[72] = x78781;
  assign FpuBasicA[73] = x78784;
  assign FpuBasicA[74] = x78787;
  assign FpuBasicA[75] = x78790;
  assign FpuBasicA[76] = x78793;
  assign FpuBasicA[77] = x78796;
  assign FpuBasicA[78] = x78799;
  assign FpuBasicA[79] = x78802;
  assign FpuBasicA[80] = x78805;
  assign FpuBasicA[81] = x78808;
  assign FpuBasicA[82] = x78811;
  assign FpuBasicA[83] = x78814;
  assign FpuBasicA[84] = x78817;
  assign FpuBasicA[85] = x78820;
  assign FpuBasicA[86] = x78823;
  assign FpuBasicA[87] = x78826;
  assign FpuBasicA[88] = x78829;
  assign FpuBasicA[89] = x78832;
  assign FpuBasicA[90] = x78835;
  assign FpuBasicA[91] = x78838;
  assign FpuBasicA[92] = x78841;
  assign FpuBasicA[93] = x78844;
  assign FpuBasicA[94] = x78847;
  assign FpuBasicA[95] = x78850;
  assign FpuBasicA[96] = x79051;
  assign FpuBasicA[97] = x79054;
  assign FpuBasicA[98] = x79057;
  assign FpuBasicA[99] = x79060;
  assign FpuBasicA[100] = x79063;
  assign FpuBasicA[101] = x79066;
  assign FpuBasicA[102] = x79069;
  assign FpuBasicA[103] = x79072;
  assign FpuBasicA[104] = x79075;
  assign FpuBasicA[105] = x79078;
  assign FpuBasicA[106] = x79081;
  assign FpuBasicA[107] = x79084;
  assign FpuBasicA[108] = x79087;
  assign FpuBasicA[109] = x79090;
  assign FpuBasicA[110] = x79093;
  assign FpuBasicA[111] = x79096;
  assign FpuBasicA[112] = x79099;
  assign FpuBasicA[113] = x79102;
  assign FpuBasicA[114] = x79105;
  assign FpuBasicA[115] = x79108;
  assign FpuBasicA[116] = x79111;
  assign FpuBasicA[117] = x79114;
  assign FpuBasicA[118] = x79117;
  assign FpuBasicA[119] = x79120;
  assign FpuBasicA[120] = x79123;
  assign FpuBasicA[121] = x79126;
  assign FpuBasicA[122] = x79129;
  assign FpuBasicA[123] = x79132;
  assign FpuBasicA[124] = x79135;
  assign FpuBasicA[125] = x79138;
  assign FpuBasicA[126] = x79141;
  assign FpuBasicA[127] = x79144;
  assign FpuBasicB[0] = x66605;
  assign FpuBasicB[1] = x66608;
  assign FpuBasicB[2] = x66611;
  assign FpuBasicB[3] = x66614;
  assign FpuBasicB[4] = x66617;
  assign FpuBasicB[5] = x66620;
  assign FpuBasicB[6] = x66623;
  assign FpuBasicB[7] = x66626;
  assign FpuBasicB[8] = x66629;
  assign FpuBasicB[9] = x66632;
  assign FpuBasicB[10] = x66635;
  assign FpuBasicB[11] = x66638;
  assign FpuBasicB[12] = x66641;
  assign FpuBasicB[13] = x66644;
  assign FpuBasicB[14] = x66647;
  assign FpuBasicB[15] = x66650;
  assign FpuBasicB[16] = x66653;
  assign FpuBasicB[17] = x66656;
  assign FpuBasicB[18] = x66659;
  assign FpuBasicB[19] = x66662;
  assign FpuBasicB[20] = x66665;
  assign FpuBasicB[21] = x66668;
  assign FpuBasicB[22] = x66671;
  assign FpuBasicB[23] = x66674;
  assign FpuBasicB[24] = x66677;
  assign FpuBasicB[25] = x66680;
  assign FpuBasicB[26] = x66683;
  assign FpuBasicB[27] = x66686;
  assign FpuBasicB[28] = x66689;
  assign FpuBasicB[29] = x66692;
  assign FpuBasicB[30] = x66695;
  assign FpuBasicB[31] = x66698;
  assign FpuBasicB[32] = x66700;
  assign FpuBasicB[33] = x66702;
  assign FpuBasicB[34] = x66704;
  assign FpuBasicB[35] = x66706;
  assign FpuBasicB[36] = x66708;
  assign FpuBasicB[37] = x66710;
  assign FpuBasicB[38] = x66712;
  assign FpuBasicB[39] = x66714;
  assign FpuBasicB[40] = x66716;
  assign FpuBasicB[41] = x66718;
  assign FpuBasicB[42] = x66720;
  assign FpuBasicB[43] = x66722;
  assign FpuBasicB[44] = x66724;
  assign FpuBasicB[45] = x66726;
  assign FpuBasicB[46] = x66728;
  assign FpuBasicB[47] = x66730;
  assign FpuBasicB[48] = x66732;
  assign FpuBasicB[49] = x66734;
  assign FpuBasicB[50] = x66736;
  assign FpuBasicB[51] = x66738;
  assign FpuBasicB[52] = x66740;
  assign FpuBasicB[53] = x66742;
  assign FpuBasicB[54] = x66744;
  assign FpuBasicB[55] = x66746;
  assign FpuBasicB[56] = x66748;
  assign FpuBasicB[57] = x66750;
  assign FpuBasicB[58] = x66752;
  assign FpuBasicB[59] = x66754;
  assign FpuBasicB[60] = x66756;
  assign FpuBasicB[61] = x66758;
  assign FpuBasicB[62] = x66760;
  assign FpuBasicB[63] = x66762;
  assign FpuBasicB[64] = x66764;
  assign FpuBasicB[65] = x66766;
  assign FpuBasicB[66] = x66768;
  assign FpuBasicB[67] = x66770;
  assign FpuBasicB[68] = x66772;
  assign FpuBasicB[69] = x66774;
  assign FpuBasicB[70] = x66776;
  assign FpuBasicB[71] = x66778;
  assign FpuBasicB[72] = x66780;
  assign FpuBasicB[73] = x66782;
  assign FpuBasicB[74] = x66784;
  assign FpuBasicB[75] = x66786;
  assign FpuBasicB[76] = x66788;
  assign FpuBasicB[77] = x66790;
  assign FpuBasicB[78] = x66792;
  assign FpuBasicB[79] = x66794;
  assign FpuBasicB[80] = x66796;
  assign FpuBasicB[81] = x66798;
  assign FpuBasicB[82] = x66800;
  assign FpuBasicB[83] = x66802;
  assign FpuBasicB[84] = x66804;
  assign FpuBasicB[85] = x66806;
  assign FpuBasicB[86] = x66808;
  assign FpuBasicB[87] = x66810;
  assign FpuBasicB[88] = x66812;
  assign FpuBasicB[89] = x66814;
  assign FpuBasicB[90] = x66816;
  assign FpuBasicB[91] = x66818;
  assign FpuBasicB[92] = x66820;
  assign FpuBasicB[93] = x66822;
  assign FpuBasicB[94] = x66824;
  assign FpuBasicB[95] = x66826;
  assign FpuBasicB[96] = x66828;
  assign FpuBasicB[97] = x66830;
  assign FpuBasicB[98] = x66832;
  assign FpuBasicB[99] = x66834;
  assign FpuBasicB[100] = x66836;
  assign FpuBasicB[101] = x66838;
  assign FpuBasicB[102] = x66840;
  assign FpuBasicB[103] = x66842;
  assign FpuBasicB[104] = x66844;
  assign FpuBasicB[105] = x66846;
  assign FpuBasicB[106] = x66848;
  assign FpuBasicB[107] = x66850;
  assign FpuBasicB[108] = x66852;
  assign FpuBasicB[109] = x66854;
  assign FpuBasicB[110] = x66856;
  assign FpuBasicB[111] = x66858;
  assign FpuBasicB[112] = x66860;
  assign FpuBasicB[113] = x66862;
  assign FpuBasicB[114] = x66864;
  assign FpuBasicB[115] = x66866;
  assign FpuBasicB[116] = x66868;
  assign FpuBasicB[117] = x66870;
  assign FpuBasicB[118] = x66872;
  assign FpuBasicB[119] = x66874;
  assign FpuBasicB[120] = x66876;
  assign FpuBasicB[121] = x66878;
  assign FpuBasicB[122] = x66880;
  assign FpuBasicB[123] = x66882;
  assign FpuBasicB[124] = x66884;
  assign FpuBasicB[125] = x66886;
  assign FpuBasicB[126] = x66888;
  assign FpuBasicB[127] = x66890;
  assign FpuBasicOp[0] = x78127;
  assign FpuBasicOp[1] = x78130;
  assign FpuBasicOp[2] = x78133;
  assign FpuBasicOp[3] = x78136;
  assign FpuBasicOp[4] = x78139;
  assign FpuBasicOp[5] = x78142;
  assign FpuBasicStall = x68742;
  assign FpuBasicValid = x83372;
  assign FpuMultA[0] = x79504;
  assign FpuMultA[1] = x79507;
  assign FpuMultA[2] = x79510;
  assign FpuMultA[3] = x79513;
  assign FpuMultA[4] = x79516;
  assign FpuMultA[5] = x79519;
  assign FpuMultA[6] = x79522;
  assign FpuMultA[7] = x79525;
  assign FpuMultA[8] = x79528;
  assign FpuMultA[9] = x79531;
  assign FpuMultA[10] = x79534;
  assign FpuMultA[11] = x79537;
  assign FpuMultA[12] = x79540;
  assign FpuMultA[13] = x79543;
  assign FpuMultA[14] = x79546;
  assign FpuMultA[15] = x79549;
  assign FpuMultA[16] = x79552;
  assign FpuMultA[17] = x79555;
  assign FpuMultA[18] = x79558;
  assign FpuMultA[19] = x79561;
  assign FpuMultA[20] = x79564;
  assign FpuMultA[21] = x79567;
  assign FpuMultA[22] = x79570;
  assign FpuMultA[23] = x79573;
  assign FpuMultA[24] = x79576;
  assign FpuMultA[25] = x79579;
  assign FpuMultA[26] = x79582;
  assign FpuMultA[27] = x79585;
  assign FpuMultA[28] = x79588;
  assign FpuMultA[29] = x79591;
  assign FpuMultA[30] = x79594;
  assign FpuMultA[31] = x79597;
  assign FpuMultA[32] = x79798;
  assign FpuMultA[33] = x79801;
  assign FpuMultA[34] = x79804;
  assign FpuMultA[35] = x79807;
  assign FpuMultA[36] = x79810;
  assign FpuMultA[37] = x79813;
  assign FpuMultA[38] = x79816;
  assign FpuMultA[39] = x79819;
  assign FpuMultA[40] = x79822;
  assign FpuMultA[41] = x79825;
  assign FpuMultA[42] = x79828;
  assign FpuMultA[43] = x79831;
  assign FpuMultA[44] = x79834;
  assign FpuMultA[45] = x79837;
  assign FpuMultA[46] = x79840;
  assign FpuMultA[47] = x79843;
  assign FpuMultA[48] = x79846;
  assign FpuMultA[49] = x79849;
  assign FpuMultA[50] = x79852;
  assign FpuMultA[51] = x79855;
  assign FpuMultA[52] = x79858;
  assign FpuMultA[53] = x79861;
  assign FpuMultA[54] = x79864;
  assign FpuMultA[55] = x79867;
  assign FpuMultA[56] = x79870;
  assign FpuMultA[57] = x79873;
  assign FpuMultA[58] = x79876;
  assign FpuMultA[59] = x79879;
  assign FpuMultA[60] = x79882;
  assign FpuMultA[61] = x79885;
  assign FpuMultA[62] = x79888;
  assign FpuMultA[63] = x79891;
  assign FpuMultA[64] = x80092;
  assign FpuMultA[65] = x80095;
  assign FpuMultA[66] = x80098;
  assign FpuMultA[67] = x80101;
  assign FpuMultA[68] = x80104;
  assign FpuMultA[69] = x80107;
  assign FpuMultA[70] = x80110;
  assign FpuMultA[71] = x80113;
  assign FpuMultA[72] = x80116;
  assign FpuMultA[73] = x80119;
  assign FpuMultA[74] = x80122;
  assign FpuMultA[75] = x80125;
  assign FpuMultA[76] = x80128;
  assign FpuMultA[77] = x80131;
  assign FpuMultA[78] = x80134;
  assign FpuMultA[79] = x80137;
  assign FpuMultA[80] = x80140;
  assign FpuMultA[81] = x80143;
  assign FpuMultA[82] = x80146;
  assign FpuMultA[83] = x80149;
  assign FpuMultA[84] = x80152;
  assign FpuMultA[85] = x80155;
  assign FpuMultA[86] = x80158;
  assign FpuMultA[87] = x80161;
  assign FpuMultA[88] = x80164;
  assign FpuMultA[89] = x80167;
  assign FpuMultA[90] = x80170;
  assign FpuMultA[91] = x80173;
  assign FpuMultA[92] = x80176;
  assign FpuMultA[93] = x80179;
  assign FpuMultA[94] = x80182;
  assign FpuMultA[95] = x80185;
  assign FpuMultA[96] = x80386;
  assign FpuMultA[97] = x80389;
  assign FpuMultA[98] = x80392;
  assign FpuMultA[99] = x80395;
  assign FpuMultA[100] = x80398;
  assign FpuMultA[101] = x80401;
  assign FpuMultA[102] = x80404;
  assign FpuMultA[103] = x80407;
  assign FpuMultA[104] = x80410;
  assign FpuMultA[105] = x80413;
  assign FpuMultA[106] = x80416;
  assign FpuMultA[107] = x80419;
  assign FpuMultA[108] = x80422;
  assign FpuMultA[109] = x80425;
  assign FpuMultA[110] = x80428;
  assign FpuMultA[111] = x80431;
  assign FpuMultA[112] = x80434;
  assign FpuMultA[113] = x80437;
  assign FpuMultA[114] = x80440;
  assign FpuMultA[115] = x80443;
  assign FpuMultA[116] = x80446;
  assign FpuMultA[117] = x80449;
  assign FpuMultA[118] = x80452;
  assign FpuMultA[119] = x80455;
  assign FpuMultA[120] = x80458;
  assign FpuMultA[121] = x80461;
  assign FpuMultA[122] = x80464;
  assign FpuMultA[123] = x80467;
  assign FpuMultA[124] = x80470;
  assign FpuMultA[125] = x80473;
  assign FpuMultA[126] = x80476;
  assign FpuMultA[127] = x80479;
  assign FpuMultB[0] = x67598;
  assign FpuMultB[1] = x67601;
  assign FpuMultB[2] = x67604;
  assign FpuMultB[3] = x67607;
  assign FpuMultB[4] = x67610;
  assign FpuMultB[5] = x67613;
  assign FpuMultB[6] = x67616;
  assign FpuMultB[7] = x67619;
  assign FpuMultB[8] = x67622;
  assign FpuMultB[9] = x67625;
  assign FpuMultB[10] = x67628;
  assign FpuMultB[11] = x67631;
  assign FpuMultB[12] = x67634;
  assign FpuMultB[13] = x67637;
  assign FpuMultB[14] = x67640;
  assign FpuMultB[15] = x67643;
  assign FpuMultB[16] = x67646;
  assign FpuMultB[17] = x67649;
  assign FpuMultB[18] = x67652;
  assign FpuMultB[19] = x67655;
  assign FpuMultB[20] = x67658;
  assign FpuMultB[21] = x67661;
  assign FpuMultB[22] = x67664;
  assign FpuMultB[23] = x67667;
  assign FpuMultB[24] = x67670;
  assign FpuMultB[25] = x67673;
  assign FpuMultB[26] = x67676;
  assign FpuMultB[27] = x67679;
  assign FpuMultB[28] = x67682;
  assign FpuMultB[29] = x67685;
  assign FpuMultB[30] = x67688;
  assign FpuMultB[31] = x67691;
  assign FpuMultB[32] = x67693;
  assign FpuMultB[33] = x67695;
  assign FpuMultB[34] = x67697;
  assign FpuMultB[35] = x67699;
  assign FpuMultB[36] = x67701;
  assign FpuMultB[37] = x67703;
  assign FpuMultB[38] = x67705;
  assign FpuMultB[39] = x67707;
  assign FpuMultB[40] = x67709;
  assign FpuMultB[41] = x67711;
  assign FpuMultB[42] = x67713;
  assign FpuMultB[43] = x67715;
  assign FpuMultB[44] = x67717;
  assign FpuMultB[45] = x67719;
  assign FpuMultB[46] = x67721;
  assign FpuMultB[47] = x67723;
  assign FpuMultB[48] = x67725;
  assign FpuMultB[49] = x67727;
  assign FpuMultB[50] = x67729;
  assign FpuMultB[51] = x67731;
  assign FpuMultB[52] = x67733;
  assign FpuMultB[53] = x67735;
  assign FpuMultB[54] = x67737;
  assign FpuMultB[55] = x67739;
  assign FpuMultB[56] = x67741;
  assign FpuMultB[57] = x67743;
  assign FpuMultB[58] = x67745;
  assign FpuMultB[59] = x67747;
  assign FpuMultB[60] = x67749;
  assign FpuMultB[61] = x67751;
  assign FpuMultB[62] = x67753;
  assign FpuMultB[63] = x67755;
  assign FpuMultB[64] = x67757;
  assign FpuMultB[65] = x67759;
  assign FpuMultB[66] = x67761;
  assign FpuMultB[67] = x67763;
  assign FpuMultB[68] = x67765;
  assign FpuMultB[69] = x67767;
  assign FpuMultB[70] = x67769;
  assign FpuMultB[71] = x67771;
  assign FpuMultB[72] = x67773;
  assign FpuMultB[73] = x67775;
  assign FpuMultB[74] = x67777;
  assign FpuMultB[75] = x67779;
  assign FpuMultB[76] = x67781;
  assign FpuMultB[77] = x67783;
  assign FpuMultB[78] = x67785;
  assign FpuMultB[79] = x67787;
  assign FpuMultB[80] = x67789;
  assign FpuMultB[81] = x67791;
  assign FpuMultB[82] = x67793;
  assign FpuMultB[83] = x67795;
  assign FpuMultB[84] = x67797;
  assign FpuMultB[85] = x67799;
  assign FpuMultB[86] = x67801;
  assign FpuMultB[87] = x67803;
  assign FpuMultB[88] = x67805;
  assign FpuMultB[89] = x67807;
  assign FpuMultB[90] = x67809;
  assign FpuMultB[91] = x67811;
  assign FpuMultB[92] = x67813;
  assign FpuMultB[93] = x67815;
  assign FpuMultB[94] = x67817;
  assign FpuMultB[95] = x67819;
  assign FpuMultB[96] = x67821;
  assign FpuMultB[97] = x67823;
  assign FpuMultB[98] = x67825;
  assign FpuMultB[99] = x67827;
  assign FpuMultB[100] = x67829;
  assign FpuMultB[101] = x67831;
  assign FpuMultB[102] = x67833;
  assign FpuMultB[103] = x67835;
  assign FpuMultB[104] = x67837;
  assign FpuMultB[105] = x67839;
  assign FpuMultB[106] = x67841;
  assign FpuMultB[107] = x67843;
  assign FpuMultB[108] = x67845;
  assign FpuMultB[109] = x67847;
  assign FpuMultB[110] = x67849;
  assign FpuMultB[111] = x67851;
  assign FpuMultB[112] = x67853;
  assign FpuMultB[113] = x67855;
  assign FpuMultB[114] = x67857;
  assign FpuMultB[115] = x67859;
  assign FpuMultB[116] = x67861;
  assign FpuMultB[117] = x67863;
  assign FpuMultB[118] = x67865;
  assign FpuMultB[119] = x67867;
  assign FpuMultB[120] = x67869;
  assign FpuMultB[121] = x67871;
  assign FpuMultB[122] = x67873;
  assign FpuMultB[123] = x67875;
  assign FpuMultB[124] = x67877;
  assign FpuMultB[125] = x67879;
  assign FpuMultB[126] = x67881;
  assign FpuMultB[127] = x67883;
  assign FpuMultOp[0] = x79462;
  assign FpuMultOp[1] = x79465;
  assign FpuMultOp[2] = x79468;
  assign FpuMultOp[3] = x79471;
  assign FpuMultOp[4] = x79474;
  assign FpuMultOp[5] = x79477;
  assign FpuMultStall = x68743;
  assign FpuMultValid = x83377;
  assign char_out = x64397;
  assign char_out_val[0] = x76834;
  assign char_out_val[1] = x76837;
  assign char_out_val[2] = x76840;
  assign char_out_val[3] = x76843;
  assign char_out_val[4] = x76846;
  assign char_out_val[5] = x76849;
  assign char_out_val[6] = x76852;
  assign reg00[0] = x2317;
  assign reg00[1] = x2321;
  assign reg00[2] = x2325;
  assign reg00[3] = x2329;
  assign reg00[4] = x2333;
  assign reg00[5] = x2337;
  assign reg00[6] = x2341;
  assign reg00[7] = x2345;
  assign reg00[8] = x2349;
  assign reg00[9] = x2353;
  assign reg00[10] = x2357;
  assign reg00[11] = x2361;
  assign reg00[12] = x2365;
  assign reg00[13] = x2369;
  assign reg00[14] = x2373;
  assign reg00[15] = x2377;
  assign reg00[16] = x2381;
  assign reg00[17] = x2385;
  assign reg00[18] = x2389;
  assign reg00[19] = x2393;
  assign reg00[20] = x2397;
  assign reg00[21] = x2401;
  assign reg00[22] = x2405;
  assign reg00[23] = x2409;
  assign reg00[24] = x2413;
  assign reg00[25] = x2417;
  assign reg00[26] = x2421;
  assign reg00[27] = x2425;
  assign reg00[28] = x2429;
  assign reg00[29] = x2433;
  assign reg00[30] = x2437;
  assign reg00[31] = x2441;
  assign reg01[0] = x2447;
  assign reg01[1] = x2451;
  assign reg01[2] = x2455;
  assign reg01[3] = x2459;
  assign reg01[4] = x2463;
  assign reg01[5] = x2467;
  assign reg01[6] = x2471;
  assign reg01[7] = x2475;
  assign reg01[8] = x2479;
  assign reg01[9] = x2483;
  assign reg01[10] = x2487;
  assign reg01[11] = x2491;
  assign reg01[12] = x2495;
  assign reg01[13] = x2499;
  assign reg01[14] = x2503;
  assign reg01[15] = x2507;
  assign reg01[16] = x2511;
  assign reg01[17] = x2515;
  assign reg01[18] = x2519;
  assign reg01[19] = x2523;
  assign reg01[20] = x2527;
  assign reg01[21] = x2531;
  assign reg01[22] = x2535;
  assign reg01[23] = x2539;
  assign reg01[24] = x2543;
  assign reg01[25] = x2547;
  assign reg01[26] = x2551;
  assign reg01[27] = x2555;
  assign reg01[28] = x2559;
  assign reg01[29] = x2563;
  assign reg01[30] = x2567;
  assign reg01[31] = x2571;
  assign reg02[0] = x2577;
  assign reg02[1] = x2581;
  assign reg02[2] = x2585;
  assign reg02[3] = x2589;
  assign reg02[4] = x2593;
  assign reg02[5] = x2597;
  assign reg02[6] = x2601;
  assign reg02[7] = x2605;
  assign reg02[8] = x2609;
  assign reg02[9] = x2613;
  assign reg02[10] = x2617;
  assign reg02[11] = x2621;
  assign reg02[12] = x2625;
  assign reg02[13] = x2629;
  assign reg02[14] = x2633;
  assign reg02[15] = x2637;
  assign reg02[16] = x2641;
  assign reg02[17] = x2645;
  assign reg02[18] = x2649;
  assign reg02[19] = x2653;
  assign reg02[20] = x2657;
  assign reg02[21] = x2661;
  assign reg02[22] = x2665;
  assign reg02[23] = x2669;
  assign reg02[24] = x2673;
  assign reg02[25] = x2677;
  assign reg02[26] = x2681;
  assign reg02[27] = x2685;
  assign reg02[28] = x2689;
  assign reg02[29] = x2693;
  assign reg02[30] = x2697;
  assign reg02[31] = x2701;
  assign reg03[0] = x2707;
  assign reg03[1] = x2711;
  assign reg03[2] = x2715;
  assign reg03[3] = x2719;
  assign reg03[4] = x2723;
  assign reg03[5] = x2727;
  assign reg03[6] = x2731;
  assign reg03[7] = x2735;
  assign reg03[8] = x2739;
  assign reg03[9] = x2743;
  assign reg03[10] = x2747;
  assign reg03[11] = x2751;
  assign reg03[12] = x2755;
  assign reg03[13] = x2759;
  assign reg03[14] = x2763;
  assign reg03[15] = x2767;
  assign reg03[16] = x2771;
  assign reg03[17] = x2775;
  assign reg03[18] = x2779;
  assign reg03[19] = x2783;
  assign reg03[20] = x2787;
  assign reg03[21] = x2791;
  assign reg03[22] = x2795;
  assign reg03[23] = x2799;
  assign reg03[24] = x2803;
  assign reg03[25] = x2807;
  assign reg03[26] = x2811;
  assign reg03[27] = x2815;
  assign reg03[28] = x2819;
  assign reg03[29] = x2823;
  assign reg03[30] = x2827;
  assign reg03[31] = x2831;
  assign reg04[0] = x2837;
  assign reg04[1] = x2841;
  assign reg04[2] = x2845;
  assign reg04[3] = x2849;
  assign reg04[4] = x2853;
  assign reg04[5] = x2857;
  assign reg04[6] = x2861;
  assign reg04[7] = x2865;
  assign reg04[8] = x2869;
  assign reg04[9] = x2873;
  assign reg04[10] = x2877;
  assign reg04[11] = x2881;
  assign reg04[12] = x2885;
  assign reg04[13] = x2889;
  assign reg04[14] = x2893;
  assign reg04[15] = x2897;
  assign reg04[16] = x2901;
  assign reg04[17] = x2905;
  assign reg04[18] = x2909;
  assign reg04[19] = x2913;
  assign reg04[20] = x2917;
  assign reg04[21] = x2921;
  assign reg04[22] = x2925;
  assign reg04[23] = x2929;
  assign reg04[24] = x2933;
  assign reg04[25] = x2937;
  assign reg04[26] = x2941;
  assign reg04[27] = x2945;
  assign reg04[28] = x2949;
  assign reg04[29] = x2953;
  assign reg04[30] = x2957;
  assign reg04[31] = x2961;
  assign reg05[0] = x2967;
  assign reg05[1] = x2971;
  assign reg05[2] = x2975;
  assign reg05[3] = x2979;
  assign reg05[4] = x2983;
  assign reg05[5] = x2987;
  assign reg05[6] = x2991;
  assign reg05[7] = x2995;
  assign reg05[8] = x2999;
  assign reg05[9] = x3003;
  assign reg05[10] = x3007;
  assign reg05[11] = x3011;
  assign reg05[12] = x3015;
  assign reg05[13] = x3019;
  assign reg05[14] = x3023;
  assign reg05[15] = x3027;
  assign reg05[16] = x3031;
  assign reg05[17] = x3035;
  assign reg05[18] = x3039;
  assign reg05[19] = x3043;
  assign reg05[20] = x3047;
  assign reg05[21] = x3051;
  assign reg05[22] = x3055;
  assign reg05[23] = x3059;
  assign reg05[24] = x3063;
  assign reg05[25] = x3067;
  assign reg05[26] = x3071;
  assign reg05[27] = x3075;
  assign reg05[28] = x3079;
  assign reg05[29] = x3083;
  assign reg05[30] = x3087;
  assign reg05[31] = x3091;
  assign reg06[0] = x3097;
  assign reg06[1] = x3101;
  assign reg06[2] = x3105;
  assign reg06[3] = x3109;
  assign reg06[4] = x3113;
  assign reg06[5] = x3117;
  assign reg06[6] = x3121;
  assign reg06[7] = x3125;
  assign reg06[8] = x3129;
  assign reg06[9] = x3133;
  assign reg06[10] = x3137;
  assign reg06[11] = x3141;
  assign reg06[12] = x3145;
  assign reg06[13] = x3149;
  assign reg06[14] = x3153;
  assign reg06[15] = x3157;
  assign reg06[16] = x3161;
  assign reg06[17] = x3165;
  assign reg06[18] = x3169;
  assign reg06[19] = x3173;
  assign reg06[20] = x3177;
  assign reg06[21] = x3181;
  assign reg06[22] = x3185;
  assign reg06[23] = x3189;
  assign reg06[24] = x3193;
  assign reg06[25] = x3197;
  assign reg06[26] = x3201;
  assign reg06[27] = x3205;
  assign reg06[28] = x3209;
  assign reg06[29] = x3213;
  assign reg06[30] = x3217;
  assign reg06[31] = x3221;
  assign reg07[0] = x3227;
  assign reg07[1] = x3231;
  assign reg07[2] = x3235;
  assign reg07[3] = x3239;
  assign reg07[4] = x3243;
  assign reg07[5] = x3247;
  assign reg07[6] = x3251;
  assign reg07[7] = x3255;
  assign reg07[8] = x3259;
  assign reg07[9] = x3263;
  assign reg07[10] = x3267;
  assign reg07[11] = x3271;
  assign reg07[12] = x3275;
  assign reg07[13] = x3279;
  assign reg07[14] = x3283;
  assign reg07[15] = x3287;
  assign reg07[16] = x3291;
  assign reg07[17] = x3295;
  assign reg07[18] = x3299;
  assign reg07[19] = x3303;
  assign reg07[20] = x3307;
  assign reg07[21] = x3311;
  assign reg07[22] = x3315;
  assign reg07[23] = x3319;
  assign reg07[24] = x3323;
  assign reg07[25] = x3327;
  assign reg07[26] = x3331;
  assign reg07[27] = x3335;
  assign reg07[28] = x3339;
  assign reg07[29] = x3343;
  assign reg07[30] = x3347;
  assign reg07[31] = x3351;

  assign x87265 = 0;

  assign ram_w0 = x63875;
  assign ram_qa0[0] = x63757;
  assign ram_da0[0] = x63757;
  assign ram_qa0[1] = x63762;
  assign ram_da0[1] = x63762;
  assign ram_qa0[2] = x63766;
  assign ram_da0[2] = x63766;
  assign ram_qa0[3] = x63771;
  assign ram_da0[3] = x63771;
  assign ram_qa0[4] = x63776;
  assign ram_da0[4] = x63776;
  assign ram_qa0[5] = x63781;
  assign ram_da0[5] = x63781;
  assign ram_qa0[6] = x63785;
  assign ram_da0[6] = x63785;
  assign ram_qa0[7] = x63790;
  assign ram_da0[7] = x63790;
  assign ram_d0[0] = x76834;
  assign ram_d0[1] = x76837;
  assign ram_d0[2] = x76840;
  assign ram_d0[3] = x76843;
  assign ram_d0[4] = x76846;
  assign ram_d0[5] = x76849;
  assign ram_d0[6] = x76852;
  assign ram_d0[7] = x76855;
  assign ram_d0[8] = x76858;
  assign ram_d0[9] = x76861;
  assign ram_d0[10] = x76864;
  assign ram_d0[11] = x76867;
  assign ram_d0[12] = x76870;
  assign ram_d0[13] = x76873;
  assign ram_d0[14] = x76876;
  assign ram_d0[15] = x76879;
  assign ram_d0[16] = x76882;
  assign ram_d0[17] = x76885;
  assign ram_d0[18] = x76888;
  assign ram_d0[19] = x76891;
  assign ram_d0[20] = x76894;
  assign ram_d0[21] = x76897;
  assign ram_d0[22] = x76900;
  assign ram_d0[23] = x76903;
  assign ram_d0[24] = x76906;
  assign ram_d0[25] = x76909;
  assign ram_d0[26] = x76912;
  assign ram_d0[27] = x76915;
  assign ram_d0[28] = x76918;
  assign ram_d0[29] = x76921;
  assign ram_d0[30] = x76924;
  assign ram_d0[31] = x76927;
  assign x63876 = ram_q0[0];
  assign x63877 = ram_q0[1];
  assign x63878 = ram_q0[2];
  assign x63879 = ram_q0[3];
  assign x63880 = ram_q0[4];
  assign x63881 = ram_q0[5];
  assign x63882 = ram_q0[6];
  assign x63883 = ram_q0[7];
  assign x63884 = ram_q0[8];
  assign x63885 = ram_q0[9];
  assign x63886 = ram_q0[10];
  assign x63887 = ram_q0[11];
  assign x63888 = ram_q0[12];
  assign x63889 = ram_q0[13];
  assign x63890 = ram_q0[14];
  assign x63891 = ram_q0[15];
  assign x63892 = ram_q0[16];
  assign x63893 = ram_q0[17];
  assign x63894 = ram_q0[18];
  assign x63895 = ram_q0[19];
  assign x63896 = ram_q0[20];
  assign x63897 = ram_q0[21];
  assign x63898 = ram_q0[22];
  assign x63899 = ram_q0[23];
  assign x63900 = ram_q0[24];
  assign x63901 = ram_q0[25];
  assign x63902 = ram_q0[26];
  assign x63903 = ram_q0[27];
  assign x63904 = ram_q0[28];
  assign x63905 = ram_q0[29];
  assign x63906 = ram_q0[30];
  assign x63907 = ram_q0[31];
  assign ram_w1 = x63875;
  assign ram_qa1[0] = x64574;
  assign ram_da1[0] = x64574;
  assign ram_qa1[1] = x64579;
  assign ram_da1[1] = x64579;
  assign ram_qa1[2] = x64583;
  assign ram_da1[2] = x64583;
  assign ram_qa1[3] = x64588;
  assign ram_da1[3] = x64588;
  assign ram_qa1[4] = x64593;
  assign ram_da1[4] = x64593;
  assign ram_qa1[5] = x64598;
  assign ram_da1[5] = x64598;
  assign ram_qa1[6] = x64602;
  assign ram_da1[6] = x64602;
  assign ram_qa1[7] = x64607;
  assign ram_da1[7] = x64607;
  assign ram_d1[0] = x77128;
  assign ram_d1[1] = x77131;
  assign ram_d1[2] = x77134;
  assign ram_d1[3] = x77137;
  assign ram_d1[4] = x77140;
  assign ram_d1[5] = x77143;
  assign ram_d1[6] = x77146;
  assign ram_d1[7] = x77149;
  assign ram_d1[8] = x77152;
  assign ram_d1[9] = x77155;
  assign ram_d1[10] = x77158;
  assign ram_d1[11] = x77161;
  assign ram_d1[12] = x77164;
  assign ram_d1[13] = x77167;
  assign ram_d1[14] = x77170;
  assign ram_d1[15] = x77173;
  assign ram_d1[16] = x77176;
  assign ram_d1[17] = x77179;
  assign ram_d1[18] = x77182;
  assign ram_d1[19] = x77185;
  assign ram_d1[20] = x77188;
  assign ram_d1[21] = x77191;
  assign ram_d1[22] = x77194;
  assign ram_d1[23] = x77197;
  assign ram_d1[24] = x77200;
  assign ram_d1[25] = x77203;
  assign ram_d1[26] = x77206;
  assign ram_d1[27] = x77209;
  assign ram_d1[28] = x77212;
  assign ram_d1[29] = x77215;
  assign ram_d1[30] = x77218;
  assign ram_d1[31] = x77221;
  assign x64608 = ram_q1[0];
  assign x64609 = ram_q1[1];
  assign x64610 = ram_q1[2];
  assign x64611 = ram_q1[3];
  assign x64612 = ram_q1[4];
  assign x64613 = ram_q1[5];
  assign x64614 = ram_q1[6];
  assign x64615 = ram_q1[7];
  assign x64616 = ram_q1[8];
  assign x64617 = ram_q1[9];
  assign x64618 = ram_q1[10];
  assign x64619 = ram_q1[11];
  assign x64620 = ram_q1[12];
  assign x64621 = ram_q1[13];
  assign x64622 = ram_q1[14];
  assign x64623 = ram_q1[15];
  assign x64624 = ram_q1[16];
  assign x64625 = ram_q1[17];
  assign x64626 = ram_q1[18];
  assign x64627 = ram_q1[19];
  assign x64628 = ram_q1[20];
  assign x64629 = ram_q1[21];
  assign x64630 = ram_q1[22];
  assign x64631 = ram_q1[23];
  assign x64632 = ram_q1[24];
  assign x64633 = ram_q1[25];
  assign x64634 = ram_q1[26];
  assign x64635 = ram_q1[27];
  assign x64636 = ram_q1[28];
  assign x64637 = ram_q1[29];
  assign x64638 = ram_q1[30];
  assign x64639 = ram_q1[31];
  assign ram_w2 = x63875;
  assign ram_qa2[0] = x65244;
  assign ram_da2[0] = x65244;
  assign ram_qa2[1] = x65249;
  assign ram_da2[1] = x65249;
  assign ram_qa2[2] = x65253;
  assign ram_da2[2] = x65253;
  assign ram_qa2[3] = x65258;
  assign ram_da2[3] = x65258;
  assign ram_qa2[4] = x65263;
  assign ram_da2[4] = x65263;
  assign ram_qa2[5] = x65268;
  assign ram_da2[5] = x65268;
  assign ram_qa2[6] = x65272;
  assign ram_da2[6] = x65272;
  assign ram_qa2[7] = x65277;
  assign ram_da2[7] = x65277;
  assign ram_d2[0] = x77422;
  assign ram_d2[1] = x77425;
  assign ram_d2[2] = x77428;
  assign ram_d2[3] = x77431;
  assign ram_d2[4] = x77434;
  assign ram_d2[5] = x77437;
  assign ram_d2[6] = x77440;
  assign ram_d2[7] = x77443;
  assign ram_d2[8] = x77446;
  assign ram_d2[9] = x77449;
  assign ram_d2[10] = x77452;
  assign ram_d2[11] = x77455;
  assign ram_d2[12] = x77458;
  assign ram_d2[13] = x77461;
  assign ram_d2[14] = x77464;
  assign ram_d2[15] = x77467;
  assign ram_d2[16] = x77470;
  assign ram_d2[17] = x77473;
  assign ram_d2[18] = x77476;
  assign ram_d2[19] = x77479;
  assign ram_d2[20] = x77482;
  assign ram_d2[21] = x77485;
  assign ram_d2[22] = x77488;
  assign ram_d2[23] = x77491;
  assign ram_d2[24] = x77494;
  assign ram_d2[25] = x77497;
  assign ram_d2[26] = x77500;
  assign ram_d2[27] = x77503;
  assign ram_d2[28] = x77506;
  assign ram_d2[29] = x77509;
  assign ram_d2[30] = x77512;
  assign ram_d2[31] = x77515;
  assign x65278 = ram_q2[0];
  assign x65279 = ram_q2[1];
  assign x65280 = ram_q2[2];
  assign x65281 = ram_q2[3];
  assign x65282 = ram_q2[4];
  assign x65283 = ram_q2[5];
  assign x65284 = ram_q2[6];
  assign x65285 = ram_q2[7];
  assign x65286 = ram_q2[8];
  assign x65287 = ram_q2[9];
  assign x65288 = ram_q2[10];
  assign x65289 = ram_q2[11];
  assign x65290 = ram_q2[12];
  assign x65291 = ram_q2[13];
  assign x65292 = ram_q2[14];
  assign x65293 = ram_q2[15];
  assign x65294 = ram_q2[16];
  assign x65295 = ram_q2[17];
  assign x65296 = ram_q2[18];
  assign x65297 = ram_q2[19];
  assign x65298 = ram_q2[20];
  assign x65299 = ram_q2[21];
  assign x65300 = ram_q2[22];
  assign x65301 = ram_q2[23];
  assign x65302 = ram_q2[24];
  assign x65303 = ram_q2[25];
  assign x65304 = ram_q2[26];
  assign x65305 = ram_q2[27];
  assign x65306 = ram_q2[28];
  assign x65307 = ram_q2[29];
  assign x65308 = ram_q2[30];
  assign x65309 = ram_q2[31];
  assign ram_w3 = x63875;
  assign ram_qa3[0] = x65914;
  assign ram_da3[0] = x65914;
  assign ram_qa3[1] = x65919;
  assign ram_da3[1] = x65919;
  assign ram_qa3[2] = x65923;
  assign ram_da3[2] = x65923;
  assign ram_qa3[3] = x65928;
  assign ram_da3[3] = x65928;
  assign ram_qa3[4] = x65933;
  assign ram_da3[4] = x65933;
  assign ram_qa3[5] = x65938;
  assign ram_da3[5] = x65938;
  assign ram_qa3[6] = x65942;
  assign ram_da3[6] = x65942;
  assign ram_qa3[7] = x65947;
  assign ram_da3[7] = x65947;
  assign ram_d3[0] = x77716;
  assign ram_d3[1] = x77719;
  assign ram_d3[2] = x77722;
  assign ram_d3[3] = x77725;
  assign ram_d3[4] = x77728;
  assign ram_d3[5] = x77731;
  assign ram_d3[6] = x77734;
  assign ram_d3[7] = x77737;
  assign ram_d3[8] = x77740;
  assign ram_d3[9] = x77743;
  assign ram_d3[10] = x77746;
  assign ram_d3[11] = x77749;
  assign ram_d3[12] = x77752;
  assign ram_d3[13] = x77755;
  assign ram_d3[14] = x77758;
  assign ram_d3[15] = x77761;
  assign ram_d3[16] = x77764;
  assign ram_d3[17] = x77767;
  assign ram_d3[18] = x77770;
  assign ram_d3[19] = x77773;
  assign ram_d3[20] = x77776;
  assign ram_d3[21] = x77779;
  assign ram_d3[22] = x77782;
  assign ram_d3[23] = x77785;
  assign ram_d3[24] = x77788;
  assign ram_d3[25] = x77791;
  assign ram_d3[26] = x77794;
  assign ram_d3[27] = x77797;
  assign ram_d3[28] = x77800;
  assign ram_d3[29] = x77803;
  assign ram_d3[30] = x77806;
  assign ram_d3[31] = x77809;
  assign x65948 = ram_q3[0];
  assign x65949 = ram_q3[1];
  assign x65950 = ram_q3[2];
  assign x65951 = ram_q3[3];
  assign x65952 = ram_q3[4];
  assign x65953 = ram_q3[5];
  assign x65954 = ram_q3[6];
  assign x65955 = ram_q3[7];
  assign x65956 = ram_q3[8];
  assign x65957 = ram_q3[9];
  assign x65958 = ram_q3[10];
  assign x65959 = ram_q3[11];
  assign x65960 = ram_q3[12];
  assign x65961 = ram_q3[13];
  assign x65962 = ram_q3[14];
  assign x65963 = ram_q3[15];
  assign x65964 = ram_q3[16];
  assign x65965 = ram_q3[17];
  assign x65966 = ram_q3[18];
  assign x65967 = ram_q3[19];
  assign x65968 = ram_q3[20];
  assign x65969 = ram_q3[21];
  assign x65970 = ram_q3[22];
  assign x65971 = ram_q3[23];
  assign x65972 = ram_q3[24];
  assign x65973 = ram_q3[25];
  assign x65974 = ram_q3[26];
  assign x65975 = ram_q3[27];
  assign x65976 = ram_q3[28];
  assign x65977 = ram_q3[29];
  assign x65978 = ram_q3[30];
  assign x65979 = ram_q3[31];

  initial
    begin
      x58 <= 0;
      x59 <= 0;
      x60 <= 0;
      x61 <= 0;
      x62 <= 0;
      x63 <= 0;
      x602 <= 0;
      x603 <= 0;
      x604 <= 0;
      x605 <= 0;
      x606 <= 0;
      x607 <= 0;
      x608 <= 0;
      x609 <= 0;
      x610 <= 0;
      x611 <= 0;
      x612 <= 0;
      x613 <= 0;
      x614 <= 0;
      x615 <= 0;
      x616 <= 0;
      x617 <= 0;
      x618 <= 0;
      x619 <= 0;
      x620 <= 0;
      x621 <= 0;
      x622 <= 0;
      x623 <= 0;
      x624 <= 0;
      x625 <= 0;
      x626 <= 0;
      x627 <= 0;
      x628 <= 0;
      x629 <= 0;
      x630 <= 0;
      x631 <= 0;
      x632 <= 0;
      x633 <= 0;
      x674 <= 0;
      x675 <= 0;
      x676 <= 0;
      x677 <= 0;
      x1232 <= 0;
      x1238 <= 0;
      x1244 <= 0;
      x1250 <= 0;
      x1256 <= 0;
      x1262 <= 0;
      x1268 <= 0;
      x1274 <= 0;
      x1281 <= 0;
      x1288 <= 0;
      x1294 <= 0;
      x1300 <= 0;
      x1306 <= 0;
      x1312 <= 0;
      x1318 <= 0;
      x1324 <= 0;
      x1330 <= 0;
      x1336 <= 0;
      x1342 <= 0;
      x1348 <= 0;
      x1354 <= 0;
      x1360 <= 0;
      x1366 <= 0;
      x1372 <= 0;
      x1379 <= 0;
      x1386 <= 0;
      x1392 <= 0;
      x1398 <= 0;
      x1404 <= 0;
      x1410 <= 0;
      x1416 <= 0;
      x1422 <= 0;
      x1758 <= 0;
      x1768 <= 0;
      x1778 <= 0;
      x1788 <= 0;
      x1798 <= 0;
      x1808 <= 0;
      x1818 <= 0;
      x1828 <= 0;
      x1914 <= 0;
      x1918 <= 0;
      x1922 <= 0;
      x1926 <= 0;
      x1930 <= 0;
      x1934 <= 0;
      x1940 <= 0;
      x1944 <= 0;
      x1948 <= 0;
      x1952 <= 0;
      x1956 <= 0;
      x1960 <= 0;
      x1966 <= 0;
      x1970 <= 0;
      x1974 <= 0;
      x1978 <= 0;
      x1982 <= 0;
      x1986 <= 0;
      x1992 <= 0;
      x1996 <= 0;
      x2000 <= 0;
      x2004 <= 0;
      x2008 <= 0;
      x2012 <= 0;
      x2018 <= 0;
      x2022 <= 0;
      x2026 <= 0;
      x2030 <= 0;
      x2034 <= 0;
      x2038 <= 0;
      x2044 <= 0;
      x2048 <= 0;
      x2052 <= 0;
      x2056 <= 0;
      x2060 <= 0;
      x2064 <= 0;
      x2070 <= 0;
      x2074 <= 0;
      x2078 <= 0;
      x2082 <= 0;
      x2086 <= 0;
      x2090 <= 0;
      x2096 <= 0;
      x2100 <= 0;
      x2104 <= 0;
      x2108 <= 0;
      x2112 <= 0;
      x2116 <= 0;
      x2317 <= 0;
      x2321 <= 0;
      x2325 <= 0;
      x2329 <= 0;
      x2333 <= 0;
      x2337 <= 0;
      x2341 <= 0;
      x2345 <= 0;
      x2349 <= 0;
      x2353 <= 0;
      x2357 <= 0;
      x2361 <= 0;
      x2365 <= 0;
      x2369 <= 0;
      x2373 <= 0;
      x2377 <= 0;
      x2381 <= 0;
      x2385 <= 0;
      x2389 <= 0;
      x2393 <= 0;
      x2397 <= 0;
      x2401 <= 0;
      x2405 <= 0;
      x2409 <= 0;
      x2413 <= 0;
      x2417 <= 0;
      x2421 <= 0;
      x2425 <= 0;
      x2429 <= 0;
      x2433 <= 0;
      x2437 <= 0;
      x2441 <= 0;
      x2447 <= 0;
      x2451 <= 0;
      x2455 <= 0;
      x2459 <= 0;
      x2463 <= 0;
      x2467 <= 0;
      x2471 <= 0;
      x2475 <= 0;
      x2479 <= 0;
      x2483 <= 0;
      x2487 <= 0;
      x2491 <= 0;
      x2495 <= 0;
      x2499 <= 0;
      x2503 <= 0;
      x2507 <= 0;
      x2511 <= 0;
      x2515 <= 0;
      x2519 <= 0;
      x2523 <= 0;
      x2527 <= 0;
      x2531 <= 0;
      x2535 <= 0;
      x2539 <= 0;
      x2543 <= 0;
      x2547 <= 0;
      x2551 <= 0;
      x2555 <= 0;
      x2559 <= 0;
      x2563 <= 0;
      x2567 <= 0;
      x2571 <= 0;
      x2577 <= 0;
      x2581 <= 0;
      x2585 <= 0;
      x2589 <= 0;
      x2593 <= 0;
      x2597 <= 0;
      x2601 <= 0;
      x2605 <= 0;
      x2609 <= 0;
      x2613 <= 0;
      x2617 <= 0;
      x2621 <= 0;
      x2625 <= 0;
      x2629 <= 0;
      x2633 <= 0;
      x2637 <= 0;
      x2641 <= 0;
      x2645 <= 0;
      x2649 <= 0;
      x2653 <= 0;
      x2657 <= 0;
      x2661 <= 0;
      x2665 <= 0;
      x2669 <= 0;
      x2673 <= 0;
      x2677 <= 0;
      x2681 <= 0;
      x2685 <= 0;
      x2689 <= 0;
      x2693 <= 0;
      x2697 <= 0;
      x2701 <= 0;
      x2707 <= 0;
      x2711 <= 0;
      x2715 <= 0;
      x2719 <= 0;
      x2723 <= 0;
      x2727 <= 0;
      x2731 <= 0;
      x2735 <= 0;
      x2739 <= 0;
      x2743 <= 0;
      x2747 <= 0;
      x2751 <= 0;
      x2755 <= 0;
      x2759 <= 0;
      x2763 <= 0;
      x2767 <= 0;
      x2771 <= 0;
      x2775 <= 0;
      x2779 <= 0;
      x2783 <= 0;
      x2787 <= 0;
      x2791 <= 0;
      x2795 <= 0;
      x2799 <= 0;
      x2803 <= 0;
      x2807 <= 0;
      x2811 <= 0;
      x2815 <= 0;
      x2819 <= 0;
      x2823 <= 0;
      x2827 <= 0;
      x2831 <= 0;
      x2837 <= 0;
      x2841 <= 0;
      x2845 <= 0;
      x2849 <= 0;
      x2853 <= 0;
      x2857 <= 0;
      x2861 <= 0;
      x2865 <= 0;
      x2869 <= 0;
      x2873 <= 0;
      x2877 <= 0;
      x2881 <= 0;
      x2885 <= 0;
      x2889 <= 0;
      x2893 <= 0;
      x2897 <= 0;
      x2901 <= 0;
      x2905 <= 0;
      x2909 <= 0;
      x2913 <= 0;
      x2917 <= 0;
      x2921 <= 0;
      x2925 <= 0;
      x2929 <= 0;
      x2933 <= 0;
      x2937 <= 0;
      x2941 <= 0;
      x2945 <= 0;
      x2949 <= 0;
      x2953 <= 0;
      x2957 <= 0;
      x2961 <= 0;
      x2967 <= 0;
      x2971 <= 0;
      x2975 <= 0;
      x2979 <= 0;
      x2983 <= 0;
      x2987 <= 0;
      x2991 <= 0;
      x2995 <= 0;
      x2999 <= 0;
      x3003 <= 0;
      x3007 <= 0;
      x3011 <= 0;
      x3015 <= 0;
      x3019 <= 0;
      x3023 <= 0;
      x3027 <= 0;
      x3031 <= 0;
      x3035 <= 0;
      x3039 <= 0;
      x3043 <= 0;
      x3047 <= 0;
      x3051 <= 0;
      x3055 <= 0;
      x3059 <= 0;
      x3063 <= 0;
      x3067 <= 0;
      x3071 <= 0;
      x3075 <= 0;
      x3079 <= 0;
      x3083 <= 0;
      x3087 <= 0;
      x3091 <= 0;
      x3097 <= 0;
      x3101 <= 0;
      x3105 <= 0;
      x3109 <= 0;
      x3113 <= 0;
      x3117 <= 0;
      x3121 <= 0;
      x3125 <= 0;
      x3129 <= 0;
      x3133 <= 0;
      x3137 <= 0;
      x3141 <= 0;
      x3145 <= 0;
      x3149 <= 0;
      x3153 <= 0;
      x3157 <= 0;
      x3161 <= 0;
      x3165 <= 0;
      x3169 <= 0;
      x3173 <= 0;
      x3177 <= 0;
      x3181 <= 0;
      x3185 <= 0;
      x3189 <= 0;
      x3193 <= 0;
      x3197 <= 0;
      x3201 <= 0;
      x3205 <= 0;
      x3209 <= 0;
      x3213 <= 0;
      x3217 <= 0;
      x3221 <= 0;
      x3227 <= 0;
      x3231 <= 0;
      x3235 <= 0;
      x3239 <= 0;
      x3243 <= 0;
      x3247 <= 0;
      x3251 <= 0;
      x3255 <= 0;
      x3259 <= 0;
      x3263 <= 0;
      x3267 <= 0;
      x3271 <= 0;
      x3275 <= 0;
      x3279 <= 0;
      x3283 <= 0;
      x3287 <= 0;
      x3291 <= 0;
      x3295 <= 0;
      x3299 <= 0;
      x3303 <= 0;
      x3307 <= 0;
      x3311 <= 0;
      x3315 <= 0;
      x3319 <= 0;
      x3323 <= 0;
      x3327 <= 0;
      x3331 <= 0;
      x3335 <= 0;
      x3339 <= 0;
      x3343 <= 0;
      x3347 <= 0;
      x3351 <= 0;
      x3358 <= 0;
      x3363 <= 0;
      x3367 <= 0;
      x3371 <= 0;
      x3375 <= 0;
      x3379 <= 0;
      x3383 <= 0;
      x3387 <= 0;
      x3391 <= 0;
      x3395 <= 0;
      x3399 <= 0;
      x3403 <= 0;
      x3407 <= 0;
      x3411 <= 0;
      x3415 <= 0;
      x3419 <= 0;
      x3423 <= 0;
      x3427 <= 0;
      x3431 <= 0;
      x3435 <= 0;
      x3439 <= 0;
      x3443 <= 0;
      x3447 <= 0;
      x3451 <= 0;
      x3455 <= 0;
      x3459 <= 0;
      x3463 <= 0;
      x3467 <= 0;
      x3471 <= 0;
      x3475 <= 0;
      x3479 <= 0;
      x3483 <= 0;
      x3489 <= 0;
      x3493 <= 0;
      x3497 <= 0;
      x3501 <= 0;
      x3505 <= 0;
      x3509 <= 0;
      x3513 <= 0;
      x3517 <= 0;
      x3521 <= 0;
      x3525 <= 0;
      x3529 <= 0;
      x3533 <= 0;
      x3537 <= 0;
      x3541 <= 0;
      x3545 <= 0;
      x3549 <= 0;
      x3553 <= 0;
      x3557 <= 0;
      x3561 <= 0;
      x3565 <= 0;
      x3569 <= 0;
      x3573 <= 0;
      x3577 <= 0;
      x3581 <= 0;
      x3585 <= 0;
      x3589 <= 0;
      x3593 <= 0;
      x3597 <= 0;
      x3601 <= 0;
      x3605 <= 0;
      x3609 <= 0;
      x3613 <= 0;
      x3619 <= 0;
      x3623 <= 0;
      x3627 <= 0;
      x3631 <= 0;
      x3635 <= 0;
      x3639 <= 0;
      x3643 <= 0;
      x3647 <= 0;
      x3651 <= 0;
      x3655 <= 0;
      x3659 <= 0;
      x3663 <= 0;
      x3667 <= 0;
      x3671 <= 0;
      x3675 <= 0;
      x3679 <= 0;
      x3683 <= 0;
      x3687 <= 0;
      x3691 <= 0;
      x3695 <= 0;
      x3699 <= 0;
      x3703 <= 0;
      x3707 <= 0;
      x3711 <= 0;
      x3715 <= 0;
      x3719 <= 0;
      x3723 <= 0;
      x3727 <= 0;
      x3731 <= 0;
      x3735 <= 0;
      x3739 <= 0;
      x3743 <= 0;
      x3749 <= 0;
      x3753 <= 0;
      x3757 <= 0;
      x3761 <= 0;
      x3765 <= 0;
      x3769 <= 0;
      x3773 <= 0;
      x3777 <= 0;
      x3781 <= 0;
      x3785 <= 0;
      x3789 <= 0;
      x3793 <= 0;
      x3797 <= 0;
      x3801 <= 0;
      x3805 <= 0;
      x3809 <= 0;
      x3813 <= 0;
      x3817 <= 0;
      x3821 <= 0;
      x3825 <= 0;
      x3829 <= 0;
      x3833 <= 0;
      x3837 <= 0;
      x3841 <= 0;
      x3845 <= 0;
      x3849 <= 0;
      x3853 <= 0;
      x3857 <= 0;
      x3861 <= 0;
      x3865 <= 0;
      x3869 <= 0;
      x3873 <= 0;
      x3879 <= 0;
      x3883 <= 0;
      x3887 <= 0;
      x3891 <= 0;
      x3895 <= 0;
      x3899 <= 0;
      x3903 <= 0;
      x3907 <= 0;
      x3911 <= 0;
      x3915 <= 0;
      x3919 <= 0;
      x3923 <= 0;
      x3927 <= 0;
      x3931 <= 0;
      x3935 <= 0;
      x3939 <= 0;
      x3943 <= 0;
      x3947 <= 0;
      x3951 <= 0;
      x3955 <= 0;
      x3959 <= 0;
      x3963 <= 0;
      x3967 <= 0;
      x3971 <= 0;
      x3975 <= 0;
      x3979 <= 0;
      x3983 <= 0;
      x3987 <= 0;
      x3991 <= 0;
      x3995 <= 0;
      x3999 <= 0;
      x4003 <= 0;
      x4009 <= 0;
      x4013 <= 0;
      x4017 <= 0;
      x4021 <= 0;
      x4025 <= 0;
      x4029 <= 0;
      x4033 <= 0;
      x4037 <= 0;
      x4041 <= 0;
      x4045 <= 0;
      x4049 <= 0;
      x4053 <= 0;
      x4057 <= 0;
      x4061 <= 0;
      x4065 <= 0;
      x4069 <= 0;
      x4073 <= 0;
      x4077 <= 0;
      x4081 <= 0;
      x4085 <= 0;
      x4089 <= 0;
      x4093 <= 0;
      x4097 <= 0;
      x4101 <= 0;
      x4105 <= 0;
      x4109 <= 0;
      x4113 <= 0;
      x4117 <= 0;
      x4121 <= 0;
      x4125 <= 0;
      x4129 <= 0;
      x4133 <= 0;
      x4139 <= 0;
      x4143 <= 0;
      x4147 <= 0;
      x4151 <= 0;
      x4155 <= 0;
      x4159 <= 0;
      x4163 <= 0;
      x4167 <= 0;
      x4171 <= 0;
      x4175 <= 0;
      x4179 <= 0;
      x4183 <= 0;
      x4187 <= 0;
      x4191 <= 0;
      x4195 <= 0;
      x4199 <= 0;
      x4203 <= 0;
      x4207 <= 0;
      x4211 <= 0;
      x4215 <= 0;
      x4219 <= 0;
      x4223 <= 0;
      x4227 <= 0;
      x4231 <= 0;
      x4235 <= 0;
      x4239 <= 0;
      x4243 <= 0;
      x4247 <= 0;
      x4251 <= 0;
      x4255 <= 0;
      x4259 <= 0;
      x4263 <= 0;
      x4269 <= 0;
      x4273 <= 0;
      x4277 <= 0;
      x4281 <= 0;
      x4285 <= 0;
      x4289 <= 0;
      x4293 <= 0;
      x4297 <= 0;
      x4301 <= 0;
      x4305 <= 0;
      x4309 <= 0;
      x4313 <= 0;
      x4317 <= 0;
      x4321 <= 0;
      x4325 <= 0;
      x4329 <= 0;
      x4333 <= 0;
      x4337 <= 0;
      x4341 <= 0;
      x4345 <= 0;
      x4349 <= 0;
      x4353 <= 0;
      x4357 <= 0;
      x4361 <= 0;
      x4365 <= 0;
      x4369 <= 0;
      x4373 <= 0;
      x4377 <= 0;
      x4381 <= 0;
      x4385 <= 0;
      x4389 <= 0;
      x4393 <= 0;
      x4399 <= 0;
      x4404 <= 0;
      x4409 <= 0;
      x4413 <= 0;
      x4417 <= 0;
      x4421 <= 0;
      x4425 <= 0;
      x4429 <= 0;
      x4433 <= 0;
      x4437 <= 0;
      x4441 <= 0;
      x4445 <= 0;
      x4449 <= 0;
      x4453 <= 0;
      x4457 <= 0;
      x4461 <= 0;
      x4465 <= 0;
      x4469 <= 0;
      x4473 <= 0;
      x4477 <= 0;
      x4481 <= 0;
      x4485 <= 0;
      x4489 <= 0;
      x4493 <= 0;
      x4497 <= 0;
      x4501 <= 0;
      x4505 <= 0;
      x4509 <= 0;
      x4513 <= 0;
      x4517 <= 0;
      x4521 <= 0;
      x4525 <= 0;
      x4531 <= 0;
      x4535 <= 0;
      x4539 <= 0;
      x4543 <= 0;
      x4547 <= 0;
      x4551 <= 0;
      x4555 <= 0;
      x4559 <= 0;
      x4563 <= 0;
      x4567 <= 0;
      x4571 <= 0;
      x4575 <= 0;
      x4579 <= 0;
      x4583 <= 0;
      x4587 <= 0;
      x4591 <= 0;
      x4595 <= 0;
      x4599 <= 0;
      x4603 <= 0;
      x4607 <= 0;
      x4611 <= 0;
      x4615 <= 0;
      x4619 <= 0;
      x4623 <= 0;
      x4627 <= 0;
      x4631 <= 0;
      x4635 <= 0;
      x4639 <= 0;
      x4643 <= 0;
      x4647 <= 0;
      x4651 <= 0;
      x4655 <= 0;
      x4661 <= 0;
      x4665 <= 0;
      x4669 <= 0;
      x4673 <= 0;
      x4677 <= 0;
      x4681 <= 0;
      x4685 <= 0;
      x4689 <= 0;
      x4693 <= 0;
      x4697 <= 0;
      x4701 <= 0;
      x4705 <= 0;
      x4709 <= 0;
      x4713 <= 0;
      x4717 <= 0;
      x4721 <= 0;
      x4725 <= 0;
      x4729 <= 0;
      x4733 <= 0;
      x4737 <= 0;
      x4741 <= 0;
      x4745 <= 0;
      x4749 <= 0;
      x4753 <= 0;
      x4757 <= 0;
      x4761 <= 0;
      x4765 <= 0;
      x4769 <= 0;
      x4773 <= 0;
      x4777 <= 0;
      x4781 <= 0;
      x4785 <= 0;
      x4791 <= 0;
      x4795 <= 0;
      x4799 <= 0;
      x4803 <= 0;
      x4807 <= 0;
      x4811 <= 0;
      x4815 <= 0;
      x4819 <= 0;
      x4823 <= 0;
      x4827 <= 0;
      x4831 <= 0;
      x4835 <= 0;
      x4839 <= 0;
      x4843 <= 0;
      x4847 <= 0;
      x4851 <= 0;
      x4855 <= 0;
      x4859 <= 0;
      x4863 <= 0;
      x4867 <= 0;
      x4871 <= 0;
      x4875 <= 0;
      x4879 <= 0;
      x4883 <= 0;
      x4887 <= 0;
      x4891 <= 0;
      x4895 <= 0;
      x4899 <= 0;
      x4903 <= 0;
      x4907 <= 0;
      x4911 <= 0;
      x4915 <= 0;
      x4921 <= 0;
      x4925 <= 0;
      x4929 <= 0;
      x4933 <= 0;
      x4937 <= 0;
      x4941 <= 0;
      x4945 <= 0;
      x4949 <= 0;
      x4953 <= 0;
      x4957 <= 0;
      x4961 <= 0;
      x4965 <= 0;
      x4969 <= 0;
      x4973 <= 0;
      x4977 <= 0;
      x4981 <= 0;
      x4985 <= 0;
      x4989 <= 0;
      x4993 <= 0;
      x4997 <= 0;
      x5001 <= 0;
      x5005 <= 0;
      x5009 <= 0;
      x5013 <= 0;
      x5017 <= 0;
      x5021 <= 0;
      x5025 <= 0;
      x5029 <= 0;
      x5033 <= 0;
      x5037 <= 0;
      x5041 <= 0;
      x5045 <= 0;
      x5051 <= 0;
      x5055 <= 0;
      x5059 <= 0;
      x5063 <= 0;
      x5067 <= 0;
      x5071 <= 0;
      x5075 <= 0;
      x5079 <= 0;
      x5083 <= 0;
      x5087 <= 0;
      x5091 <= 0;
      x5095 <= 0;
      x5099 <= 0;
      x5103 <= 0;
      x5107 <= 0;
      x5111 <= 0;
      x5115 <= 0;
      x5119 <= 0;
      x5123 <= 0;
      x5127 <= 0;
      x5131 <= 0;
      x5135 <= 0;
      x5139 <= 0;
      x5143 <= 0;
      x5147 <= 0;
      x5151 <= 0;
      x5155 <= 0;
      x5159 <= 0;
      x5163 <= 0;
      x5167 <= 0;
      x5171 <= 0;
      x5175 <= 0;
      x5181 <= 0;
      x5185 <= 0;
      x5189 <= 0;
      x5193 <= 0;
      x5197 <= 0;
      x5201 <= 0;
      x5205 <= 0;
      x5209 <= 0;
      x5213 <= 0;
      x5217 <= 0;
      x5221 <= 0;
      x5225 <= 0;
      x5229 <= 0;
      x5233 <= 0;
      x5237 <= 0;
      x5241 <= 0;
      x5245 <= 0;
      x5249 <= 0;
      x5253 <= 0;
      x5257 <= 0;
      x5261 <= 0;
      x5265 <= 0;
      x5269 <= 0;
      x5273 <= 0;
      x5277 <= 0;
      x5281 <= 0;
      x5285 <= 0;
      x5289 <= 0;
      x5293 <= 0;
      x5297 <= 0;
      x5301 <= 0;
      x5305 <= 0;
      x5311 <= 0;
      x5315 <= 0;
      x5319 <= 0;
      x5323 <= 0;
      x5327 <= 0;
      x5331 <= 0;
      x5335 <= 0;
      x5339 <= 0;
      x5343 <= 0;
      x5347 <= 0;
      x5351 <= 0;
      x5355 <= 0;
      x5359 <= 0;
      x5363 <= 0;
      x5367 <= 0;
      x5371 <= 0;
      x5375 <= 0;
      x5379 <= 0;
      x5383 <= 0;
      x5387 <= 0;
      x5391 <= 0;
      x5395 <= 0;
      x5399 <= 0;
      x5403 <= 0;
      x5407 <= 0;
      x5411 <= 0;
      x5415 <= 0;
      x5419 <= 0;
      x5423 <= 0;
      x5427 <= 0;
      x5431 <= 0;
      x5435 <= 0;
      x5442 <= 0;
      x5448 <= 0;
      x5453 <= 0;
      x5457 <= 0;
      x5461 <= 0;
      x5465 <= 0;
      x5469 <= 0;
      x5473 <= 0;
      x5477 <= 0;
      x5481 <= 0;
      x5485 <= 0;
      x5489 <= 0;
      x5493 <= 0;
      x5497 <= 0;
      x5501 <= 0;
      x5505 <= 0;
      x5509 <= 0;
      x5513 <= 0;
      x5517 <= 0;
      x5521 <= 0;
      x5525 <= 0;
      x5529 <= 0;
      x5533 <= 0;
      x5537 <= 0;
      x5541 <= 0;
      x5545 <= 0;
      x5549 <= 0;
      x5553 <= 0;
      x5557 <= 0;
      x5561 <= 0;
      x5565 <= 0;
      x5569 <= 0;
      x5575 <= 0;
      x5579 <= 0;
      x5583 <= 0;
      x5587 <= 0;
      x5591 <= 0;
      x5595 <= 0;
      x5599 <= 0;
      x5603 <= 0;
      x5607 <= 0;
      x5611 <= 0;
      x5615 <= 0;
      x5619 <= 0;
      x5623 <= 0;
      x5627 <= 0;
      x5631 <= 0;
      x5635 <= 0;
      x5639 <= 0;
      x5643 <= 0;
      x5647 <= 0;
      x5651 <= 0;
      x5655 <= 0;
      x5659 <= 0;
      x5663 <= 0;
      x5667 <= 0;
      x5671 <= 0;
      x5675 <= 0;
      x5679 <= 0;
      x5683 <= 0;
      x5687 <= 0;
      x5691 <= 0;
      x5695 <= 0;
      x5699 <= 0;
      x5705 <= 0;
      x5709 <= 0;
      x5713 <= 0;
      x5717 <= 0;
      x5721 <= 0;
      x5725 <= 0;
      x5729 <= 0;
      x5733 <= 0;
      x5737 <= 0;
      x5741 <= 0;
      x5745 <= 0;
      x5749 <= 0;
      x5753 <= 0;
      x5757 <= 0;
      x5761 <= 0;
      x5765 <= 0;
      x5769 <= 0;
      x5773 <= 0;
      x5777 <= 0;
      x5781 <= 0;
      x5785 <= 0;
      x5789 <= 0;
      x5793 <= 0;
      x5797 <= 0;
      x5801 <= 0;
      x5805 <= 0;
      x5809 <= 0;
      x5813 <= 0;
      x5817 <= 0;
      x5821 <= 0;
      x5825 <= 0;
      x5829 <= 0;
      x5835 <= 0;
      x5839 <= 0;
      x5843 <= 0;
      x5847 <= 0;
      x5851 <= 0;
      x5855 <= 0;
      x5859 <= 0;
      x5863 <= 0;
      x5867 <= 0;
      x5871 <= 0;
      x5875 <= 0;
      x5879 <= 0;
      x5883 <= 0;
      x5887 <= 0;
      x5891 <= 0;
      x5895 <= 0;
      x5899 <= 0;
      x5903 <= 0;
      x5907 <= 0;
      x5911 <= 0;
      x5915 <= 0;
      x5919 <= 0;
      x5923 <= 0;
      x5927 <= 0;
      x5931 <= 0;
      x5935 <= 0;
      x5939 <= 0;
      x5943 <= 0;
      x5947 <= 0;
      x5951 <= 0;
      x5955 <= 0;
      x5959 <= 0;
      x5965 <= 0;
      x5969 <= 0;
      x5973 <= 0;
      x5977 <= 0;
      x5981 <= 0;
      x5985 <= 0;
      x5989 <= 0;
      x5993 <= 0;
      x5997 <= 0;
      x6001 <= 0;
      x6005 <= 0;
      x6009 <= 0;
      x6013 <= 0;
      x6017 <= 0;
      x6021 <= 0;
      x6025 <= 0;
      x6029 <= 0;
      x6033 <= 0;
      x6037 <= 0;
      x6041 <= 0;
      x6045 <= 0;
      x6049 <= 0;
      x6053 <= 0;
      x6057 <= 0;
      x6061 <= 0;
      x6065 <= 0;
      x6069 <= 0;
      x6073 <= 0;
      x6077 <= 0;
      x6081 <= 0;
      x6085 <= 0;
      x6089 <= 0;
      x6095 <= 0;
      x6099 <= 0;
      x6103 <= 0;
      x6107 <= 0;
      x6111 <= 0;
      x6115 <= 0;
      x6119 <= 0;
      x6123 <= 0;
      x6127 <= 0;
      x6131 <= 0;
      x6135 <= 0;
      x6139 <= 0;
      x6143 <= 0;
      x6147 <= 0;
      x6151 <= 0;
      x6155 <= 0;
      x6159 <= 0;
      x6163 <= 0;
      x6167 <= 0;
      x6171 <= 0;
      x6175 <= 0;
      x6179 <= 0;
      x6183 <= 0;
      x6187 <= 0;
      x6191 <= 0;
      x6195 <= 0;
      x6199 <= 0;
      x6203 <= 0;
      x6207 <= 0;
      x6211 <= 0;
      x6215 <= 0;
      x6219 <= 0;
      x6225 <= 0;
      x6229 <= 0;
      x6233 <= 0;
      x6237 <= 0;
      x6241 <= 0;
      x6245 <= 0;
      x6249 <= 0;
      x6253 <= 0;
      x6257 <= 0;
      x6261 <= 0;
      x6265 <= 0;
      x6269 <= 0;
      x6273 <= 0;
      x6277 <= 0;
      x6281 <= 0;
      x6285 <= 0;
      x6289 <= 0;
      x6293 <= 0;
      x6297 <= 0;
      x6301 <= 0;
      x6305 <= 0;
      x6309 <= 0;
      x6313 <= 0;
      x6317 <= 0;
      x6321 <= 0;
      x6325 <= 0;
      x6329 <= 0;
      x6333 <= 0;
      x6337 <= 0;
      x6341 <= 0;
      x6345 <= 0;
      x6349 <= 0;
      x6355 <= 0;
      x6359 <= 0;
      x6363 <= 0;
      x6367 <= 0;
      x6371 <= 0;
      x6375 <= 0;
      x6379 <= 0;
      x6383 <= 0;
      x6387 <= 0;
      x6391 <= 0;
      x6395 <= 0;
      x6399 <= 0;
      x6403 <= 0;
      x6407 <= 0;
      x6411 <= 0;
      x6415 <= 0;
      x6419 <= 0;
      x6423 <= 0;
      x6427 <= 0;
      x6431 <= 0;
      x6435 <= 0;
      x6439 <= 0;
      x6443 <= 0;
      x6447 <= 0;
      x6451 <= 0;
      x6455 <= 0;
      x6459 <= 0;
      x6463 <= 0;
      x6467 <= 0;
      x6471 <= 0;
      x6475 <= 0;
      x6479 <= 0;
      x14598 <= 0;
      x14608 <= 0;
      x14618 <= 0;
      x14628 <= 0;
      x14638 <= 0;
      x14648 <= 0;
      x14658 <= 0;
      x14668 <= 0;
      x14767 <= 0;
      x14771 <= 0;
      x14775 <= 0;
      x14779 <= 0;
      x14783 <= 0;
      x14787 <= 0;
      x14793 <= 0;
      x14797 <= 0;
      x14801 <= 0;
      x14805 <= 0;
      x14809 <= 0;
      x14813 <= 0;
      x14819 <= 0;
      x14823 <= 0;
      x14827 <= 0;
      x14831 <= 0;
      x14835 <= 0;
      x14839 <= 0;
      x14845 <= 0;
      x14849 <= 0;
      x14853 <= 0;
      x14857 <= 0;
      x14861 <= 0;
      x14865 <= 0;
      x14871 <= 0;
      x14875 <= 0;
      x14879 <= 0;
      x14883 <= 0;
      x14887 <= 0;
      x14891 <= 0;
      x14897 <= 0;
      x14901 <= 0;
      x14905 <= 0;
      x14909 <= 0;
      x14913 <= 0;
      x14917 <= 0;
      x14923 <= 0;
      x14927 <= 0;
      x14931 <= 0;
      x14935 <= 0;
      x14939 <= 0;
      x14943 <= 0;
      x14949 <= 0;
      x14953 <= 0;
      x14957 <= 0;
      x14961 <= 0;
      x14965 <= 0;
      x14969 <= 0;
      x27755 <= 0;
      x27759 <= 0;
      x27763 <= 0;
      x27767 <= 0;
      x27771 <= 0;
      x27775 <= 0;
      x27779 <= 0;
      x27783 <= 0;
      x27787 <= 0;
      x27791 <= 0;
      x27795 <= 0;
      x27799 <= 0;
      x27803 <= 0;
      x27807 <= 0;
      x27811 <= 0;
      x27815 <= 0;
      x27819 <= 0;
      x27823 <= 0;
      x27827 <= 0;
      x27831 <= 0;
      x27835 <= 0;
      x27839 <= 0;
      x27843 <= 0;
      x27847 <= 0;
      x27851 <= 0;
      x27855 <= 0;
      x27859 <= 0;
      x27863 <= 0;
      x27867 <= 0;
      x27871 <= 0;
      x27875 <= 0;
      x27879 <= 0;
      x38722 <= 0;
      x38726 <= 0;
      x38730 <= 0;
      x38734 <= 0;
      x38738 <= 0;
      x38742 <= 0;
      x38746 <= 0;
      x38750 <= 0;
      x38754 <= 0;
      x38758 <= 0;
      x38762 <= 0;
      x38766 <= 0;
      x38770 <= 0;
      x38774 <= 0;
      x38778 <= 0;
      x38782 <= 0;
      x38786 <= 0;
      x38790 <= 0;
      x38794 <= 0;
      x38798 <= 0;
      x38802 <= 0;
      x38806 <= 0;
      x38810 <= 0;
      x38814 <= 0;
      x38818 <= 0;
      x38822 <= 0;
      x38826 <= 0;
      x38830 <= 0;
      x38834 <= 0;
      x38838 <= 0;
      x38842 <= 0;
      x38846 <= 0;
      x49689 <= 0;
      x49693 <= 0;
      x49697 <= 0;
      x49701 <= 0;
      x49705 <= 0;
      x49709 <= 0;
      x49713 <= 0;
      x49717 <= 0;
      x49721 <= 0;
      x49725 <= 0;
      x49729 <= 0;
      x49733 <= 0;
      x49737 <= 0;
      x49741 <= 0;
      x49745 <= 0;
      x49749 <= 0;
      x49753 <= 0;
      x49757 <= 0;
      x49761 <= 0;
      x49765 <= 0;
      x49769 <= 0;
      x49773 <= 0;
      x49777 <= 0;
      x49781 <= 0;
      x49785 <= 0;
      x49789 <= 0;
      x49793 <= 0;
      x49797 <= 0;
      x49801 <= 0;
      x49805 <= 0;
      x49809 <= 0;
      x49813 <= 0;
      x60656 <= 0;
      x60660 <= 0;
      x60664 <= 0;
      x60668 <= 0;
      x60672 <= 0;
      x60676 <= 0;
      x60680 <= 0;
      x60684 <= 0;
      x60688 <= 0;
      x60692 <= 0;
      x60696 <= 0;
      x60700 <= 0;
      x60704 <= 0;
      x60708 <= 0;
      x60712 <= 0;
      x60716 <= 0;
      x60720 <= 0;
      x60724 <= 0;
      x60728 <= 0;
      x60732 <= 0;
      x60736 <= 0;
      x60740 <= 0;
      x60744 <= 0;
      x60748 <= 0;
      x60752 <= 0;
      x60756 <= 0;
      x60760 <= 0;
      x60764 <= 0;
      x60768 <= 0;
      x60772 <= 0;
      x60776 <= 0;
      x60780 <= 0;
      x60784 <= 0;
      x60788 <= 0;
      x60792 <= 0;
      x60796 <= 0;
      x60800 <= 0;
      x60804 <= 0;
      x60808 <= 0;
      x60812 <= 0;
      x60816 <= 0;
      x60820 <= 0;
      x60824 <= 0;
      x60828 <= 0;
      x60832 <= 0;
      x60836 <= 0;
      x60840 <= 0;
      x60976 <= 0;
      x61105 <= 0;
      x61234 <= 0;
      x61363 <= 0;
      x61367 <= 0;
      x61371 <= 0;
      x61375 <= 0;
      x61379 <= 0;
      x61383 <= 0;
      x61387 <= 0;
      x61391 <= 0;
      x61395 <= 0;
      x61399 <= 0;
      x61403 <= 0;
      x61407 <= 0;
      x61411 <= 0;
      x61415 <= 0;
      x61419 <= 0;
      x61423 <= 0;
      x61981 <= 0;
      x61988 <= 0;
      x61995 <= 0;
      x62002 <= 0;
      x62009 <= 0;
      x62016 <= 0;
      x62023 <= 0;
      x62030 <= 0;
      x62037 <= 0;
      x62044 <= 0;
      x62051 <= 0;
      x62058 <= 0;
      x62065 <= 0;
      x62072 <= 0;
      x62079 <= 0;
      x62086 <= 0;
      x62093 <= 0;
      x62100 <= 0;
      x62107 <= 0;
      x62114 <= 0;
      x62121 <= 0;
      x62128 <= 0;
      x62135 <= 0;
      x62142 <= 0;
      x62149 <= 0;
      x62156 <= 0;
      x62163 <= 0;
      x62170 <= 0;
      x62177 <= 0;
      x62184 <= 0;
      x62191 <= 0;
      x62198 <= 0;
      x62205 <= 0;
      x62212 <= 0;
      x62219 <= 0;
      x62226 <= 0;
      x62233 <= 0;
      x62240 <= 0;
      x62247 <= 0;
      x62254 <= 0;
      x62261 <= 0;
      x62268 <= 0;
      x62275 <= 0;
      x62282 <= 0;
      x62289 <= 0;
      x62296 <= 0;
      x62303 <= 0;
      x62310 <= 0;
      x62317 <= 0;
      x62324 <= 0;
      x62331 <= 0;
      x62338 <= 0;
      x62345 <= 0;
      x62352 <= 0;
      x62359 <= 0;
      x62366 <= 0;
      x62373 <= 0;
      x62380 <= 0;
      x62387 <= 0;
      x62394 <= 0;
      x62401 <= 0;
      x62408 <= 0;
      x62415 <= 0;
      x62422 <= 0;
      x62429 <= 0;
      x62436 <= 0;
      x62443 <= 0;
      x62450 <= 0;
      x62457 <= 0;
      x62464 <= 0;
      x62471 <= 0;
      x62478 <= 0;
      x62485 <= 0;
      x62492 <= 0;
      x62499 <= 0;
      x62506 <= 0;
      x62513 <= 0;
      x62520 <= 0;
      x62527 <= 0;
      x62534 <= 0;
      x62541 <= 0;
      x62548 <= 0;
      x62555 <= 0;
      x62562 <= 0;
      x62569 <= 0;
      x62576 <= 0;
      x62583 <= 0;
      x62590 <= 0;
      x62597 <= 0;
      x62604 <= 0;
      x62611 <= 0;
      x62618 <= 0;
      x62625 <= 0;
      x62632 <= 0;
      x62639 <= 0;
      x62646 <= 0;
      x62653 <= 0;
      x62660 <= 0;
      x62667 <= 0;
      x62674 <= 0;
      x62681 <= 0;
      x62688 <= 0;
      x62695 <= 0;
      x62702 <= 0;
      x62709 <= 0;
      x62716 <= 0;
      x62723 <= 0;
      x62730 <= 0;
      x62737 <= 0;
      x62744 <= 0;
      x62751 <= 0;
      x62758 <= 0;
      x62765 <= 0;
      x62772 <= 0;
      x62779 <= 0;
      x62786 <= 0;
      x62793 <= 0;
      x62800 <= 0;
      x62807 <= 0;
      x62814 <= 0;
      x62821 <= 0;
      x62828 <= 0;
      x62835 <= 0;
      x62842 <= 0;
      x62849 <= 0;
      x62856 <= 0;
      x62863 <= 0;
      x62870 <= 0;
      x62873 <= 0;
      x62877 <= 0;
      x62881 <= 0;
      x62885 <= 0;
      x62889 <= 0;
      x62893 <= 0;
      x62897 <= 0;
      x62901 <= 0;
      x62905 <= 0;
      x62909 <= 0;
      x62913 <= 0;
      x62917 <= 0;
      x62921 <= 0;
      x62925 <= 0;
      x62929 <= 0;
      x63908 <= 0;
      x63909 <= 0;
      x63910 <= 0;
      x63911 <= 0;
      x63912 <= 0;
      x64640 <= 0;
      x64641 <= 0;
      x64642 <= 0;
      x64643 <= 0;
      x64644 <= 0;
      x65310 <= 0;
      x65311 <= 0;
      x65312 <= 0;
      x65313 <= 0;
      x65314 <= 0;
      x65980 <= 0;
      x65981 <= 0;
      x65982 <= 0;
      x65983 <= 0;
      x65984 <= 0;
      x66413 <= 0;
      x66417 <= 0;
      x66421 <= 0;
      x66425 <= 0;
      x66429 <= 0;
      x66433 <= 0;
      x66437 <= 0;
      x66441 <= 0;
      x66445 <= 0;
      x66449 <= 0;
      x66453 <= 0;
      x66457 <= 0;
      x66461 <= 0;
      x66465 <= 0;
      x66469 <= 0;
      x66894 <= 0;
      x66898 <= 0;
      x66902 <= 0;
      x66906 <= 0;
      x66910 <= 0;
      x66914 <= 0;
      x66918 <= 0;
      x66922 <= 0;
      x66926 <= 0;
      x66930 <= 0;
      x66934 <= 0;
      x66938 <= 0;
      x66942 <= 0;
      x66946 <= 0;
      x66950 <= 0;
      x66954 <= 0;
      x66958 <= 0;
      x66962 <= 0;
      x66966 <= 0;
      x66970 <= 0;
      x66974 <= 0;
      x66978 <= 0;
      x66982 <= 0;
      x66986 <= 0;
      x66990 <= 0;
      x66994 <= 0;
      x66998 <= 0;
      x67002 <= 0;
      x67006 <= 0;
      x67010 <= 0;
      x67014 <= 0;
      x67018 <= 0;
      x67022 <= 0;
      x67026 <= 0;
      x67030 <= 0;
      x67034 <= 0;
      x67038 <= 0;
      x67042 <= 0;
      x67046 <= 0;
      x67050 <= 0;
      x67054 <= 0;
      x67058 <= 0;
      x67062 <= 0;
      x67066 <= 0;
      x67070 <= 0;
      x67074 <= 0;
      x67078 <= 0;
      x67082 <= 0;
      x67086 <= 0;
      x67090 <= 0;
      x67094 <= 0;
      x67098 <= 0;
      x67102 <= 0;
      x67106 <= 0;
      x67110 <= 0;
      x67114 <= 0;
      x67118 <= 0;
      x67122 <= 0;
      x67126 <= 0;
      x67130 <= 0;
      x67134 <= 0;
      x67138 <= 0;
      x67142 <= 0;
      x67146 <= 0;
      x67150 <= 0;
      x67154 <= 0;
      x67158 <= 0;
      x67162 <= 0;
      x67166 <= 0;
      x67170 <= 0;
      x67174 <= 0;
      x67178 <= 0;
      x67182 <= 0;
      x67186 <= 0;
      x67190 <= 0;
      x67194 <= 0;
      x67198 <= 0;
      x67202 <= 0;
      x67206 <= 0;
      x67210 <= 0;
      x67214 <= 0;
      x67218 <= 0;
      x67222 <= 0;
      x67226 <= 0;
      x67230 <= 0;
      x67234 <= 0;
      x67238 <= 0;
      x67242 <= 0;
      x67246 <= 0;
      x67250 <= 0;
      x67254 <= 0;
      x67258 <= 0;
      x67262 <= 0;
      x67266 <= 0;
      x67270 <= 0;
      x67274 <= 0;
      x67278 <= 0;
      x67282 <= 0;
      x67286 <= 0;
      x67290 <= 0;
      x67294 <= 0;
      x67298 <= 0;
      x67302 <= 0;
      x67306 <= 0;
      x67310 <= 0;
      x67314 <= 0;
      x67318 <= 0;
      x67322 <= 0;
      x67326 <= 0;
      x67330 <= 0;
      x67334 <= 0;
      x67338 <= 0;
      x67342 <= 0;
      x67346 <= 0;
      x67350 <= 0;
      x67354 <= 0;
      x67358 <= 0;
      x67362 <= 0;
      x67366 <= 0;
      x67370 <= 0;
      x67374 <= 0;
      x67378 <= 0;
      x67382 <= 0;
      x67386 <= 0;
      x67390 <= 0;
      x67394 <= 0;
      x67398 <= 0;
      x67402 <= 0;
      x67405 <= 0;
      x67409 <= 0;
      x67413 <= 0;
      x67417 <= 0;
      x67421 <= 0;
      x67425 <= 0;
      x67429 <= 0;
      x67433 <= 0;
      x67437 <= 0;
      x67441 <= 0;
      x67445 <= 0;
      x67449 <= 0;
      x67453 <= 0;
      x67457 <= 0;
      x67461 <= 0;
      x67887 <= 0;
      x67891 <= 0;
      x67895 <= 0;
      x67899 <= 0;
      x67903 <= 0;
      x67907 <= 0;
      x67911 <= 0;
      x67915 <= 0;
      x67919 <= 0;
      x67923 <= 0;
      x67927 <= 0;
      x67931 <= 0;
      x67935 <= 0;
      x67939 <= 0;
      x67943 <= 0;
      x67947 <= 0;
      x67951 <= 0;
      x67955 <= 0;
      x67959 <= 0;
      x67963 <= 0;
      x67967 <= 0;
      x67971 <= 0;
      x67975 <= 0;
      x67979 <= 0;
      x67983 <= 0;
      x67987 <= 0;
      x67991 <= 0;
      x67995 <= 0;
      x67999 <= 0;
      x68003 <= 0;
      x68007 <= 0;
      x68011 <= 0;
      x68015 <= 0;
      x68019 <= 0;
      x68023 <= 0;
      x68027 <= 0;
      x68031 <= 0;
      x68035 <= 0;
      x68039 <= 0;
      x68043 <= 0;
      x68047 <= 0;
      x68051 <= 0;
      x68055 <= 0;
      x68059 <= 0;
      x68063 <= 0;
      x68067 <= 0;
      x68071 <= 0;
      x68075 <= 0;
      x68079 <= 0;
      x68083 <= 0;
      x68087 <= 0;
      x68091 <= 0;
      x68095 <= 0;
      x68099 <= 0;
      x68103 <= 0;
      x68107 <= 0;
      x68111 <= 0;
      x68115 <= 0;
      x68119 <= 0;
      x68123 <= 0;
      x68127 <= 0;
      x68131 <= 0;
      x68135 <= 0;
      x68139 <= 0;
      x68143 <= 0;
      x68147 <= 0;
      x68151 <= 0;
      x68155 <= 0;
      x68159 <= 0;
      x68163 <= 0;
      x68167 <= 0;
      x68171 <= 0;
      x68175 <= 0;
      x68179 <= 0;
      x68183 <= 0;
      x68187 <= 0;
      x68191 <= 0;
      x68195 <= 0;
      x68199 <= 0;
      x68203 <= 0;
      x68207 <= 0;
      x68211 <= 0;
      x68215 <= 0;
      x68219 <= 0;
      x68223 <= 0;
      x68227 <= 0;
      x68231 <= 0;
      x68235 <= 0;
      x68239 <= 0;
      x68243 <= 0;
      x68247 <= 0;
      x68251 <= 0;
      x68255 <= 0;
      x68259 <= 0;
      x68263 <= 0;
      x68267 <= 0;
      x68271 <= 0;
      x68275 <= 0;
      x68279 <= 0;
      x68283 <= 0;
      x68287 <= 0;
      x68291 <= 0;
      x68295 <= 0;
      x68299 <= 0;
      x68303 <= 0;
      x68307 <= 0;
      x68311 <= 0;
      x68315 <= 0;
      x68319 <= 0;
      x68323 <= 0;
      x68327 <= 0;
      x68331 <= 0;
      x68335 <= 0;
      x68339 <= 0;
      x68343 <= 0;
      x68347 <= 0;
      x68351 <= 0;
      x68355 <= 0;
      x68359 <= 0;
      x68363 <= 0;
      x68367 <= 0;
      x68371 <= 0;
      x68375 <= 0;
      x68379 <= 0;
      x68383 <= 0;
      x68387 <= 0;
      x68391 <= 0;
      x68395 <= 0;
      x68398 <= 0;
      x68402 <= 0;
      x68406 <= 0;
      x68410 <= 0;
      x68414 <= 0;
      x68418 <= 0;
      x68422 <= 0;
      x68426 <= 0;
      x68430 <= 0;
      x68434 <= 0;
      x68438 <= 0;
      x68442 <= 0;
      x68446 <= 0;
      x68450 <= 0;
      x68454 <= 0;
      x68618 <= 0;
      x68619 <= 0;
      x68620 <= 0;
      x68621 <= 0;
      x68622 <= 0;
      x68623 <= 0;
      x71147 <= 0;
      x71152 <= 0;
      x71157 <= 0;
      x71162 <= 0;
      x71167 <= 0;
      x71172 <= 0;
      x71177 <= 0;
      x71182 <= 0;
      x71185 <= 0;
      x71188 <= 0;
      x71191 <= 0;
      x71194 <= 0;
      x71197 <= 0;
      x71202 <= 0;
      x71205 <= 0;
      x71210 <= 0;
      x71215 <= 0;
      x71220 <= 0;
      x71225 <= 0;
      x71230 <= 0;
      x71235 <= 0;
      x71240 <= 0;
      x71245 <= 0;
      x71250 <= 0;
      x71255 <= 0;
      x71260 <= 0;
      x71265 <= 0;
      x71270 <= 0;
      x71275 <= 0;
      x71277 <= 0;
      x71279 <= 0;
      x71284 <= 0;
      x71289 <= 0;
      x71294 <= 0;
      x71299 <= 0;
      x71304 <= 0;
      x71309 <= 0;
      x71314 <= 0;
      x71319 <= 0;
      x71324 <= 0;
      x71329 <= 0;
      x71334 <= 0;
      x71339 <= 0;
      x71344 <= 0;
      x71349 <= 0;
      x71354 <= 0;
      x71359 <= 0;
      x71364 <= 0;
      x71369 <= 0;
      x71374 <= 0;
      x71379 <= 0;
      x71384 <= 0;
      x71389 <= 0;
      x71394 <= 0;
      x71399 <= 0;
      x71404 <= 0;
      x71409 <= 0;
      x71414 <= 0;
      x71419 <= 0;
      x71424 <= 0;
      x71429 <= 0;
      x71434 <= 0;
      x71439 <= 0;
      x71444 <= 0;
      x71449 <= 0;
      x71454 <= 0;
      x71459 <= 0;
      x71464 <= 0;
      x71469 <= 0;
      x71474 <= 0;
      x71479 <= 0;
      x71482 <= 0;
      x71485 <= 0;
      x71490 <= 0;
      x71495 <= 0;
      x71500 <= 0;
      x71505 <= 0;
      x71510 <= 0;
      x71515 <= 0;
      x71520 <= 0;
      x71525 <= 0;
      x71530 <= 0;
      x71535 <= 0;
      x71540 <= 0;
      x71545 <= 0;
      x71550 <= 0;
      x71555 <= 0;
      x71560 <= 0;
      x71565 <= 0;
      x71570 <= 0;
      x71575 <= 0;
      x71580 <= 0;
      x71585 <= 0;
      x71590 <= 0;
      x71595 <= 0;
      x71600 <= 0;
      x71605 <= 0;
      x71610 <= 0;
      x71615 <= 0;
      x71620 <= 0;
      x71625 <= 0;
      x71630 <= 0;
      x71635 <= 0;
      x71642 <= 0;
      x71647 <= 0;
      x71652 <= 0;
      x71657 <= 0;
      x71662 <= 0;
      x71667 <= 0;
      x71672 <= 0;
      x71677 <= 0;
      x71682 <= 0;
      x71687 <= 0;
      x71692 <= 0;
      x71697 <= 0;
      x71702 <= 0;
      x71707 <= 0;
      x71712 <= 0;
      x71717 <= 0;
      x71722 <= 0;
      x71727 <= 0;
      x71732 <= 0;
      x71737 <= 0;
      x71742 <= 0;
      x71747 <= 0;
      x71752 <= 0;
      x71757 <= 0;
      x71762 <= 0;
      x71767 <= 0;
      x71772 <= 0;
      x71777 <= 0;
      x71782 <= 0;
      x71787 <= 0;
      x71792 <= 0;
      x71797 <= 0;
      x71802 <= 0;
      x71807 <= 0;
      x71812 <= 0;
      x71817 <= 0;
      x71822 <= 0;
      x71827 <= 0;
      x71832 <= 0;
      x71837 <= 0;
      x71842 <= 0;
      x71847 <= 0;
      x71852 <= 0;
      x71857 <= 0;
      x71862 <= 0;
      x71867 <= 0;
      x71872 <= 0;
      x71877 <= 0;
      x71882 <= 0;
      x71887 <= 0;
      x71892 <= 0;
      x71897 <= 0;
      x71902 <= 0;
      x71907 <= 0;
      x71910 <= 0;
      x71913 <= 0;
      x71916 <= 0;
      x71919 <= 0;
      x71922 <= 0;
      x71925 <= 0;
      x71928 <= 0;
      x71931 <= 0;
      x71934 <= 0;
      x71937 <= 0;
      x71942 <= 0;
      x71947 <= 0;
      x71952 <= 0;
      x71957 <= 0;
      x71962 <= 0;
      x71967 <= 0;
      x71972 <= 0;
      x71977 <= 0;
      x71982 <= 0;
      x71987 <= 0;
      x71992 <= 0;
      x71997 <= 0;
      x72002 <= 0;
      x72007 <= 0;
      x72012 <= 0;
      x72017 <= 0;
      x72022 <= 0;
      x72027 <= 0;
      x72032 <= 0;
      x72037 <= 0;
      x72042 <= 0;
      x72047 <= 0;
      x72052 <= 0;
      x72057 <= 0;
      x72062 <= 0;
      x72067 <= 0;
      x72072 <= 0;
      x72077 <= 0;
      x72082 <= 0;
      x72087 <= 0;
      x72092 <= 0;
      x72097 <= 0;
      x72102 <= 0;
      x72107 <= 0;
      x72112 <= 0;
      x72117 <= 0;
      x72122 <= 0;
      x72127 <= 0;
      x72132 <= 0;
      x72137 <= 0;
      x72142 <= 0;
      x72147 <= 0;
      x72152 <= 0;
      x72157 <= 0;
      x72162 <= 0;
      x72167 <= 0;
      x72172 <= 0;
      x72177 <= 0;
      x72182 <= 0;
      x72187 <= 0;
      x72192 <= 0;
      x72197 <= 0;
      x72202 <= 0;
      x72207 <= 0;
      x72212 <= 0;
      x72217 <= 0;
      x72222 <= 0;
      x72227 <= 0;
      x72232 <= 0;
      x72237 <= 0;
      x72242 <= 0;
      x72247 <= 0;
      x72252 <= 0;
      x72257 <= 0;
      x72262 <= 0;
      x72267 <= 0;
      x72272 <= 0;
      x72277 <= 0;
      x72282 <= 0;
      x72287 <= 0;
      x72292 <= 0;
      x72297 <= 0;
      x72302 <= 0;
      x72307 <= 0;
      x72312 <= 0;
      x72317 <= 0;
      x72322 <= 0;
      x72327 <= 0;
      x72332 <= 0;
      x72337 <= 0;
      x72342 <= 0;
      x72347 <= 0;
      x72352 <= 0;
      x72357 <= 0;
      x72362 <= 0;
      x72367 <= 0;
      x72372 <= 0;
      x72377 <= 0;
      x72382 <= 0;
      x72387 <= 0;
      x72392 <= 0;
      x72397 <= 0;
      x72402 <= 0;
      x72407 <= 0;
      x72412 <= 0;
      x72417 <= 0;
      x72422 <= 0;
      x72427 <= 0;
      x72432 <= 0;
      x72437 <= 0;
      x72442 <= 0;
      x72447 <= 0;
      x72452 <= 0;
      x72457 <= 0;
      x72462 <= 0;
      x72467 <= 0;
      x72472 <= 0;
      x72477 <= 0;
      x72482 <= 0;
      x72487 <= 0;
      x72492 <= 0;
      x72497 <= 0;
      x72502 <= 0;
      x72507 <= 0;
      x72512 <= 0;
      x72517 <= 0;
      x72522 <= 0;
      x72527 <= 0;
      x72532 <= 0;
      x72537 <= 0;
      x72542 <= 0;
      x72547 <= 0;
      x72552 <= 0;
      x72557 <= 0;
      x72562 <= 0;
      x72567 <= 0;
      x72572 <= 0;
      x72577 <= 0;
      x72582 <= 0;
      x72587 <= 0;
      x72592 <= 0;
      x72597 <= 0;
      x72602 <= 0;
      x72607 <= 0;
      x72612 <= 0;
      x72617 <= 0;
      x72622 <= 0;
      x72627 <= 0;
      x72632 <= 0;
      x72637 <= 0;
      x72642 <= 0;
      x72647 <= 0;
      x72652 <= 0;
      x72657 <= 0;
      x72662 <= 0;
      x72667 <= 0;
      x72672 <= 0;
      x72677 <= 0;
      x72682 <= 0;
      x72687 <= 0;
      x72692 <= 0;
      x72697 <= 0;
      x72702 <= 0;
      x72707 <= 0;
      x72712 <= 0;
      x72717 <= 0;
      x72722 <= 0;
      x72727 <= 0;
      x72732 <= 0;
      x72737 <= 0;
      x72742 <= 0;
      x72747 <= 0;
      x72752 <= 0;
      x72757 <= 0;
      x72762 <= 0;
      x72767 <= 0;
      x72772 <= 0;
      x72777 <= 0;
      x72782 <= 0;
      x72787 <= 0;
      x72792 <= 0;
      x72797 <= 0;
      x72802 <= 0;
      x72807 <= 0;
      x72812 <= 0;
      x72817 <= 0;
      x72822 <= 0;
      x72827 <= 0;
      x72832 <= 0;
      x72837 <= 0;
      x72842 <= 0;
      x72847 <= 0;
      x72852 <= 0;
      x72857 <= 0;
      x72862 <= 0;
      x72867 <= 0;
      x72872 <= 0;
      x72877 <= 0;
      x72882 <= 0;
      x72887 <= 0;
      x72892 <= 0;
      x72897 <= 0;
      x72902 <= 0;
      x72907 <= 0;
      x72912 <= 0;
      x72917 <= 0;
      x72922 <= 0;
      x72927 <= 0;
      x72932 <= 0;
      x72937 <= 0;
      x72942 <= 0;
      x72947 <= 0;
      x72952 <= 0;
      x72957 <= 0;
      x72962 <= 0;
      x72967 <= 0;
      x72972 <= 0;
      x72977 <= 0;
      x72982 <= 0;
      x72987 <= 0;
      x72992 <= 0;
      x72997 <= 0;
      x73002 <= 0;
      x73007 <= 0;
      x73012 <= 0;
      x73017 <= 0;
      x73022 <= 0;
      x73027 <= 0;
      x73032 <= 0;
      x73037 <= 0;
      x73042 <= 0;
      x73047 <= 0;
      x73052 <= 0;
      x73057 <= 0;
      x73062 <= 0;
      x73067 <= 0;
      x73072 <= 0;
      x73077 <= 0;
      x73082 <= 0;
      x73087 <= 0;
      x73092 <= 0;
      x73097 <= 0;
      x73102 <= 0;
      x73107 <= 0;
      x73112 <= 0;
      x73117 <= 0;
      x73122 <= 0;
      x73127 <= 0;
      x73132 <= 0;
      x73137 <= 0;
      x73142 <= 0;
      x73147 <= 0;
      x73152 <= 0;
      x73157 <= 0;
      x73162 <= 0;
      x73167 <= 0;
      x73172 <= 0;
      x73177 <= 0;
      x73182 <= 0;
      x73187 <= 0;
      x73192 <= 0;
      x73197 <= 0;
      x73202 <= 0;
      x73207 <= 0;
      x73212 <= 0;
      x73217 <= 0;
      x73222 <= 0;
      x73227 <= 0;
      x73232 <= 0;
      x73237 <= 0;
      x73242 <= 0;
      x73247 <= 0;
      x73252 <= 0;
      x73257 <= 0;
      x73262 <= 0;
      x73267 <= 0;
      x73272 <= 0;
      x73277 <= 0;
      x73282 <= 0;
      x73287 <= 0;
      x73292 <= 0;
      x73297 <= 0;
      x73302 <= 0;
      x73307 <= 0;
      x73312 <= 0;
      x73317 <= 0;
      x73322 <= 0;
      x73327 <= 0;
      x73332 <= 0;
      x73337 <= 0;
      x73342 <= 0;
      x73347 <= 0;
      x73352 <= 0;
      x73357 <= 0;
      x73362 <= 0;
      x73367 <= 0;
      x73372 <= 0;
      x73377 <= 0;
      x73382 <= 0;
      x73387 <= 0;
      x73392 <= 0;
      x73397 <= 0;
      x73402 <= 0;
      x73407 <= 0;
      x73412 <= 0;
      x73417 <= 0;
      x73422 <= 0;
      x73427 <= 0;
      x73432 <= 0;
      x73437 <= 0;
      x73442 <= 0;
      x73447 <= 0;
      x73452 <= 0;
      x73457 <= 0;
      x73462 <= 0;
      x73467 <= 0;
      x73472 <= 0;
      x73477 <= 0;
      x73482 <= 0;
      x73487 <= 0;
      x73492 <= 0;
      x73497 <= 0;
      x73502 <= 0;
      x73507 <= 0;
      x73512 <= 0;
      x73517 <= 0;
      x73522 <= 0;
      x73527 <= 0;
      x73532 <= 0;
      x73537 <= 0;
      x73542 <= 0;
      x73547 <= 0;
      x73552 <= 0;
      x73557 <= 0;
      x73562 <= 0;
      x73567 <= 0;
      x73572 <= 0;
      x73577 <= 0;
      x73582 <= 0;
      x73587 <= 0;
      x73592 <= 0;
      x73597 <= 0;
      x73602 <= 0;
      x73607 <= 0;
      x73612 <= 0;
      x73617 <= 0;
      x73622 <= 0;
      x73627 <= 0;
      x73632 <= 0;
      x73637 <= 0;
      x73642 <= 0;
      x73647 <= 0;
      x73652 <= 0;
      x73657 <= 0;
      x73662 <= 0;
      x73667 <= 0;
      x73672 <= 0;
      x73677 <= 0;
      x73682 <= 0;
      x73687 <= 0;
      x73692 <= 0;
      x73697 <= 0;
      x73702 <= 0;
      x73707 <= 0;
      x73712 <= 0;
      x73717 <= 0;
      x73722 <= 0;
      x73727 <= 0;
      x73732 <= 0;
      x73737 <= 0;
      x73742 <= 0;
      x73747 <= 0;
      x73752 <= 0;
      x73757 <= 0;
      x73762 <= 0;
      x73767 <= 0;
      x73772 <= 0;
      x73777 <= 0;
      x73782 <= 0;
      x73787 <= 0;
      x73792 <= 0;
      x73797 <= 0;
      x73802 <= 0;
      x73807 <= 0;
      x73812 <= 0;
      x73817 <= 0;
      x73822 <= 0;
      x73827 <= 0;
      x73832 <= 0;
      x73837 <= 0;
      x73842 <= 0;
      x73847 <= 0;
      x73852 <= 0;
      x73857 <= 0;
      x73862 <= 0;
      x73867 <= 0;
      x73872 <= 0;
      x73877 <= 0;
      x73882 <= 0;
      x73887 <= 0;
      x73892 <= 0;
      x73897 <= 0;
      x73902 <= 0;
      x73907 <= 0;
      x73912 <= 0;
      x73917 <= 0;
      x73922 <= 0;
      x73927 <= 0;
      x73932 <= 0;
      x73937 <= 0;
      x73942 <= 0;
      x73947 <= 0;
      x73952 <= 0;
      x73957 <= 0;
      x73962 <= 0;
      x73967 <= 0;
      x73972 <= 0;
      x73977 <= 0;
      x73982 <= 0;
      x73987 <= 0;
      x73992 <= 0;
      x73997 <= 0;
      x74002 <= 0;
      x74005 <= 0;
      x74008 <= 0;
      x74011 <= 0;
      x74014 <= 0;
      x74017 <= 0;
      x74020 <= 0;
      x74023 <= 0;
      x74026 <= 0;
      x74029 <= 0;
      x74032 <= 0;
      x74035 <= 0;
      x74038 <= 0;
      x74041 <= 0;
      x74044 <= 0;
      x74047 <= 0;
      x74050 <= 0;
      x74053 <= 0;
      x74056 <= 0;
      x74059 <= 0;
      x74062 <= 0;
      x74065 <= 0;
      x74068 <= 0;
      x74071 <= 0;
      x74074 <= 0;
      x74077 <= 0;
      x74080 <= 0;
      x74083 <= 0;
      x74086 <= 0;
      x74089 <= 0;
      x74092 <= 0;
      x74095 <= 0;
      x74098 <= 0;
      x74101 <= 0;
      x74104 <= 0;
      x74107 <= 0;
      x74110 <= 0;
      x74113 <= 0;
      x74116 <= 0;
      x74119 <= 0;
      x74122 <= 0;
      x74125 <= 0;
      x74128 <= 0;
      x74131 <= 0;
      x74134 <= 0;
      x74137 <= 0;
      x74140 <= 0;
      x74143 <= 0;
      x74146 <= 0;
      x74149 <= 0;
      x74152 <= 0;
      x74155 <= 0;
      x74158 <= 0;
      x74161 <= 0;
      x74164 <= 0;
      x74167 <= 0;
      x74170 <= 0;
      x74173 <= 0;
      x74176 <= 0;
      x74179 <= 0;
      x74182 <= 0;
      x74185 <= 0;
      x74188 <= 0;
      x74191 <= 0;
      x74194 <= 0;
      x74197 <= 0;
      x74200 <= 0;
      x74203 <= 0;
      x74206 <= 0;
      x74209 <= 0;
      x74212 <= 0;
      x74215 <= 0;
      x74218 <= 0;
      x74221 <= 0;
      x74224 <= 0;
      x74227 <= 0;
      x74230 <= 0;
      x74233 <= 0;
      x74236 <= 0;
      x74239 <= 0;
      x74242 <= 0;
      x74245 <= 0;
      x74248 <= 0;
      x74251 <= 0;
      x74254 <= 0;
      x74257 <= 0;
      x74260 <= 0;
      x74263 <= 0;
      x74266 <= 0;
      x74269 <= 0;
      x74272 <= 0;
      x74275 <= 0;
      x74278 <= 0;
      x74281 <= 0;
      x74284 <= 0;
      x74287 <= 0;
      x74290 <= 0;
      x74293 <= 0;
      x74296 <= 0;
      x74299 <= 0;
      x74302 <= 0;
      x74305 <= 0;
      x74308 <= 0;
      x74311 <= 0;
      x74314 <= 0;
      x74317 <= 0;
      x74320 <= 0;
      x74323 <= 0;
      x74326 <= 0;
      x74329 <= 0;
      x74332 <= 0;
      x74335 <= 0;
      x74338 <= 0;
      x74341 <= 0;
      x74344 <= 0;
      x74347 <= 0;
      x74350 <= 0;
      x74353 <= 0;
      x74356 <= 0;
      x74359 <= 0;
      x74362 <= 0;
      x74365 <= 0;
      x74368 <= 0;
      x74371 <= 0;
      x74374 <= 0;
      x74377 <= 0;
      x74380 <= 0;
      x74383 <= 0;
      x74386 <= 0;
      x74389 <= 0;
      x74392 <= 0;
      x74395 <= 0;
      x74398 <= 0;
      x74401 <= 0;
      x74404 <= 0;
      x74407 <= 0;
      x74410 <= 0;
      x74413 <= 0;
      x74416 <= 0;
      x74419 <= 0;
      x74422 <= 0;
      x74425 <= 0;
      x74428 <= 0;
      x74431 <= 0;
      x74434 <= 0;
      x74437 <= 0;
      x74440 <= 0;
      x74443 <= 0;
      x74446 <= 0;
      x74449 <= 0;
      x74452 <= 0;
      x74455 <= 0;
      x74458 <= 0;
      x74461 <= 0;
      x74464 <= 0;
      x74467 <= 0;
      x74470 <= 0;
      x74473 <= 0;
      x74476 <= 0;
      x74479 <= 0;
      x74482 <= 0;
      x74485 <= 0;
      x74488 <= 0;
      x74491 <= 0;
      x74494 <= 0;
      x74497 <= 0;
      x74500 <= 0;
      x74503 <= 0;
      x74506 <= 0;
      x74509 <= 0;
      x74512 <= 0;
      x74515 <= 0;
      x74518 <= 0;
      x74521 <= 0;
      x74524 <= 0;
      x74527 <= 0;
      x74530 <= 0;
      x74533 <= 0;
      x74536 <= 0;
      x74539 <= 0;
      x74542 <= 0;
      x74545 <= 0;
      x74548 <= 0;
      x74551 <= 0;
      x74554 <= 0;
      x74557 <= 0;
      x74560 <= 0;
      x74563 <= 0;
      x74566 <= 0;
      x74569 <= 0;
      x74572 <= 0;
      x74575 <= 0;
      x74578 <= 0;
      x74581 <= 0;
      x74584 <= 0;
      x74587 <= 0;
      x74590 <= 0;
      x74593 <= 0;
      x74596 <= 0;
      x74599 <= 0;
      x74602 <= 0;
      x74605 <= 0;
      x74608 <= 0;
      x74611 <= 0;
      x74614 <= 0;
      x74617 <= 0;
      x74620 <= 0;
      x74623 <= 0;
      x74626 <= 0;
      x74629 <= 0;
      x74632 <= 0;
      x74635 <= 0;
      x74638 <= 0;
      x74641 <= 0;
      x74644 <= 0;
      x74647 <= 0;
      x74650 <= 0;
      x74653 <= 0;
      x74656 <= 0;
      x74659 <= 0;
      x74662 <= 0;
      x74665 <= 0;
      x74668 <= 0;
      x74671 <= 0;
      x74674 <= 0;
      x74677 <= 0;
      x74680 <= 0;
      x74683 <= 0;
      x74686 <= 0;
      x74689 <= 0;
      x74692 <= 0;
      x74695 <= 0;
      x74698 <= 0;
      x74701 <= 0;
      x74704 <= 0;
      x74707 <= 0;
      x74710 <= 0;
      x74713 <= 0;
      x74716 <= 0;
      x74719 <= 0;
      x74722 <= 0;
      x74725 <= 0;
      x74728 <= 0;
      x74731 <= 0;
      x74734 <= 0;
      x74737 <= 0;
      x74740 <= 0;
      x74743 <= 0;
      x74746 <= 0;
      x74749 <= 0;
      x74752 <= 0;
      x74755 <= 0;
      x74758 <= 0;
      x74761 <= 0;
      x74764 <= 0;
      x74767 <= 0;
      x74770 <= 0;
      x74773 <= 0;
      x74776 <= 0;
      x74779 <= 0;
      x74782 <= 0;
      x74785 <= 0;
      x74788 <= 0;
      x74791 <= 0;
      x74794 <= 0;
      x74797 <= 0;
      x74800 <= 0;
      x74803 <= 0;
      x74806 <= 0;
      x74809 <= 0;
      x74812 <= 0;
      x74815 <= 0;
      x74818 <= 0;
      x74821 <= 0;
      x74824 <= 0;
      x74827 <= 0;
      x74830 <= 0;
      x74833 <= 0;
      x74836 <= 0;
      x74839 <= 0;
      x74842 <= 0;
      x74845 <= 0;
      x74848 <= 0;
      x74851 <= 0;
      x74854 <= 0;
      x74857 <= 0;
      x74860 <= 0;
      x74863 <= 0;
      x74866 <= 0;
      x74869 <= 0;
      x74872 <= 0;
      x74875 <= 0;
      x74878 <= 0;
      x74881 <= 0;
      x74884 <= 0;
      x74887 <= 0;
      x74890 <= 0;
      x74893 <= 0;
      x74896 <= 0;
      x74899 <= 0;
      x74902 <= 0;
      x74905 <= 0;
      x74908 <= 0;
      x74911 <= 0;
      x74914 <= 0;
      x74917 <= 0;
      x74920 <= 0;
      x74923 <= 0;
      x74926 <= 0;
      x74929 <= 0;
      x74932 <= 0;
      x74935 <= 0;
      x74938 <= 0;
      x74941 <= 0;
      x74944 <= 0;
      x74947 <= 0;
      x74950 <= 0;
      x74953 <= 0;
      x74956 <= 0;
      x74959 <= 0;
      x74962 <= 0;
      x74965 <= 0;
      x74968 <= 0;
      x74971 <= 0;
      x74974 <= 0;
      x74977 <= 0;
      x74980 <= 0;
      x74983 <= 0;
      x74986 <= 0;
      x74989 <= 0;
      x74992 <= 0;
      x74995 <= 0;
      x74998 <= 0;
      x75001 <= 0;
      x75004 <= 0;
      x75007 <= 0;
      x75010 <= 0;
      x75013 <= 0;
      x75016 <= 0;
      x75019 <= 0;
      x75022 <= 0;
      x75025 <= 0;
      x75028 <= 0;
      x75031 <= 0;
      x75034 <= 0;
      x75037 <= 0;
      x75040 <= 0;
      x75043 <= 0;
      x75046 <= 0;
      x75049 <= 0;
      x75052 <= 0;
      x75055 <= 0;
      x75058 <= 0;
      x75061 <= 0;
      x75064 <= 0;
      x75067 <= 0;
      x75070 <= 0;
      x75073 <= 0;
      x75076 <= 0;
      x75079 <= 0;
      x75082 <= 0;
      x75085 <= 0;
      x75088 <= 0;
      x75091 <= 0;
      x75094 <= 0;
      x75097 <= 0;
      x75100 <= 0;
      x75103 <= 0;
      x75106 <= 0;
      x75109 <= 0;
      x75112 <= 0;
      x75115 <= 0;
      x75118 <= 0;
      x75121 <= 0;
      x75124 <= 0;
      x75127 <= 0;
      x75130 <= 0;
      x75133 <= 0;
      x75136 <= 0;
      x75139 <= 0;
      x75142 <= 0;
      x75145 <= 0;
      x75148 <= 0;
      x75151 <= 0;
      x75154 <= 0;
      x75157 <= 0;
      x75160 <= 0;
      x75163 <= 0;
      x75166 <= 0;
      x75169 <= 0;
      x75172 <= 0;
      x75175 <= 0;
      x75178 <= 0;
      x75181 <= 0;
      x75184 <= 0;
      x75187 <= 0;
      x75190 <= 0;
      x75193 <= 0;
      x75196 <= 0;
      x75199 <= 0;
      x75202 <= 0;
      x75205 <= 0;
      x75208 <= 0;
      x75211 <= 0;
      x75214 <= 0;
      x75217 <= 0;
      x75220 <= 0;
      x75223 <= 0;
      x75226 <= 0;
      x75229 <= 0;
      x75232 <= 0;
      x75235 <= 0;
      x75238 <= 0;
      x75241 <= 0;
      x75244 <= 0;
      x75247 <= 0;
      x75250 <= 0;
      x75253 <= 0;
      x75256 <= 0;
      x75259 <= 0;
      x75262 <= 0;
      x75265 <= 0;
      x75268 <= 0;
      x75271 <= 0;
      x75274 <= 0;
      x75277 <= 0;
      x75280 <= 0;
      x75283 <= 0;
      x75286 <= 0;
      x75289 <= 0;
      x75292 <= 0;
      x75295 <= 0;
      x75298 <= 0;
      x75301 <= 0;
      x75304 <= 0;
      x75307 <= 0;
      x75310 <= 0;
      x75313 <= 0;
      x75316 <= 0;
      x75319 <= 0;
      x75322 <= 0;
      x75325 <= 0;
      x75328 <= 0;
      x75331 <= 0;
      x75334 <= 0;
      x75337 <= 0;
      x75340 <= 0;
      x75343 <= 0;
      x75346 <= 0;
      x75349 <= 0;
      x75352 <= 0;
      x75355 <= 0;
      x75358 <= 0;
      x75361 <= 0;
      x75364 <= 0;
      x75367 <= 0;
      x75370 <= 0;
      x75373 <= 0;
      x75376 <= 0;
      x75379 <= 0;
      x75382 <= 0;
      x75385 <= 0;
      x75388 <= 0;
      x75391 <= 0;
      x75394 <= 0;
      x75397 <= 0;
      x75400 <= 0;
      x75403 <= 0;
      x75406 <= 0;
      x75409 <= 0;
      x75412 <= 0;
      x75415 <= 0;
      x75418 <= 0;
      x75421 <= 0;
      x75424 <= 0;
      x75427 <= 0;
      x75430 <= 0;
      x75433 <= 0;
      x75436 <= 0;
      x75439 <= 0;
      x75442 <= 0;
      x75445 <= 0;
      x75448 <= 0;
      x75451 <= 0;
      x75454 <= 0;
      x75457 <= 0;
      x75460 <= 0;
      x75463 <= 0;
      x75466 <= 0;
      x75469 <= 0;
      x75472 <= 0;
      x75475 <= 0;
      x75478 <= 0;
      x75481 <= 0;
      x75484 <= 0;
      x75487 <= 0;
      x75490 <= 0;
      x75493 <= 0;
      x75496 <= 0;
      x75499 <= 0;
      x75502 <= 0;
      x75505 <= 0;
      x75508 <= 0;
      x75511 <= 0;
      x75514 <= 0;
      x75517 <= 0;
      x75520 <= 0;
      x75523 <= 0;
      x75526 <= 0;
      x75529 <= 0;
      x75532 <= 0;
      x75535 <= 0;
      x75538 <= 0;
      x75541 <= 0;
      x75544 <= 0;
      x75547 <= 0;
      x75550 <= 0;
      x75553 <= 0;
      x75556 <= 0;
      x75559 <= 0;
      x75562 <= 0;
      x75565 <= 0;
      x75568 <= 0;
      x75571 <= 0;
      x75574 <= 0;
      x75577 <= 0;
      x75580 <= 0;
      x75583 <= 0;
      x75586 <= 0;
      x75589 <= 0;
      x75592 <= 0;
      x75595 <= 0;
      x75598 <= 0;
      x75601 <= 0;
      x75604 <= 0;
      x75607 <= 0;
      x75610 <= 0;
      x75613 <= 0;
      x75616 <= 0;
      x75619 <= 0;
      x75622 <= 0;
      x75625 <= 0;
      x75628 <= 0;
      x75631 <= 0;
      x75634 <= 0;
      x75637 <= 0;
      x75640 <= 0;
      x75643 <= 0;
      x75646 <= 0;
      x75649 <= 0;
      x75652 <= 0;
      x75655 <= 0;
      x75658 <= 0;
      x75661 <= 0;
      x75664 <= 0;
      x75667 <= 0;
      x75670 <= 0;
      x75673 <= 0;
      x75676 <= 0;
      x75679 <= 0;
      x75682 <= 0;
      x75685 <= 0;
      x75688 <= 0;
      x75691 <= 0;
      x75694 <= 0;
      x75697 <= 0;
      x75700 <= 0;
      x75703 <= 0;
      x75706 <= 0;
      x75709 <= 0;
      x75712 <= 0;
      x75715 <= 0;
      x75718 <= 0;
      x75721 <= 0;
      x75724 <= 0;
      x75727 <= 0;
      x75730 <= 0;
      x75733 <= 0;
      x75736 <= 0;
      x75739 <= 0;
      x75742 <= 0;
      x75745 <= 0;
      x75748 <= 0;
      x75751 <= 0;
      x75754 <= 0;
      x75757 <= 0;
      x75760 <= 0;
      x75763 <= 0;
      x75766 <= 0;
      x75769 <= 0;
      x75772 <= 0;
      x75775 <= 0;
      x75778 <= 0;
      x75781 <= 0;
      x75784 <= 0;
      x75787 <= 0;
      x75790 <= 0;
      x75793 <= 0;
      x75796 <= 0;
      x75799 <= 0;
      x75802 <= 0;
      x75805 <= 0;
      x75808 <= 0;
      x75811 <= 0;
      x75814 <= 0;
      x75817 <= 0;
      x75820 <= 0;
      x75823 <= 0;
      x75826 <= 0;
      x75829 <= 0;
      x75832 <= 0;
      x75835 <= 0;
      x75838 <= 0;
      x75841 <= 0;
      x75844 <= 0;
      x75847 <= 0;
      x75850 <= 0;
      x75853 <= 0;
      x75856 <= 0;
      x75859 <= 0;
      x75862 <= 0;
      x75865 <= 0;
      x75868 <= 0;
      x75871 <= 0;
      x75874 <= 0;
      x75877 <= 0;
      x75880 <= 0;
      x75883 <= 0;
      x75886 <= 0;
      x75889 <= 0;
      x75892 <= 0;
      x75895 <= 0;
      x75898 <= 0;
      x75901 <= 0;
      x75904 <= 0;
      x75907 <= 0;
      x75910 <= 0;
      x75913 <= 0;
      x75916 <= 0;
      x75919 <= 0;
      x75922 <= 0;
      x75925 <= 0;
      x75928 <= 0;
      x75931 <= 0;
      x75934 <= 0;
      x75937 <= 0;
      x75940 <= 0;
      x75943 <= 0;
      x75946 <= 0;
      x75949 <= 0;
      x75952 <= 0;
      x75955 <= 0;
      x75958 <= 0;
      x75961 <= 0;
      x75964 <= 0;
      x75967 <= 0;
      x75970 <= 0;
      x75973 <= 0;
      x75976 <= 0;
      x75979 <= 0;
      x75982 <= 0;
      x75985 <= 0;
      x75988 <= 0;
      x75991 <= 0;
      x75994 <= 0;
      x75997 <= 0;
      x76000 <= 0;
      x76003 <= 0;
      x76006 <= 0;
      x76009 <= 0;
      x76012 <= 0;
      x76015 <= 0;
      x76018 <= 0;
      x76021 <= 0;
      x76024 <= 0;
      x76027 <= 0;
      x76030 <= 0;
      x76033 <= 0;
      x76036 <= 0;
      x76039 <= 0;
      x76042 <= 0;
      x76045 <= 0;
      x76048 <= 0;
      x76051 <= 0;
      x76054 <= 0;
      x76057 <= 0;
      x76060 <= 0;
      x76063 <= 0;
      x76066 <= 0;
      x76069 <= 0;
      x76072 <= 0;
      x76075 <= 0;
      x76078 <= 0;
      x76081 <= 0;
      x76084 <= 0;
      x76087 <= 0;
      x76090 <= 0;
      x76093 <= 0;
      x76096 <= 0;
      x76099 <= 0;
      x76102 <= 0;
      x76105 <= 0;
      x76108 <= 0;
      x76111 <= 0;
      x76114 <= 0;
      x76117 <= 0;
      x76120 <= 0;
      x76123 <= 0;
      x76126 <= 0;
      x76129 <= 0;
      x76132 <= 0;
      x76135 <= 0;
      x76138 <= 0;
      x76141 <= 0;
      x76144 <= 0;
      x76147 <= 0;
      x76150 <= 0;
      x76153 <= 0;
      x76156 <= 0;
      x76159 <= 0;
      x76162 <= 0;
      x76165 <= 0;
      x76168 <= 0;
      x76171 <= 0;
      x76174 <= 0;
      x76177 <= 0;
      x76180 <= 0;
      x76183 <= 0;
      x76186 <= 0;
      x76189 <= 0;
      x76192 <= 0;
      x76195 <= 0;
      x76198 <= 0;
      x76201 <= 0;
      x76204 <= 0;
      x76207 <= 0;
      x76210 <= 0;
      x76213 <= 0;
      x76216 <= 0;
      x76219 <= 0;
      x76222 <= 0;
      x76225 <= 0;
      x76228 <= 0;
      x76231 <= 0;
      x76234 <= 0;
      x76237 <= 0;
      x76240 <= 0;
      x76243 <= 0;
      x76246 <= 0;
      x76249 <= 0;
      x76252 <= 0;
      x76255 <= 0;
      x76258 <= 0;
      x76261 <= 0;
      x76264 <= 0;
      x76267 <= 0;
      x76270 <= 0;
      x76273 <= 0;
      x76276 <= 0;
      x76279 <= 0;
      x76282 <= 0;
      x76285 <= 0;
      x76288 <= 0;
      x76291 <= 0;
      x76294 <= 0;
      x76297 <= 0;
      x76300 <= 0;
      x76303 <= 0;
      x76306 <= 0;
      x76309 <= 0;
      x76312 <= 0;
      x76315 <= 0;
      x76318 <= 0;
      x76321 <= 0;
      x76324 <= 0;
      x76327 <= 0;
      x76330 <= 0;
      x76333 <= 0;
      x76336 <= 0;
      x76339 <= 0;
      x76342 <= 0;
      x76345 <= 0;
      x76348 <= 0;
      x76351 <= 0;
      x76354 <= 0;
      x76357 <= 0;
      x76360 <= 0;
      x76363 <= 0;
      x76366 <= 0;
      x76369 <= 0;
      x76372 <= 0;
      x76375 <= 0;
      x76378 <= 0;
      x76381 <= 0;
      x76384 <= 0;
      x76387 <= 0;
      x76390 <= 0;
      x76393 <= 0;
      x76396 <= 0;
      x76399 <= 0;
      x76402 <= 0;
      x76405 <= 0;
      x76408 <= 0;
      x76411 <= 0;
      x76414 <= 0;
      x76417 <= 0;
      x76420 <= 0;
      x76423 <= 0;
      x76426 <= 0;
      x76429 <= 0;
      x76432 <= 0;
      x76435 <= 0;
      x76438 <= 0;
      x76441 <= 0;
      x76444 <= 0;
      x76447 <= 0;
      x76450 <= 0;
      x76453 <= 0;
      x76456 <= 0;
      x76459 <= 0;
      x76462 <= 0;
      x76465 <= 0;
      x76468 <= 0;
      x76471 <= 0;
      x76474 <= 0;
      x76477 <= 0;
      x76480 <= 0;
      x76483 <= 0;
      x76486 <= 0;
      x76489 <= 0;
      x76492 <= 0;
      x76495 <= 0;
      x76498 <= 0;
      x76501 <= 0;
      x76504 <= 0;
      x76507 <= 0;
      x76510 <= 0;
      x76513 <= 0;
      x76516 <= 0;
      x76519 <= 0;
      x76522 <= 0;
      x76525 <= 0;
      x76528 <= 0;
      x76531 <= 0;
      x76534 <= 0;
      x76537 <= 0;
      x76540 <= 0;
      x76543 <= 0;
      x76546 <= 0;
      x76549 <= 0;
      x76552 <= 0;
      x76555 <= 0;
      x76558 <= 0;
      x76561 <= 0;
      x76564 <= 0;
      x76567 <= 0;
      x76570 <= 0;
      x76573 <= 0;
      x76576 <= 0;
      x76579 <= 0;
      x76582 <= 0;
      x76585 <= 0;
      x76588 <= 0;
      x76591 <= 0;
      x76594 <= 0;
      x76597 <= 0;
      x76600 <= 0;
      x76603 <= 0;
      x76606 <= 0;
      x76609 <= 0;
      x76612 <= 0;
      x76615 <= 0;
      x76618 <= 0;
      x76621 <= 0;
      x76624 <= 0;
      x76627 <= 0;
      x76630 <= 0;
      x76633 <= 0;
      x76636 <= 0;
      x76639 <= 0;
      x76642 <= 0;
      x76645 <= 0;
      x76648 <= 0;
      x76651 <= 0;
      x76654 <= 0;
      x76657 <= 0;
      x76660 <= 0;
      x76663 <= 0;
      x76666 <= 0;
      x76669 <= 0;
      x76672 <= 0;
      x76675 <= 0;
      x76678 <= 0;
      x76681 <= 0;
      x76684 <= 0;
      x76687 <= 0;
      x76690 <= 0;
      x76693 <= 0;
      x76696 <= 0;
      x76699 <= 0;
      x76702 <= 0;
      x76705 <= 0;
      x76708 <= 0;
      x76711 <= 0;
      x76714 <= 0;
      x76717 <= 0;
      x76720 <= 0;
      x76723 <= 0;
      x76726 <= 0;
      x76729 <= 0;
      x76732 <= 0;
      x76735 <= 0;
      x76738 <= 0;
      x76741 <= 0;
      x76744 <= 0;
      x76747 <= 0;
      x76750 <= 0;
      x76753 <= 0;
      x76756 <= 0;
      x76759 <= 0;
      x76762 <= 0;
      x76765 <= 0;
      x76768 <= 0;
      x76771 <= 0;
      x76774 <= 0;
      x76777 <= 0;
      x76780 <= 0;
      x76783 <= 0;
      x76786 <= 0;
      x76789 <= 0;
      x76792 <= 0;
      x76795 <= 0;
      x76798 <= 0;
      x76801 <= 0;
      x76804 <= 0;
      x76807 <= 0;
      x76810 <= 0;
      x76813 <= 0;
      x76816 <= 0;
      x76819 <= 0;
      x76822 <= 0;
      x76825 <= 0;
      x76828 <= 0;
      x76831 <= 0;
      x76834 <= 0;
      x76837 <= 0;
      x76840 <= 0;
      x76843 <= 0;
      x76846 <= 0;
      x76849 <= 0;
      x76852 <= 0;
      x76855 <= 0;
      x76858 <= 0;
      x76861 <= 0;
      x76864 <= 0;
      x76867 <= 0;
      x76870 <= 0;
      x76873 <= 0;
      x76876 <= 0;
      x76879 <= 0;
      x76882 <= 0;
      x76885 <= 0;
      x76888 <= 0;
      x76891 <= 0;
      x76894 <= 0;
      x76897 <= 0;
      x76900 <= 0;
      x76903 <= 0;
      x76906 <= 0;
      x76909 <= 0;
      x76912 <= 0;
      x76915 <= 0;
      x76918 <= 0;
      x76921 <= 0;
      x76924 <= 0;
      x76927 <= 0;
      x76930 <= 0;
      x76933 <= 0;
      x76936 <= 0;
      x76939 <= 0;
      x76942 <= 0;
      x76945 <= 0;
      x76948 <= 0;
      x76951 <= 0;
      x76954 <= 0;
      x76957 <= 0;
      x76960 <= 0;
      x76963 <= 0;
      x76966 <= 0;
      x76969 <= 0;
      x76972 <= 0;
      x76975 <= 0;
      x76978 <= 0;
      x76981 <= 0;
      x76984 <= 0;
      x76987 <= 0;
      x76990 <= 0;
      x76993 <= 0;
      x76996 <= 0;
      x76999 <= 0;
      x77002 <= 0;
      x77005 <= 0;
      x77008 <= 0;
      x77011 <= 0;
      x77014 <= 0;
      x77017 <= 0;
      x77020 <= 0;
      x77023 <= 0;
      x77026 <= 0;
      x77029 <= 0;
      x77032 <= 0;
      x77035 <= 0;
      x77038 <= 0;
      x77041 <= 0;
      x77044 <= 0;
      x77047 <= 0;
      x77050 <= 0;
      x77053 <= 0;
      x77056 <= 0;
      x77059 <= 0;
      x77062 <= 0;
      x77065 <= 0;
      x77068 <= 0;
      x77071 <= 0;
      x77074 <= 0;
      x77077 <= 0;
      x77080 <= 0;
      x77083 <= 0;
      x77086 <= 0;
      x77089 <= 0;
      x77092 <= 0;
      x77095 <= 0;
      x77098 <= 0;
      x77101 <= 0;
      x77104 <= 0;
      x77107 <= 0;
      x77110 <= 0;
      x77113 <= 0;
      x77116 <= 0;
      x77119 <= 0;
      x77122 <= 0;
      x77125 <= 0;
      x77128 <= 0;
      x77131 <= 0;
      x77134 <= 0;
      x77137 <= 0;
      x77140 <= 0;
      x77143 <= 0;
      x77146 <= 0;
      x77149 <= 0;
      x77152 <= 0;
      x77155 <= 0;
      x77158 <= 0;
      x77161 <= 0;
      x77164 <= 0;
      x77167 <= 0;
      x77170 <= 0;
      x77173 <= 0;
      x77176 <= 0;
      x77179 <= 0;
      x77182 <= 0;
      x77185 <= 0;
      x77188 <= 0;
      x77191 <= 0;
      x77194 <= 0;
      x77197 <= 0;
      x77200 <= 0;
      x77203 <= 0;
      x77206 <= 0;
      x77209 <= 0;
      x77212 <= 0;
      x77215 <= 0;
      x77218 <= 0;
      x77221 <= 0;
      x77224 <= 0;
      x77227 <= 0;
      x77230 <= 0;
      x77233 <= 0;
      x77236 <= 0;
      x77239 <= 0;
      x77242 <= 0;
      x77245 <= 0;
      x77248 <= 0;
      x77251 <= 0;
      x77254 <= 0;
      x77257 <= 0;
      x77260 <= 0;
      x77263 <= 0;
      x77266 <= 0;
      x77269 <= 0;
      x77272 <= 0;
      x77275 <= 0;
      x77278 <= 0;
      x77281 <= 0;
      x77284 <= 0;
      x77287 <= 0;
      x77290 <= 0;
      x77293 <= 0;
      x77296 <= 0;
      x77299 <= 0;
      x77302 <= 0;
      x77305 <= 0;
      x77308 <= 0;
      x77311 <= 0;
      x77314 <= 0;
      x77317 <= 0;
      x77320 <= 0;
      x77323 <= 0;
      x77326 <= 0;
      x77329 <= 0;
      x77332 <= 0;
      x77335 <= 0;
      x77338 <= 0;
      x77341 <= 0;
      x77344 <= 0;
      x77347 <= 0;
      x77350 <= 0;
      x77353 <= 0;
      x77356 <= 0;
      x77359 <= 0;
      x77362 <= 0;
      x77365 <= 0;
      x77368 <= 0;
      x77371 <= 0;
      x77374 <= 0;
      x77377 <= 0;
      x77380 <= 0;
      x77383 <= 0;
      x77386 <= 0;
      x77389 <= 0;
      x77392 <= 0;
      x77395 <= 0;
      x77398 <= 0;
      x77401 <= 0;
      x77404 <= 0;
      x77407 <= 0;
      x77410 <= 0;
      x77413 <= 0;
      x77416 <= 0;
      x77419 <= 0;
      x77422 <= 0;
      x77425 <= 0;
      x77428 <= 0;
      x77431 <= 0;
      x77434 <= 0;
      x77437 <= 0;
      x77440 <= 0;
      x77443 <= 0;
      x77446 <= 0;
      x77449 <= 0;
      x77452 <= 0;
      x77455 <= 0;
      x77458 <= 0;
      x77461 <= 0;
      x77464 <= 0;
      x77467 <= 0;
      x77470 <= 0;
      x77473 <= 0;
      x77476 <= 0;
      x77479 <= 0;
      x77482 <= 0;
      x77485 <= 0;
      x77488 <= 0;
      x77491 <= 0;
      x77494 <= 0;
      x77497 <= 0;
      x77500 <= 0;
      x77503 <= 0;
      x77506 <= 0;
      x77509 <= 0;
      x77512 <= 0;
      x77515 <= 0;
      x77518 <= 0;
      x77521 <= 0;
      x77524 <= 0;
      x77527 <= 0;
      x77530 <= 0;
      x77533 <= 0;
      x77536 <= 0;
      x77539 <= 0;
      x77542 <= 0;
      x77545 <= 0;
      x77548 <= 0;
      x77551 <= 0;
      x77554 <= 0;
      x77557 <= 0;
      x77560 <= 0;
      x77563 <= 0;
      x77566 <= 0;
      x77569 <= 0;
      x77572 <= 0;
      x77575 <= 0;
      x77578 <= 0;
      x77581 <= 0;
      x77584 <= 0;
      x77587 <= 0;
      x77590 <= 0;
      x77593 <= 0;
      x77596 <= 0;
      x77599 <= 0;
      x77602 <= 0;
      x77605 <= 0;
      x77608 <= 0;
      x77611 <= 0;
      x77614 <= 0;
      x77617 <= 0;
      x77620 <= 0;
      x77623 <= 0;
      x77626 <= 0;
      x77629 <= 0;
      x77632 <= 0;
      x77635 <= 0;
      x77638 <= 0;
      x77641 <= 0;
      x77644 <= 0;
      x77647 <= 0;
      x77650 <= 0;
      x77653 <= 0;
      x77656 <= 0;
      x77659 <= 0;
      x77662 <= 0;
      x77665 <= 0;
      x77668 <= 0;
      x77671 <= 0;
      x77674 <= 0;
      x77677 <= 0;
      x77680 <= 0;
      x77683 <= 0;
      x77686 <= 0;
      x77689 <= 0;
      x77692 <= 0;
      x77695 <= 0;
      x77698 <= 0;
      x77701 <= 0;
      x77704 <= 0;
      x77707 <= 0;
      x77710 <= 0;
      x77713 <= 0;
      x77716 <= 0;
      x77719 <= 0;
      x77722 <= 0;
      x77725 <= 0;
      x77728 <= 0;
      x77731 <= 0;
      x77734 <= 0;
      x77737 <= 0;
      x77740 <= 0;
      x77743 <= 0;
      x77746 <= 0;
      x77749 <= 0;
      x77752 <= 0;
      x77755 <= 0;
      x77758 <= 0;
      x77761 <= 0;
      x77764 <= 0;
      x77767 <= 0;
      x77770 <= 0;
      x77773 <= 0;
      x77776 <= 0;
      x77779 <= 0;
      x77782 <= 0;
      x77785 <= 0;
      x77788 <= 0;
      x77791 <= 0;
      x77794 <= 0;
      x77797 <= 0;
      x77800 <= 0;
      x77803 <= 0;
      x77806 <= 0;
      x77809 <= 0;
      x77812 <= 0;
      x77815 <= 0;
      x77818 <= 0;
      x77821 <= 0;
      x77824 <= 0;
      x77827 <= 0;
      x77830 <= 0;
      x77833 <= 0;
      x77836 <= 0;
      x77839 <= 0;
      x77842 <= 0;
      x77845 <= 0;
      x77848 <= 0;
      x77851 <= 0;
      x77854 <= 0;
      x77857 <= 0;
      x77860 <= 0;
      x77863 <= 0;
      x77866 <= 0;
      x77869 <= 0;
      x77872 <= 0;
      x77875 <= 0;
      x77878 <= 0;
      x77881 <= 0;
      x77884 <= 0;
      x77887 <= 0;
      x77890 <= 0;
      x77893 <= 0;
      x77896 <= 0;
      x77899 <= 0;
      x77902 <= 0;
      x77905 <= 0;
      x77908 <= 0;
      x77911 <= 0;
      x77914 <= 0;
      x77917 <= 0;
      x77920 <= 0;
      x77923 <= 0;
      x77926 <= 0;
      x77929 <= 0;
      x77932 <= 0;
      x77935 <= 0;
      x77938 <= 0;
      x77941 <= 0;
      x77944 <= 0;
      x77947 <= 0;
      x77950 <= 0;
      x77953 <= 0;
      x77956 <= 0;
      x77959 <= 0;
      x77962 <= 0;
      x77965 <= 0;
      x77968 <= 0;
      x77971 <= 0;
      x77974 <= 0;
      x77977 <= 0;
      x77980 <= 0;
      x77983 <= 0;
      x77986 <= 0;
      x77989 <= 0;
      x77992 <= 0;
      x77995 <= 0;
      x77998 <= 0;
      x78001 <= 0;
      x78004 <= 0;
      x78007 <= 0;
      x78010 <= 0;
      x78013 <= 0;
      x78016 <= 0;
      x78019 <= 0;
      x78022 <= 0;
      x78025 <= 0;
      x78028 <= 0;
      x78031 <= 0;
      x78034 <= 0;
      x78037 <= 0;
      x78040 <= 0;
      x78043 <= 0;
      x78046 <= 0;
      x78049 <= 0;
      x78052 <= 0;
      x78055 <= 0;
      x78058 <= 0;
      x78061 <= 0;
      x78064 <= 0;
      x78067 <= 0;
      x78070 <= 0;
      x78073 <= 0;
      x78076 <= 0;
      x78079 <= 0;
      x78082 <= 0;
      x78085 <= 0;
      x78088 <= 0;
      x78091 <= 0;
      x78094 <= 0;
      x78097 <= 0;
      x78100 <= 0;
      x78103 <= 0;
      x78106 <= 0;
      x78109 <= 0;
      x78112 <= 0;
      x78115 <= 0;
      x78118 <= 0;
      x78121 <= 0;
      x78124 <= 0;
      x78127 <= 0;
      x78130 <= 0;
      x78133 <= 0;
      x78136 <= 0;
      x78139 <= 0;
      x78142 <= 0;
      x78145 <= 0;
      x78148 <= 0;
      x78151 <= 0;
      x78154 <= 0;
      x78157 <= 0;
      x78160 <= 0;
      x78163 <= 0;
      x78166 <= 0;
      x78169 <= 0;
      x78172 <= 0;
      x78175 <= 0;
      x78178 <= 0;
      x78181 <= 0;
      x78184 <= 0;
      x78187 <= 0;
      x78190 <= 0;
      x78193 <= 0;
      x78196 <= 0;
      x78199 <= 0;
      x78202 <= 0;
      x78205 <= 0;
      x78208 <= 0;
      x78211 <= 0;
      x78214 <= 0;
      x78217 <= 0;
      x78220 <= 0;
      x78223 <= 0;
      x78226 <= 0;
      x78229 <= 0;
      x78232 <= 0;
      x78235 <= 0;
      x78238 <= 0;
      x78241 <= 0;
      x78244 <= 0;
      x78247 <= 0;
      x78250 <= 0;
      x78253 <= 0;
      x78256 <= 0;
      x78259 <= 0;
      x78262 <= 0;
      x78265 <= 0;
      x78268 <= 0;
      x78271 <= 0;
      x78274 <= 0;
      x78277 <= 0;
      x78280 <= 0;
      x78283 <= 0;
      x78286 <= 0;
      x78289 <= 0;
      x78292 <= 0;
      x78295 <= 0;
      x78298 <= 0;
      x78301 <= 0;
      x78304 <= 0;
      x78307 <= 0;
      x78310 <= 0;
      x78313 <= 0;
      x78316 <= 0;
      x78319 <= 0;
      x78322 <= 0;
      x78325 <= 0;
      x78328 <= 0;
      x78331 <= 0;
      x78334 <= 0;
      x78337 <= 0;
      x78340 <= 0;
      x78343 <= 0;
      x78346 <= 0;
      x78349 <= 0;
      x78352 <= 0;
      x78355 <= 0;
      x78358 <= 0;
      x78361 <= 0;
      x78364 <= 0;
      x78367 <= 0;
      x78370 <= 0;
      x78373 <= 0;
      x78376 <= 0;
      x78379 <= 0;
      x78382 <= 0;
      x78385 <= 0;
      x78388 <= 0;
      x78391 <= 0;
      x78394 <= 0;
      x78397 <= 0;
      x78400 <= 0;
      x78403 <= 0;
      x78406 <= 0;
      x78409 <= 0;
      x78412 <= 0;
      x78415 <= 0;
      x78418 <= 0;
      x78421 <= 0;
      x78424 <= 0;
      x78427 <= 0;
      x78430 <= 0;
      x78433 <= 0;
      x78436 <= 0;
      x78439 <= 0;
      x78442 <= 0;
      x78445 <= 0;
      x78448 <= 0;
      x78451 <= 0;
      x78454 <= 0;
      x78457 <= 0;
      x78460 <= 0;
      x78463 <= 0;
      x78466 <= 0;
      x78469 <= 0;
      x78472 <= 0;
      x78475 <= 0;
      x78478 <= 0;
      x78481 <= 0;
      x78484 <= 0;
      x78487 <= 0;
      x78490 <= 0;
      x78493 <= 0;
      x78496 <= 0;
      x78499 <= 0;
      x78502 <= 0;
      x78505 <= 0;
      x78508 <= 0;
      x78511 <= 0;
      x78514 <= 0;
      x78517 <= 0;
      x78520 <= 0;
      x78523 <= 0;
      x78526 <= 0;
      x78529 <= 0;
      x78532 <= 0;
      x78535 <= 0;
      x78538 <= 0;
      x78541 <= 0;
      x78544 <= 0;
      x78547 <= 0;
      x78550 <= 0;
      x78553 <= 0;
      x78556 <= 0;
      x78559 <= 0;
      x78562 <= 0;
      x78565 <= 0;
      x78568 <= 0;
      x78571 <= 0;
      x78574 <= 0;
      x78577 <= 0;
      x78580 <= 0;
      x78583 <= 0;
      x78586 <= 0;
      x78589 <= 0;
      x78592 <= 0;
      x78595 <= 0;
      x78598 <= 0;
      x78601 <= 0;
      x78604 <= 0;
      x78607 <= 0;
      x78610 <= 0;
      x78613 <= 0;
      x78616 <= 0;
      x78619 <= 0;
      x78622 <= 0;
      x78625 <= 0;
      x78628 <= 0;
      x78631 <= 0;
      x78634 <= 0;
      x78637 <= 0;
      x78640 <= 0;
      x78643 <= 0;
      x78646 <= 0;
      x78649 <= 0;
      x78652 <= 0;
      x78655 <= 0;
      x78658 <= 0;
      x78661 <= 0;
      x78664 <= 0;
      x78667 <= 0;
      x78670 <= 0;
      x78673 <= 0;
      x78676 <= 0;
      x78679 <= 0;
      x78682 <= 0;
      x78685 <= 0;
      x78688 <= 0;
      x78691 <= 0;
      x78694 <= 0;
      x78697 <= 0;
      x78700 <= 0;
      x78703 <= 0;
      x78706 <= 0;
      x78709 <= 0;
      x78712 <= 0;
      x78715 <= 0;
      x78718 <= 0;
      x78721 <= 0;
      x78724 <= 0;
      x78727 <= 0;
      x78730 <= 0;
      x78733 <= 0;
      x78736 <= 0;
      x78739 <= 0;
      x78742 <= 0;
      x78745 <= 0;
      x78748 <= 0;
      x78751 <= 0;
      x78754 <= 0;
      x78757 <= 0;
      x78760 <= 0;
      x78763 <= 0;
      x78766 <= 0;
      x78769 <= 0;
      x78772 <= 0;
      x78775 <= 0;
      x78778 <= 0;
      x78781 <= 0;
      x78784 <= 0;
      x78787 <= 0;
      x78790 <= 0;
      x78793 <= 0;
      x78796 <= 0;
      x78799 <= 0;
      x78802 <= 0;
      x78805 <= 0;
      x78808 <= 0;
      x78811 <= 0;
      x78814 <= 0;
      x78817 <= 0;
      x78820 <= 0;
      x78823 <= 0;
      x78826 <= 0;
      x78829 <= 0;
      x78832 <= 0;
      x78835 <= 0;
      x78838 <= 0;
      x78841 <= 0;
      x78844 <= 0;
      x78847 <= 0;
      x78850 <= 0;
      x78853 <= 0;
      x78856 <= 0;
      x78859 <= 0;
      x78862 <= 0;
      x78865 <= 0;
      x78868 <= 0;
      x78871 <= 0;
      x78874 <= 0;
      x78877 <= 0;
      x78880 <= 0;
      x78883 <= 0;
      x78886 <= 0;
      x78889 <= 0;
      x78892 <= 0;
      x78895 <= 0;
      x78898 <= 0;
      x78901 <= 0;
      x78904 <= 0;
      x78907 <= 0;
      x78910 <= 0;
      x78913 <= 0;
      x78916 <= 0;
      x78919 <= 0;
      x78922 <= 0;
      x78925 <= 0;
      x78928 <= 0;
      x78931 <= 0;
      x78934 <= 0;
      x78937 <= 0;
      x78940 <= 0;
      x78943 <= 0;
      x78946 <= 0;
      x78949 <= 0;
      x78952 <= 0;
      x78955 <= 0;
      x78958 <= 0;
      x78961 <= 0;
      x78964 <= 0;
      x78967 <= 0;
      x78970 <= 0;
      x78973 <= 0;
      x78976 <= 0;
      x78979 <= 0;
      x78982 <= 0;
      x78985 <= 0;
      x78988 <= 0;
      x78991 <= 0;
      x78994 <= 0;
      x78997 <= 0;
      x79000 <= 0;
      x79003 <= 0;
      x79006 <= 0;
      x79009 <= 0;
      x79012 <= 0;
      x79015 <= 0;
      x79018 <= 0;
      x79021 <= 0;
      x79024 <= 0;
      x79027 <= 0;
      x79030 <= 0;
      x79033 <= 0;
      x79036 <= 0;
      x79039 <= 0;
      x79042 <= 0;
      x79045 <= 0;
      x79048 <= 0;
      x79051 <= 0;
      x79054 <= 0;
      x79057 <= 0;
      x79060 <= 0;
      x79063 <= 0;
      x79066 <= 0;
      x79069 <= 0;
      x79072 <= 0;
      x79075 <= 0;
      x79078 <= 0;
      x79081 <= 0;
      x79084 <= 0;
      x79087 <= 0;
      x79090 <= 0;
      x79093 <= 0;
      x79096 <= 0;
      x79099 <= 0;
      x79102 <= 0;
      x79105 <= 0;
      x79108 <= 0;
      x79111 <= 0;
      x79114 <= 0;
      x79117 <= 0;
      x79120 <= 0;
      x79123 <= 0;
      x79126 <= 0;
      x79129 <= 0;
      x79132 <= 0;
      x79135 <= 0;
      x79138 <= 0;
      x79141 <= 0;
      x79144 <= 0;
      x79147 <= 0;
      x79150 <= 0;
      x79153 <= 0;
      x79156 <= 0;
      x79159 <= 0;
      x79162 <= 0;
      x79165 <= 0;
      x79168 <= 0;
      x79171 <= 0;
      x79174 <= 0;
      x79177 <= 0;
      x79180 <= 0;
      x79183 <= 0;
      x79186 <= 0;
      x79189 <= 0;
      x79192 <= 0;
      x79195 <= 0;
      x79198 <= 0;
      x79201 <= 0;
      x79204 <= 0;
      x79207 <= 0;
      x79210 <= 0;
      x79213 <= 0;
      x79216 <= 0;
      x79219 <= 0;
      x79222 <= 0;
      x79225 <= 0;
      x79228 <= 0;
      x79231 <= 0;
      x79234 <= 0;
      x79237 <= 0;
      x79240 <= 0;
      x79243 <= 0;
      x79246 <= 0;
      x79249 <= 0;
      x79252 <= 0;
      x79255 <= 0;
      x79258 <= 0;
      x79261 <= 0;
      x79264 <= 0;
      x79267 <= 0;
      x79270 <= 0;
      x79273 <= 0;
      x79276 <= 0;
      x79279 <= 0;
      x79282 <= 0;
      x79285 <= 0;
      x79288 <= 0;
      x79291 <= 0;
      x79294 <= 0;
      x79297 <= 0;
      x79300 <= 0;
      x79303 <= 0;
      x79306 <= 0;
      x79309 <= 0;
      x79312 <= 0;
      x79315 <= 0;
      x79318 <= 0;
      x79321 <= 0;
      x79324 <= 0;
      x79327 <= 0;
      x79330 <= 0;
      x79333 <= 0;
      x79336 <= 0;
      x79339 <= 0;
      x79342 <= 0;
      x79345 <= 0;
      x79348 <= 0;
      x79351 <= 0;
      x79354 <= 0;
      x79357 <= 0;
      x79360 <= 0;
      x79363 <= 0;
      x79366 <= 0;
      x79369 <= 0;
      x79372 <= 0;
      x79375 <= 0;
      x79378 <= 0;
      x79381 <= 0;
      x79384 <= 0;
      x79387 <= 0;
      x79390 <= 0;
      x79393 <= 0;
      x79396 <= 0;
      x79399 <= 0;
      x79402 <= 0;
      x79405 <= 0;
      x79408 <= 0;
      x79411 <= 0;
      x79414 <= 0;
      x79417 <= 0;
      x79420 <= 0;
      x79423 <= 0;
      x79426 <= 0;
      x79429 <= 0;
      x79432 <= 0;
      x79435 <= 0;
      x79438 <= 0;
      x79441 <= 0;
      x79444 <= 0;
      x79447 <= 0;
      x79450 <= 0;
      x79453 <= 0;
      x79456 <= 0;
      x79459 <= 0;
      x79462 <= 0;
      x79465 <= 0;
      x79468 <= 0;
      x79471 <= 0;
      x79474 <= 0;
      x79477 <= 0;
      x79480 <= 0;
      x79483 <= 0;
      x79486 <= 0;
      x79489 <= 0;
      x79492 <= 0;
      x79495 <= 0;
      x79498 <= 0;
      x79501 <= 0;
      x79504 <= 0;
      x79507 <= 0;
      x79510 <= 0;
      x79513 <= 0;
      x79516 <= 0;
      x79519 <= 0;
      x79522 <= 0;
      x79525 <= 0;
      x79528 <= 0;
      x79531 <= 0;
      x79534 <= 0;
      x79537 <= 0;
      x79540 <= 0;
      x79543 <= 0;
      x79546 <= 0;
      x79549 <= 0;
      x79552 <= 0;
      x79555 <= 0;
      x79558 <= 0;
      x79561 <= 0;
      x79564 <= 0;
      x79567 <= 0;
      x79570 <= 0;
      x79573 <= 0;
      x79576 <= 0;
      x79579 <= 0;
      x79582 <= 0;
      x79585 <= 0;
      x79588 <= 0;
      x79591 <= 0;
      x79594 <= 0;
      x79597 <= 0;
      x79600 <= 0;
      x79603 <= 0;
      x79606 <= 0;
      x79609 <= 0;
      x79612 <= 0;
      x79615 <= 0;
      x79618 <= 0;
      x79621 <= 0;
      x79624 <= 0;
      x79627 <= 0;
      x79630 <= 0;
      x79633 <= 0;
      x79636 <= 0;
      x79639 <= 0;
      x79642 <= 0;
      x79645 <= 0;
      x79648 <= 0;
      x79651 <= 0;
      x79654 <= 0;
      x79657 <= 0;
      x79660 <= 0;
      x79663 <= 0;
      x79666 <= 0;
      x79669 <= 0;
      x79672 <= 0;
      x79675 <= 0;
      x79678 <= 0;
      x79681 <= 0;
      x79684 <= 0;
      x79687 <= 0;
      x79690 <= 0;
      x79693 <= 0;
      x79696 <= 0;
      x79699 <= 0;
      x79702 <= 0;
      x79705 <= 0;
      x79708 <= 0;
      x79711 <= 0;
      x79714 <= 0;
      x79717 <= 0;
      x79720 <= 0;
      x79723 <= 0;
      x79726 <= 0;
      x79729 <= 0;
      x79732 <= 0;
      x79735 <= 0;
      x79738 <= 0;
      x79741 <= 0;
      x79744 <= 0;
      x79747 <= 0;
      x79750 <= 0;
      x79753 <= 0;
      x79756 <= 0;
      x79759 <= 0;
      x79762 <= 0;
      x79765 <= 0;
      x79768 <= 0;
      x79771 <= 0;
      x79774 <= 0;
      x79777 <= 0;
      x79780 <= 0;
      x79783 <= 0;
      x79786 <= 0;
      x79789 <= 0;
      x79792 <= 0;
      x79795 <= 0;
      x79798 <= 0;
      x79801 <= 0;
      x79804 <= 0;
      x79807 <= 0;
      x79810 <= 0;
      x79813 <= 0;
      x79816 <= 0;
      x79819 <= 0;
      x79822 <= 0;
      x79825 <= 0;
      x79828 <= 0;
      x79831 <= 0;
      x79834 <= 0;
      x79837 <= 0;
      x79840 <= 0;
      x79843 <= 0;
      x79846 <= 0;
      x79849 <= 0;
      x79852 <= 0;
      x79855 <= 0;
      x79858 <= 0;
      x79861 <= 0;
      x79864 <= 0;
      x79867 <= 0;
      x79870 <= 0;
      x79873 <= 0;
      x79876 <= 0;
      x79879 <= 0;
      x79882 <= 0;
      x79885 <= 0;
      x79888 <= 0;
      x79891 <= 0;
      x79894 <= 0;
      x79897 <= 0;
      x79900 <= 0;
      x79903 <= 0;
      x79906 <= 0;
      x79909 <= 0;
      x79912 <= 0;
      x79915 <= 0;
      x79918 <= 0;
      x79921 <= 0;
      x79924 <= 0;
      x79927 <= 0;
      x79930 <= 0;
      x79933 <= 0;
      x79936 <= 0;
      x79939 <= 0;
      x79942 <= 0;
      x79945 <= 0;
      x79948 <= 0;
      x79951 <= 0;
      x79954 <= 0;
      x79957 <= 0;
      x79960 <= 0;
      x79963 <= 0;
      x79966 <= 0;
      x79969 <= 0;
      x79972 <= 0;
      x79975 <= 0;
      x79978 <= 0;
      x79981 <= 0;
      x79984 <= 0;
      x79987 <= 0;
      x79990 <= 0;
      x79993 <= 0;
      x79996 <= 0;
      x79999 <= 0;
      x80002 <= 0;
      x80005 <= 0;
      x80008 <= 0;
      x80011 <= 0;
      x80014 <= 0;
      x80017 <= 0;
      x80020 <= 0;
      x80023 <= 0;
      x80026 <= 0;
      x80029 <= 0;
      x80032 <= 0;
      x80035 <= 0;
      x80038 <= 0;
      x80041 <= 0;
      x80044 <= 0;
      x80047 <= 0;
      x80050 <= 0;
      x80053 <= 0;
      x80056 <= 0;
      x80059 <= 0;
      x80062 <= 0;
      x80065 <= 0;
      x80068 <= 0;
      x80071 <= 0;
      x80074 <= 0;
      x80077 <= 0;
      x80080 <= 0;
      x80083 <= 0;
      x80086 <= 0;
      x80089 <= 0;
      x80092 <= 0;
      x80095 <= 0;
      x80098 <= 0;
      x80101 <= 0;
      x80104 <= 0;
      x80107 <= 0;
      x80110 <= 0;
      x80113 <= 0;
      x80116 <= 0;
      x80119 <= 0;
      x80122 <= 0;
      x80125 <= 0;
      x80128 <= 0;
      x80131 <= 0;
      x80134 <= 0;
      x80137 <= 0;
      x80140 <= 0;
      x80143 <= 0;
      x80146 <= 0;
      x80149 <= 0;
      x80152 <= 0;
      x80155 <= 0;
      x80158 <= 0;
      x80161 <= 0;
      x80164 <= 0;
      x80167 <= 0;
      x80170 <= 0;
      x80173 <= 0;
      x80176 <= 0;
      x80179 <= 0;
      x80182 <= 0;
      x80185 <= 0;
      x80188 <= 0;
      x80191 <= 0;
      x80194 <= 0;
      x80197 <= 0;
      x80200 <= 0;
      x80203 <= 0;
      x80206 <= 0;
      x80209 <= 0;
      x80212 <= 0;
      x80215 <= 0;
      x80218 <= 0;
      x80221 <= 0;
      x80224 <= 0;
      x80227 <= 0;
      x80230 <= 0;
      x80233 <= 0;
      x80236 <= 0;
      x80239 <= 0;
      x80242 <= 0;
      x80245 <= 0;
      x80248 <= 0;
      x80251 <= 0;
      x80254 <= 0;
      x80257 <= 0;
      x80260 <= 0;
      x80263 <= 0;
      x80266 <= 0;
      x80269 <= 0;
      x80272 <= 0;
      x80275 <= 0;
      x80278 <= 0;
      x80281 <= 0;
      x80284 <= 0;
      x80287 <= 0;
      x80290 <= 0;
      x80293 <= 0;
      x80296 <= 0;
      x80299 <= 0;
      x80302 <= 0;
      x80305 <= 0;
      x80308 <= 0;
      x80311 <= 0;
      x80314 <= 0;
      x80317 <= 0;
      x80320 <= 0;
      x80323 <= 0;
      x80326 <= 0;
      x80329 <= 0;
      x80332 <= 0;
      x80335 <= 0;
      x80338 <= 0;
      x80341 <= 0;
      x80344 <= 0;
      x80347 <= 0;
      x80350 <= 0;
      x80353 <= 0;
      x80356 <= 0;
      x80359 <= 0;
      x80362 <= 0;
      x80365 <= 0;
      x80368 <= 0;
      x80371 <= 0;
      x80374 <= 0;
      x80377 <= 0;
      x80380 <= 0;
      x80383 <= 0;
      x80386 <= 0;
      x80389 <= 0;
      x80392 <= 0;
      x80395 <= 0;
      x80398 <= 0;
      x80401 <= 0;
      x80404 <= 0;
      x80407 <= 0;
      x80410 <= 0;
      x80413 <= 0;
      x80416 <= 0;
      x80419 <= 0;
      x80422 <= 0;
      x80425 <= 0;
      x80428 <= 0;
      x80431 <= 0;
      x80434 <= 0;
      x80437 <= 0;
      x80440 <= 0;
      x80443 <= 0;
      x80446 <= 0;
      x80449 <= 0;
      x80452 <= 0;
      x80455 <= 0;
      x80458 <= 0;
      x80461 <= 0;
      x80464 <= 0;
      x80467 <= 0;
      x80470 <= 0;
      x80473 <= 0;
      x80476 <= 0;
      x80479 <= 0;
      x80482 <= 0;
      x80485 <= 0;
      x80488 <= 0;
      x80491 <= 0;
      x80494 <= 0;
      x80497 <= 0;
      x80500 <= 0;
      x80503 <= 0;
      x80506 <= 0;
      x80509 <= 0;
      x80512 <= 0;
      x80515 <= 0;
      x80518 <= 0;
      x80521 <= 0;
      x80524 <= 0;
      x80527 <= 0;
      x80530 <= 0;
      x80533 <= 0;
      x80536 <= 0;
      x80539 <= 0;
      x80542 <= 0;
      x80545 <= 0;
      x80548 <= 0;
      x80551 <= 0;
      x80554 <= 0;
      x80557 <= 0;
      x80560 <= 0;
      x80563 <= 0;
      x80566 <= 0;
      x80569 <= 0;
      x80572 <= 0;
      x80575 <= 0;
      x80578 <= 0;
      x80581 <= 0;
      x80584 <= 0;
      x80587 <= 0;
      x80590 <= 0;
      x80593 <= 0;
      x80596 <= 0;
      x80599 <= 0;
      x80602 <= 0;
      x80605 <= 0;
      x80608 <= 0;
      x80611 <= 0;
      x80614 <= 0;
      x80617 <= 0;
      x80620 <= 0;
      x80623 <= 0;
      x80626 <= 0;
      x80629 <= 0;
      x80632 <= 0;
      x80635 <= 0;
      x80638 <= 0;
      x80641 <= 0;
      x80644 <= 0;
      x80647 <= 0;
      x80650 <= 0;
      x80653 <= 0;
      x80656 <= 0;
      x80659 <= 0;
      x80662 <= 0;
      x80665 <= 0;
      x80668 <= 0;
      x80671 <= 0;
      x80674 <= 0;
      x80677 <= 0;
      x80680 <= 0;
      x80683 <= 0;
      x80686 <= 0;
      x80689 <= 0;
      x80692 <= 0;
      x80695 <= 0;
      x80698 <= 0;
      x80701 <= 0;
      x80704 <= 0;
      x80707 <= 0;
      x80710 <= 0;
      x80713 <= 0;
      x80716 <= 0;
      x80719 <= 0;
      x80722 <= 0;
      x80725 <= 0;
      x80728 <= 0;
      x80731 <= 0;
      x80734 <= 0;
      x80737 <= 0;
      x80740 <= 0;
      x80743 <= 0;
      x80746 <= 0;
      x80749 <= 0;
      x80752 <= 0;
      x80755 <= 0;
      x80758 <= 0;
      x80761 <= 0;
      x80764 <= 0;
      x80767 <= 0;
      x80770 <= 0;
      x80773 <= 0;
      x80776 <= 0;
      x80779 <= 0;
      x80782 <= 0;
      x80785 <= 0;
      x80788 <= 0;
      x80791 <= 0;
      x80794 <= 0;
      x80797 <= 0;
      x80800 <= 0;
      x80803 <= 0;
      x80806 <= 0;
      x80809 <= 0;
      x80812 <= 0;
      x80815 <= 0;
      x80818 <= 0;
      x80821 <= 0;
      x80824 <= 0;
      x80827 <= 0;
      x80830 <= 0;
      x80833 <= 0;
      x80836 <= 0;
      x80839 <= 0;
      x80842 <= 0;
      x80845 <= 0;
      x80848 <= 0;
      x80851 <= 0;
      x80854 <= 0;
      x80857 <= 0;
      x80860 <= 0;
      x80863 <= 0;
      x80866 <= 0;
      x80869 <= 0;
      x80872 <= 0;
      x80875 <= 0;
      x80878 <= 0;
      x80881 <= 0;
      x80884 <= 0;
      x80887 <= 0;
      x80890 <= 0;
      x80893 <= 0;
      x80896 <= 0;
      x80899 <= 0;
      x80902 <= 0;
      x80905 <= 0;
      x80908 <= 0;
      x80911 <= 0;
      x80914 <= 0;
      x80917 <= 0;
      x80920 <= 0;
      x80923 <= 0;
      x80926 <= 0;
      x80929 <= 0;
      x80932 <= 0;
      x80935 <= 0;
      x80938 <= 0;
      x80941 <= 0;
      x80944 <= 0;
      x80947 <= 0;
      x80950 <= 0;
      x80953 <= 0;
      x80956 <= 0;
      x80959 <= 0;
      x80962 <= 0;
      x80965 <= 0;
      x80968 <= 0;
      x80971 <= 0;
      x80974 <= 0;
      x80977 <= 0;
      x80980 <= 0;
      x80983 <= 0;
      x80986 <= 0;
      x80989 <= 0;
      x80992 <= 0;
      x80995 <= 0;
      x80998 <= 0;
      x81001 <= 0;
      x81004 <= 0;
      x81007 <= 0;
      x81010 <= 0;
      x81013 <= 0;
      x81016 <= 0;
      x81019 <= 0;
      x81022 <= 0;
      x81025 <= 0;
      x81028 <= 0;
      x81031 <= 0;
      x81034 <= 0;
      x81037 <= 0;
      x81040 <= 0;
      x81043 <= 0;
      x81046 <= 0;
      x81049 <= 0;
      x81052 <= 0;
      x81055 <= 0;
      x81058 <= 0;
      x81061 <= 0;
      x81064 <= 0;
      x81067 <= 0;
      x81070 <= 0;
      x81073 <= 0;
      x81076 <= 0;
      x81079 <= 0;
      x81082 <= 0;
      x81085 <= 0;
      x81088 <= 0;
      x81091 <= 0;
      x81094 <= 0;
      x81097 <= 0;
      x81100 <= 0;
      x81103 <= 0;
      x81106 <= 0;
      x81109 <= 0;
      x81112 <= 0;
      x81115 <= 0;
      x81118 <= 0;
      x81121 <= 0;
      x81124 <= 0;
      x81127 <= 0;
      x81130 <= 0;
      x81133 <= 0;
      x81136 <= 0;
      x81139 <= 0;
      x81142 <= 0;
      x81145 <= 0;
      x81148 <= 0;
      x81151 <= 0;
      x81154 <= 0;
      x81157 <= 0;
      x81160 <= 0;
      x81163 <= 0;
      x81166 <= 0;
      x81169 <= 0;
      x81172 <= 0;
      x81175 <= 0;
      x81178 <= 0;
      x81181 <= 0;
      x81184 <= 0;
      x81187 <= 0;
      x81190 <= 0;
      x81193 <= 0;
      x81196 <= 0;
      x81199 <= 0;
      x81202 <= 0;
      x81205 <= 0;
      x81208 <= 0;
      x81211 <= 0;
      x81214 <= 0;
      x81217 <= 0;
      x81220 <= 0;
      x81223 <= 0;
      x81226 <= 0;
      x81229 <= 0;
      x81232 <= 0;
      x81235 <= 0;
      x81238 <= 0;
      x81241 <= 0;
      x81244 <= 0;
      x81247 <= 0;
      x81250 <= 0;
      x81253 <= 0;
      x81256 <= 0;
      x81259 <= 0;
      x81262 <= 0;
      x81265 <= 0;
      x81268 <= 0;
      x81271 <= 0;
      x81274 <= 0;
      x81277 <= 0;
      x81280 <= 0;
      x81283 <= 0;
      x81286 <= 0;
      x81289 <= 0;
      x81292 <= 0;
      x81295 <= 0;
      x81298 <= 0;
      x81301 <= 0;
      x81304 <= 0;
      x81307 <= 0;
      x81310 <= 0;
      x81313 <= 0;
      x81316 <= 0;
      x81319 <= 0;
      x81322 <= 0;
      x81325 <= 0;
      x81328 <= 0;
      x81331 <= 0;
      x81334 <= 0;
      x81337 <= 0;
      x81340 <= 0;
      x81343 <= 0;
      x81346 <= 0;
      x81349 <= 0;
      x81352 <= 0;
      x81355 <= 0;
      x81358 <= 0;
      x81361 <= 0;
      x81364 <= 0;
      x81367 <= 0;
      x81370 <= 0;
      x81373 <= 0;
      x81376 <= 0;
      x81379 <= 0;
      x81382 <= 0;
      x81385 <= 0;
      x81388 <= 0;
      x81391 <= 0;
      x81394 <= 0;
      x81397 <= 0;
      x81400 <= 0;
      x81403 <= 0;
      x81406 <= 0;
      x81409 <= 0;
      x81412 <= 0;
      x81415 <= 0;
      x81418 <= 0;
      x81421 <= 0;
      x81424 <= 0;
      x81427 <= 0;
      x81430 <= 0;
      x81433 <= 0;
      x81436 <= 0;
      x81439 <= 0;
      x81442 <= 0;
      x81445 <= 0;
      x81448 <= 0;
      x81451 <= 0;
      x81454 <= 0;
      x81457 <= 0;
      x81460 <= 0;
      x81463 <= 0;
      x81466 <= 0;
      x81469 <= 0;
      x81472 <= 0;
      x81475 <= 0;
      x81478 <= 0;
      x81481 <= 0;
      x81484 <= 0;
      x81487 <= 0;
      x81490 <= 0;
      x81493 <= 0;
      x81496 <= 0;
      x81499 <= 0;
      x81502 <= 0;
      x81505 <= 0;
      x81508 <= 0;
      x81511 <= 0;
      x81514 <= 0;
      x81517 <= 0;
      x81520 <= 0;
      x81523 <= 0;
      x81526 <= 0;
      x81529 <= 0;
      x81532 <= 0;
      x81535 <= 0;
      x81538 <= 0;
      x81541 <= 0;
      x81544 <= 0;
      x81547 <= 0;
      x81550 <= 0;
      x81553 <= 0;
      x81556 <= 0;
      x81559 <= 0;
      x81562 <= 0;
      x81565 <= 0;
      x81568 <= 0;
      x81571 <= 0;
      x81574 <= 0;
      x81577 <= 0;
      x81580 <= 0;
      x81583 <= 0;
      x81586 <= 0;
      x81589 <= 0;
      x81592 <= 0;
      x81595 <= 0;
      x81598 <= 0;
      x81601 <= 0;
      x81604 <= 0;
      x81607 <= 0;
      x81610 <= 0;
      x81613 <= 0;
      x81616 <= 0;
      x81619 <= 0;
      x81622 <= 0;
      x81625 <= 0;
      x81628 <= 0;
      x81631 <= 0;
      x81634 <= 0;
      x81637 <= 0;
      x81640 <= 0;
      x81643 <= 0;
      x81646 <= 0;
      x81649 <= 0;
      x81652 <= 0;
      x81655 <= 0;
      x81658 <= 0;
      x81661 <= 0;
      x81664 <= 0;
      x81667 <= 0;
      x81670 <= 0;
      x81673 <= 0;
      x81676 <= 0;
      x81679 <= 0;
      x81682 <= 0;
      x81685 <= 0;
      x81688 <= 0;
      x81691 <= 0;
      x81694 <= 0;
      x81697 <= 0;
      x81700 <= 0;
      x81703 <= 0;
      x81706 <= 0;
      x81709 <= 0;
      x81712 <= 0;
      x81715 <= 0;
      x81718 <= 0;
      x81721 <= 0;
      x81724 <= 0;
      x81727 <= 0;
      x81730 <= 0;
      x81733 <= 0;
      x81736 <= 0;
      x81739 <= 0;
      x81742 <= 0;
      x81745 <= 0;
      x81748 <= 0;
      x81751 <= 0;
      x81754 <= 0;
      x81757 <= 0;
      x81760 <= 0;
      x81763 <= 0;
      x81766 <= 0;
      x81769 <= 0;
      x81772 <= 0;
      x81775 <= 0;
      x81778 <= 0;
      x81781 <= 0;
      x81784 <= 0;
      x81787 <= 0;
      x81790 <= 0;
      x81793 <= 0;
      x81796 <= 0;
      x81799 <= 0;
      x81802 <= 0;
      x81805 <= 0;
      x81808 <= 0;
      x81811 <= 0;
      x81814 <= 0;
      x81817 <= 0;
      x81820 <= 0;
      x81823 <= 0;
      x81826 <= 0;
      x81829 <= 0;
      x81832 <= 0;
      x81835 <= 0;
      x81838 <= 0;
      x81841 <= 0;
      x81844 <= 0;
      x81847 <= 0;
      x81850 <= 0;
      x81853 <= 0;
      x81856 <= 0;
      x81859 <= 0;
      x81862 <= 0;
      x81865 <= 0;
      x81868 <= 0;
      x81871 <= 0;
      x81874 <= 0;
      x81877 <= 0;
      x81880 <= 0;
      x81883 <= 0;
      x81886 <= 0;
      x81889 <= 0;
      x81892 <= 0;
      x81895 <= 0;
      x81898 <= 0;
      x81901 <= 0;
      x81904 <= 0;
      x81907 <= 0;
      x81910 <= 0;
      x81913 <= 0;
      x81916 <= 0;
      x81919 <= 0;
      x81922 <= 0;
      x81925 <= 0;
      x81928 <= 0;
      x81931 <= 0;
      x81934 <= 0;
      x81937 <= 0;
      x81940 <= 0;
      x81943 <= 0;
      x81946 <= 0;
      x81949 <= 0;
      x81952 <= 0;
      x81955 <= 0;
      x81958 <= 0;
      x81961 <= 0;
      x81964 <= 0;
      x81967 <= 0;
      x81970 <= 0;
      x81973 <= 0;
      x81976 <= 0;
      x81979 <= 0;
      x81982 <= 0;
      x81985 <= 0;
      x81988 <= 0;
      x81991 <= 0;
      x81994 <= 0;
      x81997 <= 0;
      x82000 <= 0;
      x82003 <= 0;
      x82006 <= 0;
      x82009 <= 0;
      x82012 <= 0;
      x82015 <= 0;
      x82018 <= 0;
      x82021 <= 0;
      x82024 <= 0;
      x82027 <= 0;
      x82030 <= 0;
      x82033 <= 0;
      x82036 <= 0;
      x82039 <= 0;
      x82042 <= 0;
      x82045 <= 0;
      x82048 <= 0;
      x82051 <= 0;
      x82054 <= 0;
      x82057 <= 0;
      x82060 <= 0;
      x82063 <= 0;
      x82066 <= 0;
      x82069 <= 0;
      x82072 <= 0;
      x82075 <= 0;
      x82078 <= 0;
      x82081 <= 0;
      x82084 <= 0;
      x82087 <= 0;
      x82090 <= 0;
      x82093 <= 0;
      x82096 <= 0;
      x82099 <= 0;
      x82102 <= 0;
      x82105 <= 0;
      x82108 <= 0;
      x82111 <= 0;
      x82114 <= 0;
      x82117 <= 0;
      x82120 <= 0;
      x82123 <= 0;
      x82126 <= 0;
      x82129 <= 0;
      x82132 <= 0;
      x82135 <= 0;
      x82138 <= 0;
      x82141 <= 0;
      x82144 <= 0;
      x82147 <= 0;
      x82150 <= 0;
      x82153 <= 0;
      x82156 <= 0;
      x82159 <= 0;
      x82162 <= 0;
      x82165 <= 0;
      x82168 <= 0;
      x82171 <= 0;
      x82174 <= 0;
      x82177 <= 0;
      x82180 <= 0;
      x82183 <= 0;
      x82186 <= 0;
      x82189 <= 0;
      x82192 <= 0;
      x82195 <= 0;
      x82198 <= 0;
      x82201 <= 0;
      x82204 <= 0;
      x82207 <= 0;
      x82210 <= 0;
      x82213 <= 0;
      x82216 <= 0;
      x82219 <= 0;
      x82222 <= 0;
      x82225 <= 0;
      x82228 <= 0;
      x82231 <= 0;
      x82234 <= 0;
      x82237 <= 0;
      x82240 <= 0;
      x82243 <= 0;
      x82246 <= 0;
      x82249 <= 0;
      x82252 <= 0;
      x82255 <= 0;
      x82258 <= 0;
      x82261 <= 0;
      x82264 <= 0;
      x82267 <= 0;
      x82270 <= 0;
      x82273 <= 0;
      x82276 <= 0;
      x82279 <= 0;
      x82282 <= 0;
      x82285 <= 0;
      x82288 <= 0;
      x82291 <= 0;
      x82294 <= 0;
      x82297 <= 0;
      x82300 <= 0;
      x82303 <= 0;
      x82306 <= 0;
      x82309 <= 0;
      x82312 <= 0;
      x82315 <= 0;
      x82318 <= 0;
      x82321 <= 0;
      x82324 <= 0;
      x82327 <= 0;
      x82330 <= 0;
      x82333 <= 0;
      x82336 <= 0;
      x82339 <= 0;
      x82342 <= 0;
      x82345 <= 0;
      x82348 <= 0;
      x82351 <= 0;
      x82354 <= 0;
      x82357 <= 0;
      x82360 <= 0;
      x82363 <= 0;
      x82366 <= 0;
      x82369 <= 0;
      x82372 <= 0;
      x82375 <= 0;
      x82378 <= 0;
      x82381 <= 0;
      x82384 <= 0;
      x82387 <= 0;
      x82390 <= 0;
      x82393 <= 0;
      x82396 <= 0;
      x82399 <= 0;
      x82402 <= 0;
      x82405 <= 0;
      x82408 <= 0;
      x82411 <= 0;
      x82414 <= 0;
      x82417 <= 0;
      x82420 <= 0;
      x82423 <= 0;
      x82426 <= 0;
      x82429 <= 0;
      x82432 <= 0;
      x82435 <= 0;
      x82438 <= 0;
      x82441 <= 0;
      x82444 <= 0;
      x82447 <= 0;
      x82450 <= 0;
      x82453 <= 0;
      x82456 <= 0;
      x82459 <= 0;
      x82462 <= 0;
      x82465 <= 0;
      x82468 <= 0;
      x82471 <= 0;
      x82474 <= 0;
      x82477 <= 0;
      x82480 <= 0;
      x82483 <= 0;
      x82486 <= 0;
      x82489 <= 0;
      x82492 <= 0;
      x82495 <= 0;
      x82498 <= 0;
      x82501 <= 0;
      x82504 <= 0;
      x82507 <= 0;
      x82510 <= 0;
      x82513 <= 0;
      x82516 <= 0;
      x82519 <= 0;
      x82522 <= 0;
      x82525 <= 0;
      x82528 <= 0;
      x82531 <= 0;
      x82534 <= 0;
      x82537 <= 0;
      x82540 <= 0;
      x82543 <= 0;
      x82546 <= 0;
      x82549 <= 0;
      x82552 <= 0;
      x82555 <= 0;
      x82558 <= 0;
      x82561 <= 0;
      x82564 <= 0;
      x82567 <= 0;
      x82570 <= 0;
      x82573 <= 0;
      x82576 <= 0;
      x82579 <= 0;
      x82582 <= 0;
      x82585 <= 0;
      x82588 <= 0;
      x82591 <= 0;
      x82594 <= 0;
      x82597 <= 0;
      x82600 <= 0;
      x82603 <= 0;
      x82606 <= 0;
      x82609 <= 0;
      x82612 <= 0;
      x82615 <= 0;
      x82618 <= 0;
      x82621 <= 0;
      x82624 <= 0;
      x82627 <= 0;
      x82630 <= 0;
      x82633 <= 0;
      x82636 <= 0;
      x82639 <= 0;
      x82642 <= 0;
      x82645 <= 0;
      x82648 <= 0;
      x82651 <= 0;
      x82654 <= 0;
      x82657 <= 0;
      x82660 <= 0;
      x82663 <= 0;
      x82666 <= 0;
      x82669 <= 0;
      x82672 <= 0;
      x82675 <= 0;
      x82678 <= 0;
      x82681 <= 0;
      x82684 <= 0;
      x82687 <= 0;
      x82690 <= 0;
      x82693 <= 0;
      x82696 <= 0;
      x82699 <= 0;
      x82702 <= 0;
      x82705 <= 0;
      x82708 <= 0;
      x82711 <= 0;
      x82714 <= 0;
      x82717 <= 0;
      x82720 <= 0;
      x82723 <= 0;
      x82726 <= 0;
      x82729 <= 0;
      x82732 <= 0;
      x82735 <= 0;
      x82738 <= 0;
      x82741 <= 0;
      x82744 <= 0;
      x82747 <= 0;
      x82750 <= 0;
      x82753 <= 0;
      x82756 <= 0;
      x82759 <= 0;
      x82762 <= 0;
      x82765 <= 0;
      x82768 <= 0;
      x82771 <= 0;
      x82774 <= 0;
      x82777 <= 0;
      x82780 <= 0;
      x82783 <= 0;
      x82786 <= 0;
      x82789 <= 0;
      x82792 <= 0;
      x82795 <= 0;
      x82798 <= 0;
      x82801 <= 0;
      x82804 <= 0;
      x82807 <= 0;
      x82810 <= 0;
      x82813 <= 0;
      x82816 <= 0;
      x82819 <= 0;
      x82822 <= 0;
      x82825 <= 0;
      x82828 <= 0;
      x82831 <= 0;
      x82834 <= 0;
      x82837 <= 0;
      x82840 <= 0;
      x82843 <= 0;
      x82846 <= 0;
      x82849 <= 0;
      x82852 <= 0;
      x82855 <= 0;
      x82858 <= 0;
      x82861 <= 0;
      x82864 <= 0;
      x82867 <= 0;
      x82870 <= 0;
      x82873 <= 0;
      x82876 <= 0;
      x82879 <= 0;
      x82882 <= 0;
      x82885 <= 0;
      x82888 <= 0;
      x82891 <= 0;
      x82894 <= 0;
      x82897 <= 0;
      x82900 <= 0;
      x82903 <= 0;
      x82906 <= 0;
      x82909 <= 0;
      x82912 <= 0;
      x82915 <= 0;
      x82918 <= 0;
      x82921 <= 0;
      x82924 <= 0;
      x82927 <= 0;
      x82930 <= 0;
      x82933 <= 0;
      x82936 <= 0;
      x82939 <= 0;
      x82942 <= 0;
      x82945 <= 0;
      x82948 <= 0;
      x82951 <= 0;
      x82954 <= 0;
      x82957 <= 0;
      x82960 <= 0;
      x82963 <= 0;
      x82966 <= 0;
      x82969 <= 0;
      x82972 <= 0;
      x82975 <= 0;
      x82978 <= 0;
      x82981 <= 0;
      x82984 <= 0;
      x82987 <= 0;
      x82990 <= 0;
      x82993 <= 0;
      x82996 <= 0;
      x82999 <= 0;
      x83002 <= 0;
      x83005 <= 0;
      x83008 <= 0;
      x83011 <= 0;
      x83014 <= 0;
      x83017 <= 0;
      x83020 <= 0;
      x83023 <= 0;
      x83026 <= 0;
      x83029 <= 0;
      x83032 <= 0;
      x83035 <= 0;
      x83038 <= 0;
      x83041 <= 0;
      x83044 <= 0;
      x83047 <= 0;
      x83050 <= 0;
      x83053 <= 0;
      x83056 <= 0;
      x83059 <= 0;
      x83062 <= 0;
      x83065 <= 0;
      x83068 <= 0;
      x83071 <= 0;
      x83074 <= 0;
      x83077 <= 0;
      x83080 <= 0;
      x83083 <= 0;
      x83086 <= 0;
      x83089 <= 0;
      x83092 <= 0;
      x83095 <= 0;
      x83098 <= 0;
      x83101 <= 0;
      x83104 <= 0;
      x83107 <= 0;
      x83110 <= 0;
      x83113 <= 0;
      x83116 <= 0;
      x83119 <= 0;
      x83122 <= 0;
      x83125 <= 0;
      x83128 <= 0;
      x83131 <= 0;
      x83134 <= 0;
      x83137 <= 0;
      x83140 <= 0;
      x83143 <= 0;
      x83146 <= 0;
      x83149 <= 0;
      x83152 <= 0;
      x83155 <= 0;
      x83158 <= 0;
      x83161 <= 0;
      x83164 <= 0;
      x83167 <= 0;
      x83170 <= 0;
      x83173 <= 0;
      x83176 <= 0;
      x83179 <= 0;
      x83182 <= 0;
      x83185 <= 0;
      x83188 <= 0;
      x83191 <= 0;
      x83194 <= 0;
      x83197 <= 0;
      x83200 <= 0;
      x83203 <= 0;
      x83206 <= 0;
      x83209 <= 0;
      x83212 <= 0;
      x83215 <= 0;
      x83218 <= 0;
      x83221 <= 0;
      x83224 <= 0;
      x83227 <= 0;
      x83230 <= 0;
      x83233 <= 0;
      x83236 <= 0;
      x83239 <= 0;
      x83242 <= 0;
      x83245 <= 0;
      x83248 <= 0;
      x83251 <= 0;
      x83254 <= 0;
      x83257 <= 0;
      x83260 <= 0;
      x83263 <= 0;
      x83266 <= 0;
      x83269 <= 0;
      x83272 <= 0;
      x83275 <= 0;
      x83278 <= 0;
      x83281 <= 0;
      x83284 <= 0;
      x83287 <= 0;
      x83290 <= 0;
      x83293 <= 0;
      x83296 <= 0;
      x83299 <= 0;
      x83302 <= 0;
      x83305 <= 0;
      x83308 <= 0;
      x83311 <= 0;
      x83314 <= 0;
      x83317 <= 0;
      x83320 <= 0;
      x83323 <= 0;
      x83326 <= 0;
      x83329 <= 0;
      x83332 <= 0;
      x83335 <= 0;
      x83338 <= 0;
      x83341 <= 0;
      x83344 <= 0;
      x83347 <= 0;
      x83352 <= 0;
      x83357 <= 0;
      x83362 <= 0;
      x83367 <= 0;
      x83372 <= 0;
      x83377 <= 0;
      x83382 <= 0;
    end

  always @ (posedge phi)
    begin
       x58 <= x42;
       x59 <= x45;
       x60 <= x48;
       x61 <= x51;
       x62 <= x54;
       x63 <= x57;
       x602 <= x508;
       x603 <= x511;
       x604 <= x514;
       x605 <= x517;
       x606 <= x520;
       x607 <= x523;
       x608 <= x526;
       x609 <= x529;
       x610 <= x532;
       x611 <= x535;
       x612 <= x538;
       x613 <= x541;
       x614 <= x544;
       x615 <= x547;
       x616 <= x550;
       x617 <= x553;
       x618 <= x556;
       x619 <= x559;
       x620 <= x562;
       x621 <= x565;
       x622 <= x568;
       x623 <= x571;
       x624 <= x574;
       x625 <= x577;
       x626 <= x580;
       x627 <= x583;
       x628 <= x586;
       x629 <= x589;
       x630 <= x592;
       x631 <= x595;
       x632 <= x598;
       x633 <= x601;
       x674 <= x664;
       x675 <= x667;
       x676 <= x670;
       x677 <= x673;
       x1232 <= x1231;
       x1238 <= x1237;
       x1244 <= x1243;
       x1250 <= x1249;
       x1256 <= x1255;
       x1262 <= x1261;
       x1268 <= x1267;
       x1274 <= x1273;
       x1281 <= x1280;
       x1288 <= x1287;
       x1294 <= x1293;
       x1300 <= x1299;
       x1306 <= x1305;
       x1312 <= x1311;
       x1318 <= x1317;
       x1324 <= x1323;
       x1330 <= x1329;
       x1336 <= x1335;
       x1342 <= x1341;
       x1348 <= x1347;
       x1354 <= x1353;
       x1360 <= x1359;
       x1366 <= x1365;
       x1372 <= x1371;
       x1379 <= x1378;
       x1386 <= x1385;
       x1392 <= x1391;
       x1398 <= x1397;
       x1404 <= x1403;
       x1410 <= x1409;
       x1416 <= x1415;
       x1422 <= x1421;
       x1758 <= x1757;
       x1768 <= x1767;
       x1778 <= x1777;
       x1788 <= x1787;
       x1798 <= x1797;
       x1808 <= x1807;
       x1818 <= x1817;
       x1828 <= x1827;
       x1914 <= x1913;
       x1918 <= x1917;
       x1922 <= x1921;
       x1926 <= x1925;
       x1930 <= x1929;
       x1934 <= x1933;
       x1940 <= x1939;
       x1944 <= x1943;
       x1948 <= x1947;
       x1952 <= x1951;
       x1956 <= x1955;
       x1960 <= x1959;
       x1966 <= x1965;
       x1970 <= x1969;
       x1974 <= x1973;
       x1978 <= x1977;
       x1982 <= x1981;
       x1986 <= x1985;
       x1992 <= x1991;
       x1996 <= x1995;
       x2000 <= x1999;
       x2004 <= x2003;
       x2008 <= x2007;
       x2012 <= x2011;
       x2018 <= x2017;
       x2022 <= x2021;
       x2026 <= x2025;
       x2030 <= x2029;
       x2034 <= x2033;
       x2038 <= x2037;
       x2044 <= x2043;
       x2048 <= x2047;
       x2052 <= x2051;
       x2056 <= x2055;
       x2060 <= x2059;
       x2064 <= x2063;
       x2070 <= x2069;
       x2074 <= x2073;
       x2078 <= x2077;
       x2082 <= x2081;
       x2086 <= x2085;
       x2090 <= x2089;
       x2096 <= x2095;
       x2100 <= x2099;
       x2104 <= x2103;
       x2108 <= x2107;
       x2112 <= x2111;
       x2116 <= x2115;
       x2317 <= x2316;
       x2321 <= x2320;
       x2325 <= x2324;
       x2329 <= x2328;
       x2333 <= x2332;
       x2337 <= x2336;
       x2341 <= x2340;
       x2345 <= x2344;
       x2349 <= x2348;
       x2353 <= x2352;
       x2357 <= x2356;
       x2361 <= x2360;
       x2365 <= x2364;
       x2369 <= x2368;
       x2373 <= x2372;
       x2377 <= x2376;
       x2381 <= x2380;
       x2385 <= x2384;
       x2389 <= x2388;
       x2393 <= x2392;
       x2397 <= x2396;
       x2401 <= x2400;
       x2405 <= x2404;
       x2409 <= x2408;
       x2413 <= x2412;
       x2417 <= x2416;
       x2421 <= x2420;
       x2425 <= x2424;
       x2429 <= x2428;
       x2433 <= x2432;
       x2437 <= x2436;
       x2441 <= x2440;
       x2447 <= x2446;
       x2451 <= x2450;
       x2455 <= x2454;
       x2459 <= x2458;
       x2463 <= x2462;
       x2467 <= x2466;
       x2471 <= x2470;
       x2475 <= x2474;
       x2479 <= x2478;
       x2483 <= x2482;
       x2487 <= x2486;
       x2491 <= x2490;
       x2495 <= x2494;
       x2499 <= x2498;
       x2503 <= x2502;
       x2507 <= x2506;
       x2511 <= x2510;
       x2515 <= x2514;
       x2519 <= x2518;
       x2523 <= x2522;
       x2527 <= x2526;
       x2531 <= x2530;
       x2535 <= x2534;
       x2539 <= x2538;
       x2543 <= x2542;
       x2547 <= x2546;
       x2551 <= x2550;
       x2555 <= x2554;
       x2559 <= x2558;
       x2563 <= x2562;
       x2567 <= x2566;
       x2571 <= x2570;
       x2577 <= x2576;
       x2581 <= x2580;
       x2585 <= x2584;
       x2589 <= x2588;
       x2593 <= x2592;
       x2597 <= x2596;
       x2601 <= x2600;
       x2605 <= x2604;
       x2609 <= x2608;
       x2613 <= x2612;
       x2617 <= x2616;
       x2621 <= x2620;
       x2625 <= x2624;
       x2629 <= x2628;
       x2633 <= x2632;
       x2637 <= x2636;
       x2641 <= x2640;
       x2645 <= x2644;
       x2649 <= x2648;
       x2653 <= x2652;
       x2657 <= x2656;
       x2661 <= x2660;
       x2665 <= x2664;
       x2669 <= x2668;
       x2673 <= x2672;
       x2677 <= x2676;
       x2681 <= x2680;
       x2685 <= x2684;
       x2689 <= x2688;
       x2693 <= x2692;
       x2697 <= x2696;
       x2701 <= x2700;
       x2707 <= x2706;
       x2711 <= x2710;
       x2715 <= x2714;
       x2719 <= x2718;
       x2723 <= x2722;
       x2727 <= x2726;
       x2731 <= x2730;
       x2735 <= x2734;
       x2739 <= x2738;
       x2743 <= x2742;
       x2747 <= x2746;
       x2751 <= x2750;
       x2755 <= x2754;
       x2759 <= x2758;
       x2763 <= x2762;
       x2767 <= x2766;
       x2771 <= x2770;
       x2775 <= x2774;
       x2779 <= x2778;
       x2783 <= x2782;
       x2787 <= x2786;
       x2791 <= x2790;
       x2795 <= x2794;
       x2799 <= x2798;
       x2803 <= x2802;
       x2807 <= x2806;
       x2811 <= x2810;
       x2815 <= x2814;
       x2819 <= x2818;
       x2823 <= x2822;
       x2827 <= x2826;
       x2831 <= x2830;
       x2837 <= x2836;
       x2841 <= x2840;
       x2845 <= x2844;
       x2849 <= x2848;
       x2853 <= x2852;
       x2857 <= x2856;
       x2861 <= x2860;
       x2865 <= x2864;
       x2869 <= x2868;
       x2873 <= x2872;
       x2877 <= x2876;
       x2881 <= x2880;
       x2885 <= x2884;
       x2889 <= x2888;
       x2893 <= x2892;
       x2897 <= x2896;
       x2901 <= x2900;
       x2905 <= x2904;
       x2909 <= x2908;
       x2913 <= x2912;
       x2917 <= x2916;
       x2921 <= x2920;
       x2925 <= x2924;
       x2929 <= x2928;
       x2933 <= x2932;
       x2937 <= x2936;
       x2941 <= x2940;
       x2945 <= x2944;
       x2949 <= x2948;
       x2953 <= x2952;
       x2957 <= x2956;
       x2961 <= x2960;
       x2967 <= x2966;
       x2971 <= x2970;
       x2975 <= x2974;
       x2979 <= x2978;
       x2983 <= x2982;
       x2987 <= x2986;
       x2991 <= x2990;
       x2995 <= x2994;
       x2999 <= x2998;
       x3003 <= x3002;
       x3007 <= x3006;
       x3011 <= x3010;
       x3015 <= x3014;
       x3019 <= x3018;
       x3023 <= x3022;
       x3027 <= x3026;
       x3031 <= x3030;
       x3035 <= x3034;
       x3039 <= x3038;
       x3043 <= x3042;
       x3047 <= x3046;
       x3051 <= x3050;
       x3055 <= x3054;
       x3059 <= x3058;
       x3063 <= x3062;
       x3067 <= x3066;
       x3071 <= x3070;
       x3075 <= x3074;
       x3079 <= x3078;
       x3083 <= x3082;
       x3087 <= x3086;
       x3091 <= x3090;
       x3097 <= x3096;
       x3101 <= x3100;
       x3105 <= x3104;
       x3109 <= x3108;
       x3113 <= x3112;
       x3117 <= x3116;
       x3121 <= x3120;
       x3125 <= x3124;
       x3129 <= x3128;
       x3133 <= x3132;
       x3137 <= x3136;
       x3141 <= x3140;
       x3145 <= x3144;
       x3149 <= x3148;
       x3153 <= x3152;
       x3157 <= x3156;
       x3161 <= x3160;
       x3165 <= x3164;
       x3169 <= x3168;
       x3173 <= x3172;
       x3177 <= x3176;
       x3181 <= x3180;
       x3185 <= x3184;
       x3189 <= x3188;
       x3193 <= x3192;
       x3197 <= x3196;
       x3201 <= x3200;
       x3205 <= x3204;
       x3209 <= x3208;
       x3213 <= x3212;
       x3217 <= x3216;
       x3221 <= x3220;
       x3227 <= x3226;
       x3231 <= x3230;
       x3235 <= x3234;
       x3239 <= x3238;
       x3243 <= x3242;
       x3247 <= x3246;
       x3251 <= x3250;
       x3255 <= x3254;
       x3259 <= x3258;
       x3263 <= x3262;
       x3267 <= x3266;
       x3271 <= x3270;
       x3275 <= x3274;
       x3279 <= x3278;
       x3283 <= x3282;
       x3287 <= x3286;
       x3291 <= x3290;
       x3295 <= x3294;
       x3299 <= x3298;
       x3303 <= x3302;
       x3307 <= x3306;
       x3311 <= x3310;
       x3315 <= x3314;
       x3319 <= x3318;
       x3323 <= x3322;
       x3327 <= x3326;
       x3331 <= x3330;
       x3335 <= x3334;
       x3339 <= x3338;
       x3343 <= x3342;
       x3347 <= x3346;
       x3351 <= x3350;
       x3358 <= x3357;
       x3363 <= x3362;
       x3367 <= x3366;
       x3371 <= x3370;
       x3375 <= x3374;
       x3379 <= x3378;
       x3383 <= x3382;
       x3387 <= x3386;
       x3391 <= x3390;
       x3395 <= x3394;
       x3399 <= x3398;
       x3403 <= x3402;
       x3407 <= x3406;
       x3411 <= x3410;
       x3415 <= x3414;
       x3419 <= x3418;
       x3423 <= x3422;
       x3427 <= x3426;
       x3431 <= x3430;
       x3435 <= x3434;
       x3439 <= x3438;
       x3443 <= x3442;
       x3447 <= x3446;
       x3451 <= x3450;
       x3455 <= x3454;
       x3459 <= x3458;
       x3463 <= x3462;
       x3467 <= x3466;
       x3471 <= x3470;
       x3475 <= x3474;
       x3479 <= x3478;
       x3483 <= x3482;
       x3489 <= x3488;
       x3493 <= x3492;
       x3497 <= x3496;
       x3501 <= x3500;
       x3505 <= x3504;
       x3509 <= x3508;
       x3513 <= x3512;
       x3517 <= x3516;
       x3521 <= x3520;
       x3525 <= x3524;
       x3529 <= x3528;
       x3533 <= x3532;
       x3537 <= x3536;
       x3541 <= x3540;
       x3545 <= x3544;
       x3549 <= x3548;
       x3553 <= x3552;
       x3557 <= x3556;
       x3561 <= x3560;
       x3565 <= x3564;
       x3569 <= x3568;
       x3573 <= x3572;
       x3577 <= x3576;
       x3581 <= x3580;
       x3585 <= x3584;
       x3589 <= x3588;
       x3593 <= x3592;
       x3597 <= x3596;
       x3601 <= x3600;
       x3605 <= x3604;
       x3609 <= x3608;
       x3613 <= x3612;
       x3619 <= x3618;
       x3623 <= x3622;
       x3627 <= x3626;
       x3631 <= x3630;
       x3635 <= x3634;
       x3639 <= x3638;
       x3643 <= x3642;
       x3647 <= x3646;
       x3651 <= x3650;
       x3655 <= x3654;
       x3659 <= x3658;
       x3663 <= x3662;
       x3667 <= x3666;
       x3671 <= x3670;
       x3675 <= x3674;
       x3679 <= x3678;
       x3683 <= x3682;
       x3687 <= x3686;
       x3691 <= x3690;
       x3695 <= x3694;
       x3699 <= x3698;
       x3703 <= x3702;
       x3707 <= x3706;
       x3711 <= x3710;
       x3715 <= x3714;
       x3719 <= x3718;
       x3723 <= x3722;
       x3727 <= x3726;
       x3731 <= x3730;
       x3735 <= x3734;
       x3739 <= x3738;
       x3743 <= x3742;
       x3749 <= x3748;
       x3753 <= x3752;
       x3757 <= x3756;
       x3761 <= x3760;
       x3765 <= x3764;
       x3769 <= x3768;
       x3773 <= x3772;
       x3777 <= x3776;
       x3781 <= x3780;
       x3785 <= x3784;
       x3789 <= x3788;
       x3793 <= x3792;
       x3797 <= x3796;
       x3801 <= x3800;
       x3805 <= x3804;
       x3809 <= x3808;
       x3813 <= x3812;
       x3817 <= x3816;
       x3821 <= x3820;
       x3825 <= x3824;
       x3829 <= x3828;
       x3833 <= x3832;
       x3837 <= x3836;
       x3841 <= x3840;
       x3845 <= x3844;
       x3849 <= x3848;
       x3853 <= x3852;
       x3857 <= x3856;
       x3861 <= x3860;
       x3865 <= x3864;
       x3869 <= x3868;
       x3873 <= x3872;
       x3879 <= x3878;
       x3883 <= x3882;
       x3887 <= x3886;
       x3891 <= x3890;
       x3895 <= x3894;
       x3899 <= x3898;
       x3903 <= x3902;
       x3907 <= x3906;
       x3911 <= x3910;
       x3915 <= x3914;
       x3919 <= x3918;
       x3923 <= x3922;
       x3927 <= x3926;
       x3931 <= x3930;
       x3935 <= x3934;
       x3939 <= x3938;
       x3943 <= x3942;
       x3947 <= x3946;
       x3951 <= x3950;
       x3955 <= x3954;
       x3959 <= x3958;
       x3963 <= x3962;
       x3967 <= x3966;
       x3971 <= x3970;
       x3975 <= x3974;
       x3979 <= x3978;
       x3983 <= x3982;
       x3987 <= x3986;
       x3991 <= x3990;
       x3995 <= x3994;
       x3999 <= x3998;
       x4003 <= x4002;
       x4009 <= x4008;
       x4013 <= x4012;
       x4017 <= x4016;
       x4021 <= x4020;
       x4025 <= x4024;
       x4029 <= x4028;
       x4033 <= x4032;
       x4037 <= x4036;
       x4041 <= x4040;
       x4045 <= x4044;
       x4049 <= x4048;
       x4053 <= x4052;
       x4057 <= x4056;
       x4061 <= x4060;
       x4065 <= x4064;
       x4069 <= x4068;
       x4073 <= x4072;
       x4077 <= x4076;
       x4081 <= x4080;
       x4085 <= x4084;
       x4089 <= x4088;
       x4093 <= x4092;
       x4097 <= x4096;
       x4101 <= x4100;
       x4105 <= x4104;
       x4109 <= x4108;
       x4113 <= x4112;
       x4117 <= x4116;
       x4121 <= x4120;
       x4125 <= x4124;
       x4129 <= x4128;
       x4133 <= x4132;
       x4139 <= x4138;
       x4143 <= x4142;
       x4147 <= x4146;
       x4151 <= x4150;
       x4155 <= x4154;
       x4159 <= x4158;
       x4163 <= x4162;
       x4167 <= x4166;
       x4171 <= x4170;
       x4175 <= x4174;
       x4179 <= x4178;
       x4183 <= x4182;
       x4187 <= x4186;
       x4191 <= x4190;
       x4195 <= x4194;
       x4199 <= x4198;
       x4203 <= x4202;
       x4207 <= x4206;
       x4211 <= x4210;
       x4215 <= x4214;
       x4219 <= x4218;
       x4223 <= x4222;
       x4227 <= x4226;
       x4231 <= x4230;
       x4235 <= x4234;
       x4239 <= x4238;
       x4243 <= x4242;
       x4247 <= x4246;
       x4251 <= x4250;
       x4255 <= x4254;
       x4259 <= x4258;
       x4263 <= x4262;
       x4269 <= x4268;
       x4273 <= x4272;
       x4277 <= x4276;
       x4281 <= x4280;
       x4285 <= x4284;
       x4289 <= x4288;
       x4293 <= x4292;
       x4297 <= x4296;
       x4301 <= x4300;
       x4305 <= x4304;
       x4309 <= x4308;
       x4313 <= x4312;
       x4317 <= x4316;
       x4321 <= x4320;
       x4325 <= x4324;
       x4329 <= x4328;
       x4333 <= x4332;
       x4337 <= x4336;
       x4341 <= x4340;
       x4345 <= x4344;
       x4349 <= x4348;
       x4353 <= x4352;
       x4357 <= x4356;
       x4361 <= x4360;
       x4365 <= x4364;
       x4369 <= x4368;
       x4373 <= x4372;
       x4377 <= x4376;
       x4381 <= x4380;
       x4385 <= x4384;
       x4389 <= x4388;
       x4393 <= x4392;
       x4399 <= x4398;
       x4404 <= x4403;
       x4409 <= x4408;
       x4413 <= x4412;
       x4417 <= x4416;
       x4421 <= x4420;
       x4425 <= x4424;
       x4429 <= x4428;
       x4433 <= x4432;
       x4437 <= x4436;
       x4441 <= x4440;
       x4445 <= x4444;
       x4449 <= x4448;
       x4453 <= x4452;
       x4457 <= x4456;
       x4461 <= x4460;
       x4465 <= x4464;
       x4469 <= x4468;
       x4473 <= x4472;
       x4477 <= x4476;
       x4481 <= x4480;
       x4485 <= x4484;
       x4489 <= x4488;
       x4493 <= x4492;
       x4497 <= x4496;
       x4501 <= x4500;
       x4505 <= x4504;
       x4509 <= x4508;
       x4513 <= x4512;
       x4517 <= x4516;
       x4521 <= x4520;
       x4525 <= x4524;
       x4531 <= x4530;
       x4535 <= x4534;
       x4539 <= x4538;
       x4543 <= x4542;
       x4547 <= x4546;
       x4551 <= x4550;
       x4555 <= x4554;
       x4559 <= x4558;
       x4563 <= x4562;
       x4567 <= x4566;
       x4571 <= x4570;
       x4575 <= x4574;
       x4579 <= x4578;
       x4583 <= x4582;
       x4587 <= x4586;
       x4591 <= x4590;
       x4595 <= x4594;
       x4599 <= x4598;
       x4603 <= x4602;
       x4607 <= x4606;
       x4611 <= x4610;
       x4615 <= x4614;
       x4619 <= x4618;
       x4623 <= x4622;
       x4627 <= x4626;
       x4631 <= x4630;
       x4635 <= x4634;
       x4639 <= x4638;
       x4643 <= x4642;
       x4647 <= x4646;
       x4651 <= x4650;
       x4655 <= x4654;
       x4661 <= x4660;
       x4665 <= x4664;
       x4669 <= x4668;
       x4673 <= x4672;
       x4677 <= x4676;
       x4681 <= x4680;
       x4685 <= x4684;
       x4689 <= x4688;
       x4693 <= x4692;
       x4697 <= x4696;
       x4701 <= x4700;
       x4705 <= x4704;
       x4709 <= x4708;
       x4713 <= x4712;
       x4717 <= x4716;
       x4721 <= x4720;
       x4725 <= x4724;
       x4729 <= x4728;
       x4733 <= x4732;
       x4737 <= x4736;
       x4741 <= x4740;
       x4745 <= x4744;
       x4749 <= x4748;
       x4753 <= x4752;
       x4757 <= x4756;
       x4761 <= x4760;
       x4765 <= x4764;
       x4769 <= x4768;
       x4773 <= x4772;
       x4777 <= x4776;
       x4781 <= x4780;
       x4785 <= x4784;
       x4791 <= x4790;
       x4795 <= x4794;
       x4799 <= x4798;
       x4803 <= x4802;
       x4807 <= x4806;
       x4811 <= x4810;
       x4815 <= x4814;
       x4819 <= x4818;
       x4823 <= x4822;
       x4827 <= x4826;
       x4831 <= x4830;
       x4835 <= x4834;
       x4839 <= x4838;
       x4843 <= x4842;
       x4847 <= x4846;
       x4851 <= x4850;
       x4855 <= x4854;
       x4859 <= x4858;
       x4863 <= x4862;
       x4867 <= x4866;
       x4871 <= x4870;
       x4875 <= x4874;
       x4879 <= x4878;
       x4883 <= x4882;
       x4887 <= x4886;
       x4891 <= x4890;
       x4895 <= x4894;
       x4899 <= x4898;
       x4903 <= x4902;
       x4907 <= x4906;
       x4911 <= x4910;
       x4915 <= x4914;
       x4921 <= x4920;
       x4925 <= x4924;
       x4929 <= x4928;
       x4933 <= x4932;
       x4937 <= x4936;
       x4941 <= x4940;
       x4945 <= x4944;
       x4949 <= x4948;
       x4953 <= x4952;
       x4957 <= x4956;
       x4961 <= x4960;
       x4965 <= x4964;
       x4969 <= x4968;
       x4973 <= x4972;
       x4977 <= x4976;
       x4981 <= x4980;
       x4985 <= x4984;
       x4989 <= x4988;
       x4993 <= x4992;
       x4997 <= x4996;
       x5001 <= x5000;
       x5005 <= x5004;
       x5009 <= x5008;
       x5013 <= x5012;
       x5017 <= x5016;
       x5021 <= x5020;
       x5025 <= x5024;
       x5029 <= x5028;
       x5033 <= x5032;
       x5037 <= x5036;
       x5041 <= x5040;
       x5045 <= x5044;
       x5051 <= x5050;
       x5055 <= x5054;
       x5059 <= x5058;
       x5063 <= x5062;
       x5067 <= x5066;
       x5071 <= x5070;
       x5075 <= x5074;
       x5079 <= x5078;
       x5083 <= x5082;
       x5087 <= x5086;
       x5091 <= x5090;
       x5095 <= x5094;
       x5099 <= x5098;
       x5103 <= x5102;
       x5107 <= x5106;
       x5111 <= x5110;
       x5115 <= x5114;
       x5119 <= x5118;
       x5123 <= x5122;
       x5127 <= x5126;
       x5131 <= x5130;
       x5135 <= x5134;
       x5139 <= x5138;
       x5143 <= x5142;
       x5147 <= x5146;
       x5151 <= x5150;
       x5155 <= x5154;
       x5159 <= x5158;
       x5163 <= x5162;
       x5167 <= x5166;
       x5171 <= x5170;
       x5175 <= x5174;
       x5181 <= x5180;
       x5185 <= x5184;
       x5189 <= x5188;
       x5193 <= x5192;
       x5197 <= x5196;
       x5201 <= x5200;
       x5205 <= x5204;
       x5209 <= x5208;
       x5213 <= x5212;
       x5217 <= x5216;
       x5221 <= x5220;
       x5225 <= x5224;
       x5229 <= x5228;
       x5233 <= x5232;
       x5237 <= x5236;
       x5241 <= x5240;
       x5245 <= x5244;
       x5249 <= x5248;
       x5253 <= x5252;
       x5257 <= x5256;
       x5261 <= x5260;
       x5265 <= x5264;
       x5269 <= x5268;
       x5273 <= x5272;
       x5277 <= x5276;
       x5281 <= x5280;
       x5285 <= x5284;
       x5289 <= x5288;
       x5293 <= x5292;
       x5297 <= x5296;
       x5301 <= x5300;
       x5305 <= x5304;
       x5311 <= x5310;
       x5315 <= x5314;
       x5319 <= x5318;
       x5323 <= x5322;
       x5327 <= x5326;
       x5331 <= x5330;
       x5335 <= x5334;
       x5339 <= x5338;
       x5343 <= x5342;
       x5347 <= x5346;
       x5351 <= x5350;
       x5355 <= x5354;
       x5359 <= x5358;
       x5363 <= x5362;
       x5367 <= x5366;
       x5371 <= x5370;
       x5375 <= x5374;
       x5379 <= x5378;
       x5383 <= x5382;
       x5387 <= x5386;
       x5391 <= x5390;
       x5395 <= x5394;
       x5399 <= x5398;
       x5403 <= x5402;
       x5407 <= x5406;
       x5411 <= x5410;
       x5415 <= x5414;
       x5419 <= x5418;
       x5423 <= x5422;
       x5427 <= x5426;
       x5431 <= x5430;
       x5435 <= x5434;
       x5442 <= x5441;
       x5448 <= x5447;
       x5453 <= x5452;
       x5457 <= x5456;
       x5461 <= x5460;
       x5465 <= x5464;
       x5469 <= x5468;
       x5473 <= x5472;
       x5477 <= x5476;
       x5481 <= x5480;
       x5485 <= x5484;
       x5489 <= x5488;
       x5493 <= x5492;
       x5497 <= x5496;
       x5501 <= x5500;
       x5505 <= x5504;
       x5509 <= x5508;
       x5513 <= x5512;
       x5517 <= x5516;
       x5521 <= x5520;
       x5525 <= x5524;
       x5529 <= x5528;
       x5533 <= x5532;
       x5537 <= x5536;
       x5541 <= x5540;
       x5545 <= x5544;
       x5549 <= x5548;
       x5553 <= x5552;
       x5557 <= x5556;
       x5561 <= x5560;
       x5565 <= x5564;
       x5569 <= x5568;
       x5575 <= x5574;
       x5579 <= x5578;
       x5583 <= x5582;
       x5587 <= x5586;
       x5591 <= x5590;
       x5595 <= x5594;
       x5599 <= x5598;
       x5603 <= x5602;
       x5607 <= x5606;
       x5611 <= x5610;
       x5615 <= x5614;
       x5619 <= x5618;
       x5623 <= x5622;
       x5627 <= x5626;
       x5631 <= x5630;
       x5635 <= x5634;
       x5639 <= x5638;
       x5643 <= x5642;
       x5647 <= x5646;
       x5651 <= x5650;
       x5655 <= x5654;
       x5659 <= x5658;
       x5663 <= x5662;
       x5667 <= x5666;
       x5671 <= x5670;
       x5675 <= x5674;
       x5679 <= x5678;
       x5683 <= x5682;
       x5687 <= x5686;
       x5691 <= x5690;
       x5695 <= x5694;
       x5699 <= x5698;
       x5705 <= x5704;
       x5709 <= x5708;
       x5713 <= x5712;
       x5717 <= x5716;
       x5721 <= x5720;
       x5725 <= x5724;
       x5729 <= x5728;
       x5733 <= x5732;
       x5737 <= x5736;
       x5741 <= x5740;
       x5745 <= x5744;
       x5749 <= x5748;
       x5753 <= x5752;
       x5757 <= x5756;
       x5761 <= x5760;
       x5765 <= x5764;
       x5769 <= x5768;
       x5773 <= x5772;
       x5777 <= x5776;
       x5781 <= x5780;
       x5785 <= x5784;
       x5789 <= x5788;
       x5793 <= x5792;
       x5797 <= x5796;
       x5801 <= x5800;
       x5805 <= x5804;
       x5809 <= x5808;
       x5813 <= x5812;
       x5817 <= x5816;
       x5821 <= x5820;
       x5825 <= x5824;
       x5829 <= x5828;
       x5835 <= x5834;
       x5839 <= x5838;
       x5843 <= x5842;
       x5847 <= x5846;
       x5851 <= x5850;
       x5855 <= x5854;
       x5859 <= x5858;
       x5863 <= x5862;
       x5867 <= x5866;
       x5871 <= x5870;
       x5875 <= x5874;
       x5879 <= x5878;
       x5883 <= x5882;
       x5887 <= x5886;
       x5891 <= x5890;
       x5895 <= x5894;
       x5899 <= x5898;
       x5903 <= x5902;
       x5907 <= x5906;
       x5911 <= x5910;
       x5915 <= x5914;
       x5919 <= x5918;
       x5923 <= x5922;
       x5927 <= x5926;
       x5931 <= x5930;
       x5935 <= x5934;
       x5939 <= x5938;
       x5943 <= x5942;
       x5947 <= x5946;
       x5951 <= x5950;
       x5955 <= x5954;
       x5959 <= x5958;
       x5965 <= x5964;
       x5969 <= x5968;
       x5973 <= x5972;
       x5977 <= x5976;
       x5981 <= x5980;
       x5985 <= x5984;
       x5989 <= x5988;
       x5993 <= x5992;
       x5997 <= x5996;
       x6001 <= x6000;
       x6005 <= x6004;
       x6009 <= x6008;
       x6013 <= x6012;
       x6017 <= x6016;
       x6021 <= x6020;
       x6025 <= x6024;
       x6029 <= x6028;
       x6033 <= x6032;
       x6037 <= x6036;
       x6041 <= x6040;
       x6045 <= x6044;
       x6049 <= x6048;
       x6053 <= x6052;
       x6057 <= x6056;
       x6061 <= x6060;
       x6065 <= x6064;
       x6069 <= x6068;
       x6073 <= x6072;
       x6077 <= x6076;
       x6081 <= x6080;
       x6085 <= x6084;
       x6089 <= x6088;
       x6095 <= x6094;
       x6099 <= x6098;
       x6103 <= x6102;
       x6107 <= x6106;
       x6111 <= x6110;
       x6115 <= x6114;
       x6119 <= x6118;
       x6123 <= x6122;
       x6127 <= x6126;
       x6131 <= x6130;
       x6135 <= x6134;
       x6139 <= x6138;
       x6143 <= x6142;
       x6147 <= x6146;
       x6151 <= x6150;
       x6155 <= x6154;
       x6159 <= x6158;
       x6163 <= x6162;
       x6167 <= x6166;
       x6171 <= x6170;
       x6175 <= x6174;
       x6179 <= x6178;
       x6183 <= x6182;
       x6187 <= x6186;
       x6191 <= x6190;
       x6195 <= x6194;
       x6199 <= x6198;
       x6203 <= x6202;
       x6207 <= x6206;
       x6211 <= x6210;
       x6215 <= x6214;
       x6219 <= x6218;
       x6225 <= x6224;
       x6229 <= x6228;
       x6233 <= x6232;
       x6237 <= x6236;
       x6241 <= x6240;
       x6245 <= x6244;
       x6249 <= x6248;
       x6253 <= x6252;
       x6257 <= x6256;
       x6261 <= x6260;
       x6265 <= x6264;
       x6269 <= x6268;
       x6273 <= x6272;
       x6277 <= x6276;
       x6281 <= x6280;
       x6285 <= x6284;
       x6289 <= x6288;
       x6293 <= x6292;
       x6297 <= x6296;
       x6301 <= x6300;
       x6305 <= x6304;
       x6309 <= x6308;
       x6313 <= x6312;
       x6317 <= x6316;
       x6321 <= x6320;
       x6325 <= x6324;
       x6329 <= x6328;
       x6333 <= x6332;
       x6337 <= x6336;
       x6341 <= x6340;
       x6345 <= x6344;
       x6349 <= x6348;
       x6355 <= x6354;
       x6359 <= x6358;
       x6363 <= x6362;
       x6367 <= x6366;
       x6371 <= x6370;
       x6375 <= x6374;
       x6379 <= x6378;
       x6383 <= x6382;
       x6387 <= x6386;
       x6391 <= x6390;
       x6395 <= x6394;
       x6399 <= x6398;
       x6403 <= x6402;
       x6407 <= x6406;
       x6411 <= x6410;
       x6415 <= x6414;
       x6419 <= x6418;
       x6423 <= x6422;
       x6427 <= x6426;
       x6431 <= x6430;
       x6435 <= x6434;
       x6439 <= x6438;
       x6443 <= x6442;
       x6447 <= x6446;
       x6451 <= x6450;
       x6455 <= x6454;
       x6459 <= x6458;
       x6463 <= x6462;
       x6467 <= x6466;
       x6471 <= x6470;
       x6475 <= x6474;
       x6479 <= x6478;
       x14598 <= x14597;
       x14608 <= x14607;
       x14618 <= x14617;
       x14628 <= x14627;
       x14638 <= x14637;
       x14648 <= x14647;
       x14658 <= x14657;
       x14668 <= x14667;
       x14767 <= x14766;
       x14771 <= x14770;
       x14775 <= x14774;
       x14779 <= x14778;
       x14783 <= x14782;
       x14787 <= x14786;
       x14793 <= x14792;
       x14797 <= x14796;
       x14801 <= x14800;
       x14805 <= x14804;
       x14809 <= x14808;
       x14813 <= x14812;
       x14819 <= x14818;
       x14823 <= x14822;
       x14827 <= x14826;
       x14831 <= x14830;
       x14835 <= x14834;
       x14839 <= x14838;
       x14845 <= x14844;
       x14849 <= x14848;
       x14853 <= x14852;
       x14857 <= x14856;
       x14861 <= x14860;
       x14865 <= x14864;
       x14871 <= x14870;
       x14875 <= x14874;
       x14879 <= x14878;
       x14883 <= x14882;
       x14887 <= x14886;
       x14891 <= x14890;
       x14897 <= x14896;
       x14901 <= x14900;
       x14905 <= x14904;
       x14909 <= x14908;
       x14913 <= x14912;
       x14917 <= x14916;
       x14923 <= x14922;
       x14927 <= x14926;
       x14931 <= x14930;
       x14935 <= x14934;
       x14939 <= x14938;
       x14943 <= x14942;
       x14949 <= x14948;
       x14953 <= x14952;
       x14957 <= x14956;
       x14961 <= x14960;
       x14965 <= x14964;
       x14969 <= x14968;
       x27755 <= x27754;
       x27759 <= x27758;
       x27763 <= x27762;
       x27767 <= x27766;
       x27771 <= x27770;
       x27775 <= x27774;
       x27779 <= x27778;
       x27783 <= x27782;
       x27787 <= x27786;
       x27791 <= x27790;
       x27795 <= x27794;
       x27799 <= x27798;
       x27803 <= x27802;
       x27807 <= x27806;
       x27811 <= x27810;
       x27815 <= x27814;
       x27819 <= x27818;
       x27823 <= x27822;
       x27827 <= x27826;
       x27831 <= x27830;
       x27835 <= x27834;
       x27839 <= x27838;
       x27843 <= x27842;
       x27847 <= x27846;
       x27851 <= x27850;
       x27855 <= x27854;
       x27859 <= x27858;
       x27863 <= x27862;
       x27867 <= x27866;
       x27871 <= x27870;
       x27875 <= x27874;
       x27879 <= x27878;
       x38722 <= x38721;
       x38726 <= x38725;
       x38730 <= x38729;
       x38734 <= x38733;
       x38738 <= x38737;
       x38742 <= x38741;
       x38746 <= x38745;
       x38750 <= x38749;
       x38754 <= x38753;
       x38758 <= x38757;
       x38762 <= x38761;
       x38766 <= x38765;
       x38770 <= x38769;
       x38774 <= x38773;
       x38778 <= x38777;
       x38782 <= x38781;
       x38786 <= x38785;
       x38790 <= x38789;
       x38794 <= x38793;
       x38798 <= x38797;
       x38802 <= x38801;
       x38806 <= x38805;
       x38810 <= x38809;
       x38814 <= x38813;
       x38818 <= x38817;
       x38822 <= x38821;
       x38826 <= x38825;
       x38830 <= x38829;
       x38834 <= x38833;
       x38838 <= x38837;
       x38842 <= x38841;
       x38846 <= x38845;
       x49689 <= x49688;
       x49693 <= x49692;
       x49697 <= x49696;
       x49701 <= x49700;
       x49705 <= x49704;
       x49709 <= x49708;
       x49713 <= x49712;
       x49717 <= x49716;
       x49721 <= x49720;
       x49725 <= x49724;
       x49729 <= x49728;
       x49733 <= x49732;
       x49737 <= x49736;
       x49741 <= x49740;
       x49745 <= x49744;
       x49749 <= x49748;
       x49753 <= x49752;
       x49757 <= x49756;
       x49761 <= x49760;
       x49765 <= x49764;
       x49769 <= x49768;
       x49773 <= x49772;
       x49777 <= x49776;
       x49781 <= x49780;
       x49785 <= x49784;
       x49789 <= x49788;
       x49793 <= x49792;
       x49797 <= x49796;
       x49801 <= x49800;
       x49805 <= x49804;
       x49809 <= x49808;
       x49813 <= x49812;
       x60656 <= x60655;
       x60660 <= x60659;
       x60664 <= x60663;
       x60668 <= x60667;
       x60672 <= x60671;
       x60676 <= x60675;
       x60680 <= x60679;
       x60684 <= x60683;
       x60688 <= x60687;
       x60692 <= x60691;
       x60696 <= x60695;
       x60700 <= x60699;
       x60704 <= x60703;
       x60708 <= x60707;
       x60712 <= x60711;
       x60716 <= x60715;
       x60720 <= x60719;
       x60724 <= x60723;
       x60728 <= x60727;
       x60732 <= x60731;
       x60736 <= x60735;
       x60740 <= x60739;
       x60744 <= x60743;
       x60748 <= x60747;
       x60752 <= x60751;
       x60756 <= x60755;
       x60760 <= x60759;
       x60764 <= x60763;
       x60768 <= x60767;
       x60772 <= x60771;
       x60776 <= x60775;
       x60780 <= x60779;
       x60784 <= x60783;
       x60788 <= x60787;
       x60792 <= x60791;
       x60796 <= x60795;
       x60800 <= x60799;
       x60804 <= x60803;
       x60808 <= x60807;
       x60812 <= x60811;
       x60816 <= x60815;
       x60820 <= x60819;
       x60824 <= x60823;
       x60828 <= x60827;
       x60832 <= x60831;
       x60836 <= x60835;
       x60840 <= x60839;
       x60976 <= x60975;
       x61105 <= x61104;
       x61234 <= x61233;
       x61363 <= x61362;
       x61367 <= x61366;
       x61371 <= x61370;
       x61375 <= x61374;
       x61379 <= x61378;
       x61383 <= x61382;
       x61387 <= x61386;
       x61391 <= x61390;
       x61395 <= x61394;
       x61399 <= x61398;
       x61403 <= x61402;
       x61407 <= x61406;
       x61411 <= x61410;
       x61415 <= x61414;
       x61419 <= x61418;
       x61423 <= x61422;
       x61981 <= x61980;
       x61988 <= x61987;
       x61995 <= x61994;
       x62002 <= x62001;
       x62009 <= x62008;
       x62016 <= x62015;
       x62023 <= x62022;
       x62030 <= x62029;
       x62037 <= x62036;
       x62044 <= x62043;
       x62051 <= x62050;
       x62058 <= x62057;
       x62065 <= x62064;
       x62072 <= x62071;
       x62079 <= x62078;
       x62086 <= x62085;
       x62093 <= x62092;
       x62100 <= x62099;
       x62107 <= x62106;
       x62114 <= x62113;
       x62121 <= x62120;
       x62128 <= x62127;
       x62135 <= x62134;
       x62142 <= x62141;
       x62149 <= x62148;
       x62156 <= x62155;
       x62163 <= x62162;
       x62170 <= x62169;
       x62177 <= x62176;
       x62184 <= x62183;
       x62191 <= x62190;
       x62198 <= x62197;
       x62205 <= x62204;
       x62212 <= x62211;
       x62219 <= x62218;
       x62226 <= x62225;
       x62233 <= x62232;
       x62240 <= x62239;
       x62247 <= x62246;
       x62254 <= x62253;
       x62261 <= x62260;
       x62268 <= x62267;
       x62275 <= x62274;
       x62282 <= x62281;
       x62289 <= x62288;
       x62296 <= x62295;
       x62303 <= x62302;
       x62310 <= x62309;
       x62317 <= x62316;
       x62324 <= x62323;
       x62331 <= x62330;
       x62338 <= x62337;
       x62345 <= x62344;
       x62352 <= x62351;
       x62359 <= x62358;
       x62366 <= x62365;
       x62373 <= x62372;
       x62380 <= x62379;
       x62387 <= x62386;
       x62394 <= x62393;
       x62401 <= x62400;
       x62408 <= x62407;
       x62415 <= x62414;
       x62422 <= x62421;
       x62429 <= x62428;
       x62436 <= x62435;
       x62443 <= x62442;
       x62450 <= x62449;
       x62457 <= x62456;
       x62464 <= x62463;
       x62471 <= x62470;
       x62478 <= x62477;
       x62485 <= x62484;
       x62492 <= x62491;
       x62499 <= x62498;
       x62506 <= x62505;
       x62513 <= x62512;
       x62520 <= x62519;
       x62527 <= x62526;
       x62534 <= x62533;
       x62541 <= x62540;
       x62548 <= x62547;
       x62555 <= x62554;
       x62562 <= x62561;
       x62569 <= x62568;
       x62576 <= x62575;
       x62583 <= x62582;
       x62590 <= x62589;
       x62597 <= x62596;
       x62604 <= x62603;
       x62611 <= x62610;
       x62618 <= x62617;
       x62625 <= x62624;
       x62632 <= x62631;
       x62639 <= x62638;
       x62646 <= x62645;
       x62653 <= x62652;
       x62660 <= x62659;
       x62667 <= x62666;
       x62674 <= x62673;
       x62681 <= x62680;
       x62688 <= x62687;
       x62695 <= x62694;
       x62702 <= x62701;
       x62709 <= x62708;
       x62716 <= x62715;
       x62723 <= x62722;
       x62730 <= x62729;
       x62737 <= x62736;
       x62744 <= x62743;
       x62751 <= x62750;
       x62758 <= x62757;
       x62765 <= x62764;
       x62772 <= x62771;
       x62779 <= x62778;
       x62786 <= x62785;
       x62793 <= x62792;
       x62800 <= x62799;
       x62807 <= x62806;
       x62814 <= x62813;
       x62821 <= x62820;
       x62828 <= x62827;
       x62835 <= x62834;
       x62842 <= x62841;
       x62849 <= x62848;
       x62856 <= x62855;
       x62863 <= x62862;
       x62870 <= x62869;
       x62873 <= x86263;
       x62877 <= x62876;
       x62881 <= x62880;
       x62885 <= x62884;
       x62889 <= x62888;
       x62893 <= x62892;
       x62897 <= x62896;
       x62901 <= x62900;
       x62905 <= x62904;
       x62909 <= x62908;
       x62913 <= x62912;
       x62917 <= x62916;
       x62921 <= x62920;
       x62925 <= x62924;
       x62929 <= x62928;
       x63908 <= x87265;
       x63909 <= x87265;
       x63910 <= x87265;
       x63911 <= x86264;
       x63912 <= x86265;
       x64640 <= x87265;
       x64641 <= x87265;
       x64642 <= x87265;
       x64643 <= x86297;
       x64644 <= x86298;
       x65310 <= x87265;
       x65311 <= x87265;
       x65312 <= x87265;
       x65313 <= x86330;
       x65314 <= x86331;
       x65980 <= x87265;
       x65981 <= x87265;
       x65982 <= x87265;
       x65983 <= x86363;
       x65984 <= x86364;
       x66413 <= x66412;
       x66417 <= x66416;
       x66421 <= x66420;
       x66425 <= x66424;
       x66429 <= x66428;
       x66433 <= x66432;
       x66437 <= x66436;
       x66441 <= x66440;
       x66445 <= x66444;
       x66449 <= x66448;
       x66453 <= x66452;
       x66457 <= x66456;
       x66461 <= x66460;
       x66465 <= x66464;
       x66469 <= x66468;
       x66894 <= x66893;
       x66898 <= x66897;
       x66902 <= x66901;
       x66906 <= x66905;
       x66910 <= x66909;
       x66914 <= x66913;
       x66918 <= x66917;
       x66922 <= x66921;
       x66926 <= x66925;
       x66930 <= x66929;
       x66934 <= x66933;
       x66938 <= x66937;
       x66942 <= x66941;
       x66946 <= x66945;
       x66950 <= x66949;
       x66954 <= x66953;
       x66958 <= x66957;
       x66962 <= x66961;
       x66966 <= x66965;
       x66970 <= x66969;
       x66974 <= x66973;
       x66978 <= x66977;
       x66982 <= x66981;
       x66986 <= x66985;
       x66990 <= x66989;
       x66994 <= x66993;
       x66998 <= x66997;
       x67002 <= x67001;
       x67006 <= x67005;
       x67010 <= x67009;
       x67014 <= x67013;
       x67018 <= x67017;
       x67022 <= x67021;
       x67026 <= x67025;
       x67030 <= x67029;
       x67034 <= x67033;
       x67038 <= x67037;
       x67042 <= x67041;
       x67046 <= x67045;
       x67050 <= x67049;
       x67054 <= x67053;
       x67058 <= x67057;
       x67062 <= x67061;
       x67066 <= x67065;
       x67070 <= x67069;
       x67074 <= x67073;
       x67078 <= x67077;
       x67082 <= x67081;
       x67086 <= x67085;
       x67090 <= x67089;
       x67094 <= x67093;
       x67098 <= x67097;
       x67102 <= x67101;
       x67106 <= x67105;
       x67110 <= x67109;
       x67114 <= x67113;
       x67118 <= x67117;
       x67122 <= x67121;
       x67126 <= x67125;
       x67130 <= x67129;
       x67134 <= x67133;
       x67138 <= x67137;
       x67142 <= x67141;
       x67146 <= x67145;
       x67150 <= x67149;
       x67154 <= x67153;
       x67158 <= x67157;
       x67162 <= x67161;
       x67166 <= x67165;
       x67170 <= x67169;
       x67174 <= x67173;
       x67178 <= x67177;
       x67182 <= x67181;
       x67186 <= x67185;
       x67190 <= x67189;
       x67194 <= x67193;
       x67198 <= x67197;
       x67202 <= x67201;
       x67206 <= x67205;
       x67210 <= x67209;
       x67214 <= x67213;
       x67218 <= x67217;
       x67222 <= x67221;
       x67226 <= x67225;
       x67230 <= x67229;
       x67234 <= x67233;
       x67238 <= x67237;
       x67242 <= x67241;
       x67246 <= x67245;
       x67250 <= x67249;
       x67254 <= x67253;
       x67258 <= x67257;
       x67262 <= x67261;
       x67266 <= x67265;
       x67270 <= x67269;
       x67274 <= x67273;
       x67278 <= x67277;
       x67282 <= x67281;
       x67286 <= x67285;
       x67290 <= x67289;
       x67294 <= x67293;
       x67298 <= x67297;
       x67302 <= x67301;
       x67306 <= x67305;
       x67310 <= x67309;
       x67314 <= x67313;
       x67318 <= x67317;
       x67322 <= x67321;
       x67326 <= x67325;
       x67330 <= x67329;
       x67334 <= x67333;
       x67338 <= x67337;
       x67342 <= x67341;
       x67346 <= x67345;
       x67350 <= x67349;
       x67354 <= x67353;
       x67358 <= x67357;
       x67362 <= x67361;
       x67366 <= x67365;
       x67370 <= x67369;
       x67374 <= x67373;
       x67378 <= x67377;
       x67382 <= x67381;
       x67386 <= x67385;
       x67390 <= x67389;
       x67394 <= x67393;
       x67398 <= x67397;
       x67402 <= x67401;
       x67405 <= x86396;
       x67409 <= x67408;
       x67413 <= x67412;
       x67417 <= x67416;
       x67421 <= x67420;
       x67425 <= x67424;
       x67429 <= x67428;
       x67433 <= x67432;
       x67437 <= x67436;
       x67441 <= x67440;
       x67445 <= x67444;
       x67449 <= x67448;
       x67453 <= x67452;
       x67457 <= x67456;
       x67461 <= x67460;
       x67887 <= x67886;
       x67891 <= x67890;
       x67895 <= x67894;
       x67899 <= x67898;
       x67903 <= x67902;
       x67907 <= x67906;
       x67911 <= x67910;
       x67915 <= x67914;
       x67919 <= x67918;
       x67923 <= x67922;
       x67927 <= x67926;
       x67931 <= x67930;
       x67935 <= x67934;
       x67939 <= x67938;
       x67943 <= x67942;
       x67947 <= x67946;
       x67951 <= x67950;
       x67955 <= x67954;
       x67959 <= x67958;
       x67963 <= x67962;
       x67967 <= x67966;
       x67971 <= x67970;
       x67975 <= x67974;
       x67979 <= x67978;
       x67983 <= x67982;
       x67987 <= x67986;
       x67991 <= x67990;
       x67995 <= x67994;
       x67999 <= x67998;
       x68003 <= x68002;
       x68007 <= x68006;
       x68011 <= x68010;
       x68015 <= x68014;
       x68019 <= x68018;
       x68023 <= x68022;
       x68027 <= x68026;
       x68031 <= x68030;
       x68035 <= x68034;
       x68039 <= x68038;
       x68043 <= x68042;
       x68047 <= x68046;
       x68051 <= x68050;
       x68055 <= x68054;
       x68059 <= x68058;
       x68063 <= x68062;
       x68067 <= x68066;
       x68071 <= x68070;
       x68075 <= x68074;
       x68079 <= x68078;
       x68083 <= x68082;
       x68087 <= x68086;
       x68091 <= x68090;
       x68095 <= x68094;
       x68099 <= x68098;
       x68103 <= x68102;
       x68107 <= x68106;
       x68111 <= x68110;
       x68115 <= x68114;
       x68119 <= x68118;
       x68123 <= x68122;
       x68127 <= x68126;
       x68131 <= x68130;
       x68135 <= x68134;
       x68139 <= x68138;
       x68143 <= x68142;
       x68147 <= x68146;
       x68151 <= x68150;
       x68155 <= x68154;
       x68159 <= x68158;
       x68163 <= x68162;
       x68167 <= x68166;
       x68171 <= x68170;
       x68175 <= x68174;
       x68179 <= x68178;
       x68183 <= x68182;
       x68187 <= x68186;
       x68191 <= x68190;
       x68195 <= x68194;
       x68199 <= x68198;
       x68203 <= x68202;
       x68207 <= x68206;
       x68211 <= x68210;
       x68215 <= x68214;
       x68219 <= x68218;
       x68223 <= x68222;
       x68227 <= x68226;
       x68231 <= x68230;
       x68235 <= x68234;
       x68239 <= x68238;
       x68243 <= x68242;
       x68247 <= x68246;
       x68251 <= x68250;
       x68255 <= x68254;
       x68259 <= x68258;
       x68263 <= x68262;
       x68267 <= x68266;
       x68271 <= x68270;
       x68275 <= x68274;
       x68279 <= x68278;
       x68283 <= x68282;
       x68287 <= x68286;
       x68291 <= x68290;
       x68295 <= x68294;
       x68299 <= x68298;
       x68303 <= x68302;
       x68307 <= x68306;
       x68311 <= x68310;
       x68315 <= x68314;
       x68319 <= x68318;
       x68323 <= x68322;
       x68327 <= x68326;
       x68331 <= x68330;
       x68335 <= x68334;
       x68339 <= x68338;
       x68343 <= x68342;
       x68347 <= x68346;
       x68351 <= x68350;
       x68355 <= x68354;
       x68359 <= x68358;
       x68363 <= x68362;
       x68367 <= x68366;
       x68371 <= x68370;
       x68375 <= x68374;
       x68379 <= x68378;
       x68383 <= x68382;
       x68387 <= x68386;
       x68391 <= x68390;
       x68395 <= x68394;
       x68398 <= x86397;
       x68402 <= x68401;
       x68406 <= x68405;
       x68410 <= x68409;
       x68414 <= x68413;
       x68418 <= x68417;
       x68422 <= x68421;
       x68426 <= x68425;
       x68430 <= x68429;
       x68434 <= x68433;
       x68438 <= x68437;
       x68442 <= x68441;
       x68446 <= x68445;
       x68450 <= x68449;
       x68454 <= x68453;
       x68618 <= x68572;
       x68619 <= x68581;
       x68620 <= x68590;
       x68621 <= x68599;
       x68622 <= x68608;
       x68623 <= x68617;
       x71147 <= x71146;
       x71152 <= x71151;
       x71157 <= x71156;
       x71162 <= x71161;
       x71167 <= x71166;
       x71172 <= x71171;
       x71177 <= x71176;
       x71182 <= x71181;
       x71185 <= x71184;
       x71188 <= x71187;
       x71191 <= x71190;
       x71194 <= x71193;
       x71197 <= x71196;
       x71202 <= x71201;
       x71205 <= x71204;
       x71210 <= x71209;
       x71215 <= x71214;
       x71220 <= x71219;
       x71225 <= x71224;
       x71230 <= x71229;
       x71235 <= x71234;
       x71240 <= x71239;
       x71245 <= x71244;
       x71250 <= x71249;
       x71255 <= x71254;
       x71260 <= x71259;
       x71265 <= x71264;
       x71270 <= x71269;
       x71275 <= x71274;
       x71277 <= x86719;
       x71279 <= x86720;
       x71284 <= x71283;
       x71289 <= x71288;
       x71294 <= x71293;
       x71299 <= x71298;
       x71304 <= x71303;
       x71309 <= x71308;
       x71314 <= x71313;
       x71319 <= x71318;
       x71324 <= x71323;
       x71329 <= x71328;
       x71334 <= x71333;
       x71339 <= x71338;
       x71344 <= x71343;
       x71349 <= x71348;
       x71354 <= x71353;
       x71359 <= x71358;
       x71364 <= x71363;
       x71369 <= x71368;
       x71374 <= x71373;
       x71379 <= x71378;
       x71384 <= x71383;
       x71389 <= x71388;
       x71394 <= x71393;
       x71399 <= x71398;
       x71404 <= x71403;
       x71409 <= x71408;
       x71414 <= x71413;
       x71419 <= x71418;
       x71424 <= x71423;
       x71429 <= x71428;
       x71434 <= x71433;
       x71439 <= x71438;
       x71444 <= x71443;
       x71449 <= x71448;
       x71454 <= x71453;
       x71459 <= x71458;
       x71464 <= x71463;
       x71469 <= x71468;
       x71474 <= x71473;
       x71479 <= x71478;
       x71482 <= x71481;
       x71485 <= x71484;
       x71490 <= x71489;
       x71495 <= x71494;
       x71500 <= x71499;
       x71505 <= x71504;
       x71510 <= x71509;
       x71515 <= x71514;
       x71520 <= x71519;
       x71525 <= x71524;
       x71530 <= x71529;
       x71535 <= x71534;
       x71540 <= x71539;
       x71545 <= x71544;
       x71550 <= x71549;
       x71555 <= x71554;
       x71560 <= x71559;
       x71565 <= x71564;
       x71570 <= x71569;
       x71575 <= x71574;
       x71580 <= x71579;
       x71585 <= x71584;
       x71590 <= x71589;
       x71595 <= x71594;
       x71600 <= x71599;
       x71605 <= x71604;
       x71610 <= x71609;
       x71615 <= x71614;
       x71620 <= x71619;
       x71625 <= x71624;
       x71630 <= x71629;
       x71635 <= x71634;
       x71642 <= x71641;
       x71647 <= x71646;
       x71652 <= x71651;
       x71657 <= x71656;
       x71662 <= x71661;
       x71667 <= x71666;
       x71672 <= x71671;
       x71677 <= x71676;
       x71682 <= x71681;
       x71687 <= x71686;
       x71692 <= x71691;
       x71697 <= x71696;
       x71702 <= x71701;
       x71707 <= x71706;
       x71712 <= x71711;
       x71717 <= x71716;
       x71722 <= x71721;
       x71727 <= x71726;
       x71732 <= x71731;
       x71737 <= x71736;
       x71742 <= x71741;
       x71747 <= x71746;
       x71752 <= x71751;
       x71757 <= x71756;
       x71762 <= x71761;
       x71767 <= x71766;
       x71772 <= x71771;
       x71777 <= x71776;
       x71782 <= x71781;
       x71787 <= x71786;
       x71792 <= x71791;
       x71797 <= x71796;
       x71802 <= x71801;
       x71807 <= x71806;
       x71812 <= x71811;
       x71817 <= x71816;
       x71822 <= x71821;
       x71827 <= x71826;
       x71832 <= x71831;
       x71837 <= x71836;
       x71842 <= x71841;
       x71847 <= x71846;
       x71852 <= x71851;
       x71857 <= x71856;
       x71862 <= x71861;
       x71867 <= x71866;
       x71872 <= x71871;
       x71877 <= x71876;
       x71882 <= x71881;
       x71887 <= x71886;
       x71892 <= x71891;
       x71897 <= x71896;
       x71902 <= x71901;
       x71907 <= x71906;
       x71910 <= x71909;
       x71913 <= x71912;
       x71916 <= x71915;
       x71919 <= x71918;
       x71922 <= x71921;
       x71925 <= x71924;
       x71928 <= x71927;
       x71931 <= x71930;
       x71934 <= x71933;
       x71937 <= x71936;
       x71942 <= x71941;
       x71947 <= x71946;
       x71952 <= x71951;
       x71957 <= x71956;
       x71962 <= x71961;
       x71967 <= x71966;
       x71972 <= x71971;
       x71977 <= x71976;
       x71982 <= x71981;
       x71987 <= x71986;
       x71992 <= x71991;
       x71997 <= x71996;
       x72002 <= x72001;
       x72007 <= x72006;
       x72012 <= x72011;
       x72017 <= x72016;
       x72022 <= x72021;
       x72027 <= x72026;
       x72032 <= x72031;
       x72037 <= x72036;
       x72042 <= x72041;
       x72047 <= x72046;
       x72052 <= x72051;
       x72057 <= x72056;
       x72062 <= x72061;
       x72067 <= x72066;
       x72072 <= x72071;
       x72077 <= x72076;
       x72082 <= x72081;
       x72087 <= x72086;
       x72092 <= x72091;
       x72097 <= x72096;
       x72102 <= x72101;
       x72107 <= x72106;
       x72112 <= x72111;
       x72117 <= x72116;
       x72122 <= x72121;
       x72127 <= x72126;
       x72132 <= x72131;
       x72137 <= x72136;
       x72142 <= x72141;
       x72147 <= x72146;
       x72152 <= x72151;
       x72157 <= x72156;
       x72162 <= x72161;
       x72167 <= x72166;
       x72172 <= x72171;
       x72177 <= x72176;
       x72182 <= x72181;
       x72187 <= x72186;
       x72192 <= x72191;
       x72197 <= x72196;
       x72202 <= x72201;
       x72207 <= x72206;
       x72212 <= x72211;
       x72217 <= x72216;
       x72222 <= x72221;
       x72227 <= x72226;
       x72232 <= x72231;
       x72237 <= x72236;
       x72242 <= x72241;
       x72247 <= x72246;
       x72252 <= x72251;
       x72257 <= x72256;
       x72262 <= x72261;
       x72267 <= x72266;
       x72272 <= x72271;
       x72277 <= x72276;
       x72282 <= x72281;
       x72287 <= x72286;
       x72292 <= x72291;
       x72297 <= x72296;
       x72302 <= x72301;
       x72307 <= x72306;
       x72312 <= x72311;
       x72317 <= x72316;
       x72322 <= x72321;
       x72327 <= x72326;
       x72332 <= x72331;
       x72337 <= x72336;
       x72342 <= x72341;
       x72347 <= x72346;
       x72352 <= x72351;
       x72357 <= x72356;
       x72362 <= x72361;
       x72367 <= x72366;
       x72372 <= x72371;
       x72377 <= x72376;
       x72382 <= x72381;
       x72387 <= x72386;
       x72392 <= x72391;
       x72397 <= x72396;
       x72402 <= x72401;
       x72407 <= x72406;
       x72412 <= x72411;
       x72417 <= x72416;
       x72422 <= x72421;
       x72427 <= x72426;
       x72432 <= x72431;
       x72437 <= x72436;
       x72442 <= x72441;
       x72447 <= x72446;
       x72452 <= x72451;
       x72457 <= x72456;
       x72462 <= x72461;
       x72467 <= x72466;
       x72472 <= x72471;
       x72477 <= x72476;
       x72482 <= x72481;
       x72487 <= x72486;
       x72492 <= x72491;
       x72497 <= x72496;
       x72502 <= x72501;
       x72507 <= x72506;
       x72512 <= x72511;
       x72517 <= x72516;
       x72522 <= x72521;
       x72527 <= x72526;
       x72532 <= x72531;
       x72537 <= x72536;
       x72542 <= x72541;
       x72547 <= x72546;
       x72552 <= x72551;
       x72557 <= x72556;
       x72562 <= x72561;
       x72567 <= x72566;
       x72572 <= x72571;
       x72577 <= x72576;
       x72582 <= x72581;
       x72587 <= x72586;
       x72592 <= x72591;
       x72597 <= x72596;
       x72602 <= x72601;
       x72607 <= x72606;
       x72612 <= x72611;
       x72617 <= x72616;
       x72622 <= x72621;
       x72627 <= x72626;
       x72632 <= x72631;
       x72637 <= x72636;
       x72642 <= x72641;
       x72647 <= x72646;
       x72652 <= x72651;
       x72657 <= x72656;
       x72662 <= x72661;
       x72667 <= x72666;
       x72672 <= x72671;
       x72677 <= x72676;
       x72682 <= x72681;
       x72687 <= x72686;
       x72692 <= x72691;
       x72697 <= x72696;
       x72702 <= x72701;
       x72707 <= x72706;
       x72712 <= x72711;
       x72717 <= x72716;
       x72722 <= x72721;
       x72727 <= x72726;
       x72732 <= x72731;
       x72737 <= x72736;
       x72742 <= x72741;
       x72747 <= x72746;
       x72752 <= x72751;
       x72757 <= x72756;
       x72762 <= x72761;
       x72767 <= x72766;
       x72772 <= x72771;
       x72777 <= x72776;
       x72782 <= x72781;
       x72787 <= x72786;
       x72792 <= x72791;
       x72797 <= x72796;
       x72802 <= x72801;
       x72807 <= x72806;
       x72812 <= x72811;
       x72817 <= x72816;
       x72822 <= x72821;
       x72827 <= x72826;
       x72832 <= x72831;
       x72837 <= x72836;
       x72842 <= x72841;
       x72847 <= x72846;
       x72852 <= x72851;
       x72857 <= x72856;
       x72862 <= x72861;
       x72867 <= x72866;
       x72872 <= x72871;
       x72877 <= x72876;
       x72882 <= x72881;
       x72887 <= x72886;
       x72892 <= x72891;
       x72897 <= x72896;
       x72902 <= x72901;
       x72907 <= x72906;
       x72912 <= x72911;
       x72917 <= x72916;
       x72922 <= x72921;
       x72927 <= x72926;
       x72932 <= x72931;
       x72937 <= x72936;
       x72942 <= x72941;
       x72947 <= x72946;
       x72952 <= x72951;
       x72957 <= x72956;
       x72962 <= x72961;
       x72967 <= x72966;
       x72972 <= x72971;
       x72977 <= x72976;
       x72982 <= x72981;
       x72987 <= x72986;
       x72992 <= x72991;
       x72997 <= x72996;
       x73002 <= x73001;
       x73007 <= x73006;
       x73012 <= x73011;
       x73017 <= x73016;
       x73022 <= x73021;
       x73027 <= x73026;
       x73032 <= x73031;
       x73037 <= x73036;
       x73042 <= x73041;
       x73047 <= x73046;
       x73052 <= x73051;
       x73057 <= x73056;
       x73062 <= x73061;
       x73067 <= x73066;
       x73072 <= x73071;
       x73077 <= x73076;
       x73082 <= x73081;
       x73087 <= x73086;
       x73092 <= x73091;
       x73097 <= x73096;
       x73102 <= x73101;
       x73107 <= x73106;
       x73112 <= x73111;
       x73117 <= x73116;
       x73122 <= x73121;
       x73127 <= x73126;
       x73132 <= x73131;
       x73137 <= x73136;
       x73142 <= x73141;
       x73147 <= x73146;
       x73152 <= x73151;
       x73157 <= x73156;
       x73162 <= x73161;
       x73167 <= x73166;
       x73172 <= x73171;
       x73177 <= x73176;
       x73182 <= x73181;
       x73187 <= x73186;
       x73192 <= x73191;
       x73197 <= x73196;
       x73202 <= x73201;
       x73207 <= x73206;
       x73212 <= x73211;
       x73217 <= x73216;
       x73222 <= x73221;
       x73227 <= x73226;
       x73232 <= x73231;
       x73237 <= x73236;
       x73242 <= x73241;
       x73247 <= x73246;
       x73252 <= x73251;
       x73257 <= x73256;
       x73262 <= x73261;
       x73267 <= x73266;
       x73272 <= x73271;
       x73277 <= x73276;
       x73282 <= x73281;
       x73287 <= x73286;
       x73292 <= x73291;
       x73297 <= x73296;
       x73302 <= x73301;
       x73307 <= x73306;
       x73312 <= x73311;
       x73317 <= x73316;
       x73322 <= x73321;
       x73327 <= x73326;
       x73332 <= x73331;
       x73337 <= x73336;
       x73342 <= x73341;
       x73347 <= x73346;
       x73352 <= x73351;
       x73357 <= x73356;
       x73362 <= x73361;
       x73367 <= x73366;
       x73372 <= x73371;
       x73377 <= x73376;
       x73382 <= x73381;
       x73387 <= x73386;
       x73392 <= x73391;
       x73397 <= x73396;
       x73402 <= x73401;
       x73407 <= x73406;
       x73412 <= x73411;
       x73417 <= x73416;
       x73422 <= x73421;
       x73427 <= x73426;
       x73432 <= x73431;
       x73437 <= x73436;
       x73442 <= x73441;
       x73447 <= x73446;
       x73452 <= x73451;
       x73457 <= x73456;
       x73462 <= x73461;
       x73467 <= x73466;
       x73472 <= x73471;
       x73477 <= x73476;
       x73482 <= x73481;
       x73487 <= x73486;
       x73492 <= x73491;
       x73497 <= x73496;
       x73502 <= x73501;
       x73507 <= x73506;
       x73512 <= x73511;
       x73517 <= x73516;
       x73522 <= x73521;
       x73527 <= x73526;
       x73532 <= x73531;
       x73537 <= x73536;
       x73542 <= x73541;
       x73547 <= x73546;
       x73552 <= x73551;
       x73557 <= x73556;
       x73562 <= x73561;
       x73567 <= x73566;
       x73572 <= x73571;
       x73577 <= x73576;
       x73582 <= x73581;
       x73587 <= x73586;
       x73592 <= x73591;
       x73597 <= x73596;
       x73602 <= x73601;
       x73607 <= x73606;
       x73612 <= x73611;
       x73617 <= x73616;
       x73622 <= x73621;
       x73627 <= x73626;
       x73632 <= x73631;
       x73637 <= x73636;
       x73642 <= x73641;
       x73647 <= x73646;
       x73652 <= x73651;
       x73657 <= x73656;
       x73662 <= x73661;
       x73667 <= x73666;
       x73672 <= x73671;
       x73677 <= x73676;
       x73682 <= x73681;
       x73687 <= x73686;
       x73692 <= x73691;
       x73697 <= x73696;
       x73702 <= x73701;
       x73707 <= x73706;
       x73712 <= x73711;
       x73717 <= x73716;
       x73722 <= x73721;
       x73727 <= x73726;
       x73732 <= x73731;
       x73737 <= x73736;
       x73742 <= x73741;
       x73747 <= x73746;
       x73752 <= x73751;
       x73757 <= x73756;
       x73762 <= x73761;
       x73767 <= x73766;
       x73772 <= x73771;
       x73777 <= x73776;
       x73782 <= x73781;
       x73787 <= x73786;
       x73792 <= x73791;
       x73797 <= x73796;
       x73802 <= x73801;
       x73807 <= x73806;
       x73812 <= x73811;
       x73817 <= x73816;
       x73822 <= x73821;
       x73827 <= x73826;
       x73832 <= x73831;
       x73837 <= x73836;
       x73842 <= x73841;
       x73847 <= x73846;
       x73852 <= x73851;
       x73857 <= x73856;
       x73862 <= x73861;
       x73867 <= x73866;
       x73872 <= x73871;
       x73877 <= x73876;
       x73882 <= x73881;
       x73887 <= x73886;
       x73892 <= x73891;
       x73897 <= x73896;
       x73902 <= x73901;
       x73907 <= x73906;
       x73912 <= x73911;
       x73917 <= x73916;
       x73922 <= x73921;
       x73927 <= x73926;
       x73932 <= x73931;
       x73937 <= x73936;
       x73942 <= x73941;
       x73947 <= x73946;
       x73952 <= x73951;
       x73957 <= x73956;
       x73962 <= x73961;
       x73967 <= x73966;
       x73972 <= x73971;
       x73977 <= x73976;
       x73982 <= x73981;
       x73987 <= x73986;
       x73992 <= x73991;
       x73997 <= x73996;
       x74002 <= x74001;
       x74005 <= x74004;
       x74008 <= x74007;
       x74011 <= x74010;
       x74014 <= x74013;
       x74017 <= x74016;
       x74020 <= x74019;
       x74023 <= x74022;
       x74026 <= x74025;
       x74029 <= x74028;
       x74032 <= x74031;
       x74035 <= x74034;
       x74038 <= x74037;
       x74041 <= x74040;
       x74044 <= x74043;
       x74047 <= x74046;
       x74050 <= x74049;
       x74053 <= x74052;
       x74056 <= x74055;
       x74059 <= x74058;
       x74062 <= x74061;
       x74065 <= x74064;
       x74068 <= x74067;
       x74071 <= x74070;
       x74074 <= x74073;
       x74077 <= x74076;
       x74080 <= x74079;
       x74083 <= x74082;
       x74086 <= x74085;
       x74089 <= x74088;
       x74092 <= x74091;
       x74095 <= x74094;
       x74098 <= x74097;
       x74101 <= x74100;
       x74104 <= x74103;
       x74107 <= x74106;
       x74110 <= x74109;
       x74113 <= x74112;
       x74116 <= x74115;
       x74119 <= x74118;
       x74122 <= x74121;
       x74125 <= x74124;
       x74128 <= x74127;
       x74131 <= x74130;
       x74134 <= x74133;
       x74137 <= x74136;
       x74140 <= x74139;
       x74143 <= x74142;
       x74146 <= x74145;
       x74149 <= x74148;
       x74152 <= x74151;
       x74155 <= x74154;
       x74158 <= x74157;
       x74161 <= x74160;
       x74164 <= x74163;
       x74167 <= x74166;
       x74170 <= x74169;
       x74173 <= x74172;
       x74176 <= x74175;
       x74179 <= x74178;
       x74182 <= x74181;
       x74185 <= x74184;
       x74188 <= x74187;
       x74191 <= x74190;
       x74194 <= x74193;
       x74197 <= x74196;
       x74200 <= x74199;
       x74203 <= x74202;
       x74206 <= x74205;
       x74209 <= x74208;
       x74212 <= x74211;
       x74215 <= x74214;
       x74218 <= x74217;
       x74221 <= x74220;
       x74224 <= x74223;
       x74227 <= x74226;
       x74230 <= x74229;
       x74233 <= x74232;
       x74236 <= x74235;
       x74239 <= x74238;
       x74242 <= x74241;
       x74245 <= x74244;
       x74248 <= x74247;
       x74251 <= x74250;
       x74254 <= x74253;
       x74257 <= x74256;
       x74260 <= x74259;
       x74263 <= x74262;
       x74266 <= x74265;
       x74269 <= x74268;
       x74272 <= x74271;
       x74275 <= x74274;
       x74278 <= x74277;
       x74281 <= x74280;
       x74284 <= x74283;
       x74287 <= x74286;
       x74290 <= x74289;
       x74293 <= x74292;
       x74296 <= x74295;
       x74299 <= x74298;
       x74302 <= x74301;
       x74305 <= x74304;
       x74308 <= x74307;
       x74311 <= x74310;
       x74314 <= x74313;
       x74317 <= x74316;
       x74320 <= x74319;
       x74323 <= x74322;
       x74326 <= x74325;
       x74329 <= x74328;
       x74332 <= x74331;
       x74335 <= x74334;
       x74338 <= x74337;
       x74341 <= x74340;
       x74344 <= x74343;
       x74347 <= x74346;
       x74350 <= x74349;
       x74353 <= x74352;
       x74356 <= x74355;
       x74359 <= x74358;
       x74362 <= x74361;
       x74365 <= x74364;
       x74368 <= x74367;
       x74371 <= x74370;
       x74374 <= x74373;
       x74377 <= x74376;
       x74380 <= x74379;
       x74383 <= x74382;
       x74386 <= x74385;
       x74389 <= x74388;
       x74392 <= x74391;
       x74395 <= x74394;
       x74398 <= x74397;
       x74401 <= x74400;
       x74404 <= x74403;
       x74407 <= x74406;
       x74410 <= x74409;
       x74413 <= x74412;
       x74416 <= x74415;
       x74419 <= x74418;
       x74422 <= x74421;
       x74425 <= x74424;
       x74428 <= x74427;
       x74431 <= x74430;
       x74434 <= x74433;
       x74437 <= x74436;
       x74440 <= x74439;
       x74443 <= x74442;
       x74446 <= x74445;
       x74449 <= x74448;
       x74452 <= x74451;
       x74455 <= x74454;
       x74458 <= x74457;
       x74461 <= x74460;
       x74464 <= x74463;
       x74467 <= x74466;
       x74470 <= x74469;
       x74473 <= x74472;
       x74476 <= x74475;
       x74479 <= x74478;
       x74482 <= x74481;
       x74485 <= x74484;
       x74488 <= x74487;
       x74491 <= x74490;
       x74494 <= x74493;
       x74497 <= x74496;
       x74500 <= x74499;
       x74503 <= x74502;
       x74506 <= x74505;
       x74509 <= x74508;
       x74512 <= x74511;
       x74515 <= x74514;
       x74518 <= x74517;
       x74521 <= x74520;
       x74524 <= x74523;
       x74527 <= x74526;
       x74530 <= x74529;
       x74533 <= x74532;
       x74536 <= x74535;
       x74539 <= x74538;
       x74542 <= x74541;
       x74545 <= x74544;
       x74548 <= x74547;
       x74551 <= x74550;
       x74554 <= x74553;
       x74557 <= x74556;
       x74560 <= x74559;
       x74563 <= x74562;
       x74566 <= x74565;
       x74569 <= x74568;
       x74572 <= x74571;
       x74575 <= x74574;
       x74578 <= x74577;
       x74581 <= x74580;
       x74584 <= x74583;
       x74587 <= x74586;
       x74590 <= x74589;
       x74593 <= x74592;
       x74596 <= x74595;
       x74599 <= x74598;
       x74602 <= x74601;
       x74605 <= x74604;
       x74608 <= x74607;
       x74611 <= x74610;
       x74614 <= x74613;
       x74617 <= x74616;
       x74620 <= x74619;
       x74623 <= x74622;
       x74626 <= x74625;
       x74629 <= x74628;
       x74632 <= x74631;
       x74635 <= x74634;
       x74638 <= x74637;
       x74641 <= x74640;
       x74644 <= x74643;
       x74647 <= x74646;
       x74650 <= x74649;
       x74653 <= x74652;
       x74656 <= x74655;
       x74659 <= x74658;
       x74662 <= x74661;
       x74665 <= x74664;
       x74668 <= x74667;
       x74671 <= x74670;
       x74674 <= x74673;
       x74677 <= x74676;
       x74680 <= x74679;
       x74683 <= x74682;
       x74686 <= x74685;
       x74689 <= x74688;
       x74692 <= x74691;
       x74695 <= x74694;
       x74698 <= x74697;
       x74701 <= x74700;
       x74704 <= x74703;
       x74707 <= x74706;
       x74710 <= x74709;
       x74713 <= x74712;
       x74716 <= x74715;
       x74719 <= x74718;
       x74722 <= x74721;
       x74725 <= x74724;
       x74728 <= x74727;
       x74731 <= x74730;
       x74734 <= x74733;
       x74737 <= x74736;
       x74740 <= x74739;
       x74743 <= x74742;
       x74746 <= x74745;
       x74749 <= x74748;
       x74752 <= x74751;
       x74755 <= x74754;
       x74758 <= x74757;
       x74761 <= x74760;
       x74764 <= x74763;
       x74767 <= x74766;
       x74770 <= x74769;
       x74773 <= x74772;
       x74776 <= x74775;
       x74779 <= x74778;
       x74782 <= x74781;
       x74785 <= x74784;
       x74788 <= x74787;
       x74791 <= x74790;
       x74794 <= x74793;
       x74797 <= x74796;
       x74800 <= x74799;
       x74803 <= x74802;
       x74806 <= x74805;
       x74809 <= x74808;
       x74812 <= x74811;
       x74815 <= x74814;
       x74818 <= x74817;
       x74821 <= x74820;
       x74824 <= x74823;
       x74827 <= x74826;
       x74830 <= x74829;
       x74833 <= x74832;
       x74836 <= x74835;
       x74839 <= x74838;
       x74842 <= x74841;
       x74845 <= x74844;
       x74848 <= x74847;
       x74851 <= x74850;
       x74854 <= x74853;
       x74857 <= x74856;
       x74860 <= x74859;
       x74863 <= x74862;
       x74866 <= x74865;
       x74869 <= x74868;
       x74872 <= x74871;
       x74875 <= x74874;
       x74878 <= x74877;
       x74881 <= x74880;
       x74884 <= x74883;
       x74887 <= x74886;
       x74890 <= x74889;
       x74893 <= x74892;
       x74896 <= x74895;
       x74899 <= x74898;
       x74902 <= x74901;
       x74905 <= x74904;
       x74908 <= x74907;
       x74911 <= x74910;
       x74914 <= x74913;
       x74917 <= x74916;
       x74920 <= x74919;
       x74923 <= x74922;
       x74926 <= x74925;
       x74929 <= x74928;
       x74932 <= x74931;
       x74935 <= x74934;
       x74938 <= x74937;
       x74941 <= x74940;
       x74944 <= x74943;
       x74947 <= x74946;
       x74950 <= x74949;
       x74953 <= x74952;
       x74956 <= x74955;
       x74959 <= x74958;
       x74962 <= x74961;
       x74965 <= x74964;
       x74968 <= x74967;
       x74971 <= x74970;
       x74974 <= x74973;
       x74977 <= x74976;
       x74980 <= x74979;
       x74983 <= x74982;
       x74986 <= x74985;
       x74989 <= x74988;
       x74992 <= x74991;
       x74995 <= x74994;
       x74998 <= x74997;
       x75001 <= x75000;
       x75004 <= x75003;
       x75007 <= x75006;
       x75010 <= x75009;
       x75013 <= x75012;
       x75016 <= x75015;
       x75019 <= x75018;
       x75022 <= x75021;
       x75025 <= x75024;
       x75028 <= x75027;
       x75031 <= x75030;
       x75034 <= x75033;
       x75037 <= x75036;
       x75040 <= x75039;
       x75043 <= x75042;
       x75046 <= x75045;
       x75049 <= x75048;
       x75052 <= x75051;
       x75055 <= x75054;
       x75058 <= x75057;
       x75061 <= x75060;
       x75064 <= x75063;
       x75067 <= x75066;
       x75070 <= x75069;
       x75073 <= x75072;
       x75076 <= x75075;
       x75079 <= x75078;
       x75082 <= x75081;
       x75085 <= x75084;
       x75088 <= x75087;
       x75091 <= x75090;
       x75094 <= x75093;
       x75097 <= x75096;
       x75100 <= x75099;
       x75103 <= x75102;
       x75106 <= x75105;
       x75109 <= x75108;
       x75112 <= x75111;
       x75115 <= x75114;
       x75118 <= x75117;
       x75121 <= x75120;
       x75124 <= x75123;
       x75127 <= x75126;
       x75130 <= x75129;
       x75133 <= x75132;
       x75136 <= x75135;
       x75139 <= x75138;
       x75142 <= x75141;
       x75145 <= x75144;
       x75148 <= x75147;
       x75151 <= x75150;
       x75154 <= x75153;
       x75157 <= x75156;
       x75160 <= x75159;
       x75163 <= x75162;
       x75166 <= x75165;
       x75169 <= x75168;
       x75172 <= x75171;
       x75175 <= x75174;
       x75178 <= x75177;
       x75181 <= x75180;
       x75184 <= x75183;
       x75187 <= x75186;
       x75190 <= x75189;
       x75193 <= x75192;
       x75196 <= x75195;
       x75199 <= x75198;
       x75202 <= x75201;
       x75205 <= x75204;
       x75208 <= x75207;
       x75211 <= x75210;
       x75214 <= x75213;
       x75217 <= x75216;
       x75220 <= x75219;
       x75223 <= x75222;
       x75226 <= x75225;
       x75229 <= x75228;
       x75232 <= x75231;
       x75235 <= x75234;
       x75238 <= x75237;
       x75241 <= x75240;
       x75244 <= x75243;
       x75247 <= x75246;
       x75250 <= x75249;
       x75253 <= x75252;
       x75256 <= x75255;
       x75259 <= x75258;
       x75262 <= x75261;
       x75265 <= x75264;
       x75268 <= x75267;
       x75271 <= x75270;
       x75274 <= x75273;
       x75277 <= x75276;
       x75280 <= x75279;
       x75283 <= x75282;
       x75286 <= x75285;
       x75289 <= x75288;
       x75292 <= x75291;
       x75295 <= x75294;
       x75298 <= x75297;
       x75301 <= x75300;
       x75304 <= x75303;
       x75307 <= x75306;
       x75310 <= x75309;
       x75313 <= x75312;
       x75316 <= x75315;
       x75319 <= x75318;
       x75322 <= x75321;
       x75325 <= x75324;
       x75328 <= x75327;
       x75331 <= x75330;
       x75334 <= x75333;
       x75337 <= x75336;
       x75340 <= x75339;
       x75343 <= x75342;
       x75346 <= x75345;
       x75349 <= x75348;
       x75352 <= x75351;
       x75355 <= x75354;
       x75358 <= x75357;
       x75361 <= x75360;
       x75364 <= x75363;
       x75367 <= x75366;
       x75370 <= x75369;
       x75373 <= x75372;
       x75376 <= x75375;
       x75379 <= x75378;
       x75382 <= x75381;
       x75385 <= x75384;
       x75388 <= x75387;
       x75391 <= x75390;
       x75394 <= x75393;
       x75397 <= x75396;
       x75400 <= x75399;
       x75403 <= x75402;
       x75406 <= x75405;
       x75409 <= x75408;
       x75412 <= x75411;
       x75415 <= x75414;
       x75418 <= x75417;
       x75421 <= x75420;
       x75424 <= x75423;
       x75427 <= x75426;
       x75430 <= x75429;
       x75433 <= x75432;
       x75436 <= x75435;
       x75439 <= x75438;
       x75442 <= x75441;
       x75445 <= x75444;
       x75448 <= x75447;
       x75451 <= x75450;
       x75454 <= x75453;
       x75457 <= x75456;
       x75460 <= x75459;
       x75463 <= x75462;
       x75466 <= x75465;
       x75469 <= x75468;
       x75472 <= x75471;
       x75475 <= x75474;
       x75478 <= x75477;
       x75481 <= x75480;
       x75484 <= x75483;
       x75487 <= x75486;
       x75490 <= x75489;
       x75493 <= x75492;
       x75496 <= x75495;
       x75499 <= x75498;
       x75502 <= x75501;
       x75505 <= x75504;
       x75508 <= x75507;
       x75511 <= x75510;
       x75514 <= x75513;
       x75517 <= x75516;
       x75520 <= x75519;
       x75523 <= x75522;
       x75526 <= x75525;
       x75529 <= x75528;
       x75532 <= x75531;
       x75535 <= x75534;
       x75538 <= x75537;
       x75541 <= x75540;
       x75544 <= x75543;
       x75547 <= x75546;
       x75550 <= x75549;
       x75553 <= x75552;
       x75556 <= x75555;
       x75559 <= x75558;
       x75562 <= x75561;
       x75565 <= x75564;
       x75568 <= x75567;
       x75571 <= x75570;
       x75574 <= x75573;
       x75577 <= x75576;
       x75580 <= x75579;
       x75583 <= x75582;
       x75586 <= x75585;
       x75589 <= x75588;
       x75592 <= x75591;
       x75595 <= x75594;
       x75598 <= x75597;
       x75601 <= x75600;
       x75604 <= x75603;
       x75607 <= x75606;
       x75610 <= x75609;
       x75613 <= x75612;
       x75616 <= x75615;
       x75619 <= x75618;
       x75622 <= x75621;
       x75625 <= x75624;
       x75628 <= x75627;
       x75631 <= x75630;
       x75634 <= x75633;
       x75637 <= x75636;
       x75640 <= x75639;
       x75643 <= x75642;
       x75646 <= x75645;
       x75649 <= x75648;
       x75652 <= x75651;
       x75655 <= x75654;
       x75658 <= x75657;
       x75661 <= x75660;
       x75664 <= x75663;
       x75667 <= x75666;
       x75670 <= x75669;
       x75673 <= x75672;
       x75676 <= x75675;
       x75679 <= x75678;
       x75682 <= x75681;
       x75685 <= x75684;
       x75688 <= x75687;
       x75691 <= x75690;
       x75694 <= x75693;
       x75697 <= x75696;
       x75700 <= x75699;
       x75703 <= x75702;
       x75706 <= x75705;
       x75709 <= x75708;
       x75712 <= x75711;
       x75715 <= x75714;
       x75718 <= x75717;
       x75721 <= x75720;
       x75724 <= x75723;
       x75727 <= x75726;
       x75730 <= x75729;
       x75733 <= x75732;
       x75736 <= x75735;
       x75739 <= x75738;
       x75742 <= x75741;
       x75745 <= x75744;
       x75748 <= x75747;
       x75751 <= x75750;
       x75754 <= x75753;
       x75757 <= x75756;
       x75760 <= x75759;
       x75763 <= x75762;
       x75766 <= x75765;
       x75769 <= x75768;
       x75772 <= x75771;
       x75775 <= x75774;
       x75778 <= x75777;
       x75781 <= x75780;
       x75784 <= x75783;
       x75787 <= x75786;
       x75790 <= x75789;
       x75793 <= x75792;
       x75796 <= x75795;
       x75799 <= x75798;
       x75802 <= x75801;
       x75805 <= x75804;
       x75808 <= x75807;
       x75811 <= x75810;
       x75814 <= x75813;
       x75817 <= x75816;
       x75820 <= x75819;
       x75823 <= x75822;
       x75826 <= x75825;
       x75829 <= x75828;
       x75832 <= x75831;
       x75835 <= x75834;
       x75838 <= x75837;
       x75841 <= x75840;
       x75844 <= x75843;
       x75847 <= x75846;
       x75850 <= x75849;
       x75853 <= x75852;
       x75856 <= x75855;
       x75859 <= x75858;
       x75862 <= x75861;
       x75865 <= x75864;
       x75868 <= x75867;
       x75871 <= x75870;
       x75874 <= x75873;
       x75877 <= x75876;
       x75880 <= x75879;
       x75883 <= x75882;
       x75886 <= x75885;
       x75889 <= x75888;
       x75892 <= x75891;
       x75895 <= x75894;
       x75898 <= x75897;
       x75901 <= x75900;
       x75904 <= x75903;
       x75907 <= x75906;
       x75910 <= x75909;
       x75913 <= x75912;
       x75916 <= x75915;
       x75919 <= x75918;
       x75922 <= x75921;
       x75925 <= x75924;
       x75928 <= x75927;
       x75931 <= x75930;
       x75934 <= x75933;
       x75937 <= x75936;
       x75940 <= x75939;
       x75943 <= x75942;
       x75946 <= x75945;
       x75949 <= x75948;
       x75952 <= x75951;
       x75955 <= x75954;
       x75958 <= x75957;
       x75961 <= x75960;
       x75964 <= x75963;
       x75967 <= x75966;
       x75970 <= x75969;
       x75973 <= x75972;
       x75976 <= x75975;
       x75979 <= x75978;
       x75982 <= x75981;
       x75985 <= x75984;
       x75988 <= x75987;
       x75991 <= x75990;
       x75994 <= x75993;
       x75997 <= x75996;
       x76000 <= x75999;
       x76003 <= x76002;
       x76006 <= x76005;
       x76009 <= x76008;
       x76012 <= x76011;
       x76015 <= x76014;
       x76018 <= x76017;
       x76021 <= x76020;
       x76024 <= x76023;
       x76027 <= x76026;
       x76030 <= x76029;
       x76033 <= x76032;
       x76036 <= x76035;
       x76039 <= x76038;
       x76042 <= x76041;
       x76045 <= x76044;
       x76048 <= x76047;
       x76051 <= x76050;
       x76054 <= x76053;
       x76057 <= x76056;
       x76060 <= x76059;
       x76063 <= x76062;
       x76066 <= x76065;
       x76069 <= x76068;
       x76072 <= x76071;
       x76075 <= x76074;
       x76078 <= x76077;
       x76081 <= x76080;
       x76084 <= x76083;
       x76087 <= x76086;
       x76090 <= x76089;
       x76093 <= x76092;
       x76096 <= x76095;
       x76099 <= x76098;
       x76102 <= x76101;
       x76105 <= x76104;
       x76108 <= x76107;
       x76111 <= x76110;
       x76114 <= x76113;
       x76117 <= x76116;
       x76120 <= x76119;
       x76123 <= x76122;
       x76126 <= x76125;
       x76129 <= x76128;
       x76132 <= x76131;
       x76135 <= x76134;
       x76138 <= x76137;
       x76141 <= x76140;
       x76144 <= x76143;
       x76147 <= x76146;
       x76150 <= x76149;
       x76153 <= x76152;
       x76156 <= x76155;
       x76159 <= x76158;
       x76162 <= x76161;
       x76165 <= x76164;
       x76168 <= x76167;
       x76171 <= x76170;
       x76174 <= x76173;
       x76177 <= x76176;
       x76180 <= x76179;
       x76183 <= x76182;
       x76186 <= x76185;
       x76189 <= x76188;
       x76192 <= x76191;
       x76195 <= x76194;
       x76198 <= x76197;
       x76201 <= x76200;
       x76204 <= x76203;
       x76207 <= x76206;
       x76210 <= x76209;
       x76213 <= x76212;
       x76216 <= x76215;
       x76219 <= x76218;
       x76222 <= x76221;
       x76225 <= x76224;
       x76228 <= x76227;
       x76231 <= x76230;
       x76234 <= x76233;
       x76237 <= x76236;
       x76240 <= x76239;
       x76243 <= x76242;
       x76246 <= x76245;
       x76249 <= x76248;
       x76252 <= x76251;
       x76255 <= x76254;
       x76258 <= x76257;
       x76261 <= x76260;
       x76264 <= x76263;
       x76267 <= x76266;
       x76270 <= x76269;
       x76273 <= x76272;
       x76276 <= x76275;
       x76279 <= x76278;
       x76282 <= x76281;
       x76285 <= x76284;
       x76288 <= x76287;
       x76291 <= x76290;
       x76294 <= x76293;
       x76297 <= x76296;
       x76300 <= x76299;
       x76303 <= x76302;
       x76306 <= x76305;
       x76309 <= x76308;
       x76312 <= x76311;
       x76315 <= x76314;
       x76318 <= x76317;
       x76321 <= x76320;
       x76324 <= x76323;
       x76327 <= x76326;
       x76330 <= x76329;
       x76333 <= x76332;
       x76336 <= x76335;
       x76339 <= x76338;
       x76342 <= x76341;
       x76345 <= x76344;
       x76348 <= x76347;
       x76351 <= x76350;
       x76354 <= x76353;
       x76357 <= x76356;
       x76360 <= x76359;
       x76363 <= x76362;
       x76366 <= x76365;
       x76369 <= x76368;
       x76372 <= x76371;
       x76375 <= x76374;
       x76378 <= x76377;
       x76381 <= x76380;
       x76384 <= x76383;
       x76387 <= x76386;
       x76390 <= x76389;
       x76393 <= x76392;
       x76396 <= x76395;
       x76399 <= x76398;
       x76402 <= x76401;
       x76405 <= x76404;
       x76408 <= x76407;
       x76411 <= x76410;
       x76414 <= x76413;
       x76417 <= x76416;
       x76420 <= x76419;
       x76423 <= x76422;
       x76426 <= x76425;
       x76429 <= x76428;
       x76432 <= x76431;
       x76435 <= x76434;
       x76438 <= x76437;
       x76441 <= x76440;
       x76444 <= x76443;
       x76447 <= x76446;
       x76450 <= x76449;
       x76453 <= x76452;
       x76456 <= x76455;
       x76459 <= x76458;
       x76462 <= x76461;
       x76465 <= x76464;
       x76468 <= x76467;
       x76471 <= x76470;
       x76474 <= x76473;
       x76477 <= x76476;
       x76480 <= x76479;
       x76483 <= x76482;
       x76486 <= x76485;
       x76489 <= x76488;
       x76492 <= x76491;
       x76495 <= x76494;
       x76498 <= x76497;
       x76501 <= x76500;
       x76504 <= x76503;
       x76507 <= x76506;
       x76510 <= x76509;
       x76513 <= x76512;
       x76516 <= x76515;
       x76519 <= x76518;
       x76522 <= x76521;
       x76525 <= x76524;
       x76528 <= x76527;
       x76531 <= x76530;
       x76534 <= x76533;
       x76537 <= x76536;
       x76540 <= x76539;
       x76543 <= x76542;
       x76546 <= x76545;
       x76549 <= x76548;
       x76552 <= x76551;
       x76555 <= x76554;
       x76558 <= x76557;
       x76561 <= x76560;
       x76564 <= x76563;
       x76567 <= x76566;
       x76570 <= x76569;
       x76573 <= x76572;
       x76576 <= x76575;
       x76579 <= x76578;
       x76582 <= x76581;
       x76585 <= x76584;
       x76588 <= x76587;
       x76591 <= x76590;
       x76594 <= x76593;
       x76597 <= x76596;
       x76600 <= x76599;
       x76603 <= x76602;
       x76606 <= x76605;
       x76609 <= x76608;
       x76612 <= x76611;
       x76615 <= x76614;
       x76618 <= x76617;
       x76621 <= x76620;
       x76624 <= x76623;
       x76627 <= x76626;
       x76630 <= x76629;
       x76633 <= x76632;
       x76636 <= x76635;
       x76639 <= x76638;
       x76642 <= x76641;
       x76645 <= x76644;
       x76648 <= x76647;
       x76651 <= x76650;
       x76654 <= x76653;
       x76657 <= x76656;
       x76660 <= x76659;
       x76663 <= x76662;
       x76666 <= x76665;
       x76669 <= x76668;
       x76672 <= x76671;
       x76675 <= x76674;
       x76678 <= x76677;
       x76681 <= x76680;
       x76684 <= x76683;
       x76687 <= x76686;
       x76690 <= x76689;
       x76693 <= x76692;
       x76696 <= x76695;
       x76699 <= x76698;
       x76702 <= x76701;
       x76705 <= x76704;
       x76708 <= x76707;
       x76711 <= x76710;
       x76714 <= x76713;
       x76717 <= x76716;
       x76720 <= x76719;
       x76723 <= x76722;
       x76726 <= x76725;
       x76729 <= x76728;
       x76732 <= x76731;
       x76735 <= x76734;
       x76738 <= x76737;
       x76741 <= x76740;
       x76744 <= x76743;
       x76747 <= x76746;
       x76750 <= x76749;
       x76753 <= x76752;
       x76756 <= x76755;
       x76759 <= x76758;
       x76762 <= x76761;
       x76765 <= x76764;
       x76768 <= x76767;
       x76771 <= x76770;
       x76774 <= x76773;
       x76777 <= x76776;
       x76780 <= x76779;
       x76783 <= x76782;
       x76786 <= x76785;
       x76789 <= x76788;
       x76792 <= x76791;
       x76795 <= x76794;
       x76798 <= x76797;
       x76801 <= x76800;
       x76804 <= x76803;
       x76807 <= x76806;
       x76810 <= x76809;
       x76813 <= x76812;
       x76816 <= x76815;
       x76819 <= x76818;
       x76822 <= x76821;
       x76825 <= x76824;
       x76828 <= x76827;
       x76831 <= x76830;
       x76834 <= x76833;
       x76837 <= x76836;
       x76840 <= x76839;
       x76843 <= x76842;
       x76846 <= x76845;
       x76849 <= x76848;
       x76852 <= x76851;
       x76855 <= x76854;
       x76858 <= x76857;
       x76861 <= x76860;
       x76864 <= x76863;
       x76867 <= x76866;
       x76870 <= x76869;
       x76873 <= x76872;
       x76876 <= x76875;
       x76879 <= x76878;
       x76882 <= x76881;
       x76885 <= x76884;
       x76888 <= x76887;
       x76891 <= x76890;
       x76894 <= x76893;
       x76897 <= x76896;
       x76900 <= x76899;
       x76903 <= x76902;
       x76906 <= x76905;
       x76909 <= x76908;
       x76912 <= x76911;
       x76915 <= x76914;
       x76918 <= x76917;
       x76921 <= x76920;
       x76924 <= x76923;
       x76927 <= x76926;
       x76930 <= x76929;
       x76933 <= x76932;
       x76936 <= x76935;
       x76939 <= x76938;
       x76942 <= x76941;
       x76945 <= x76944;
       x76948 <= x76947;
       x76951 <= x76950;
       x76954 <= x76953;
       x76957 <= x76956;
       x76960 <= x76959;
       x76963 <= x76962;
       x76966 <= x76965;
       x76969 <= x76968;
       x76972 <= x76971;
       x76975 <= x76974;
       x76978 <= x76977;
       x76981 <= x76980;
       x76984 <= x76983;
       x76987 <= x76986;
       x76990 <= x76989;
       x76993 <= x76992;
       x76996 <= x76995;
       x76999 <= x76998;
       x77002 <= x77001;
       x77005 <= x77004;
       x77008 <= x77007;
       x77011 <= x77010;
       x77014 <= x77013;
       x77017 <= x77016;
       x77020 <= x77019;
       x77023 <= x77022;
       x77026 <= x77025;
       x77029 <= x77028;
       x77032 <= x77031;
       x77035 <= x77034;
       x77038 <= x77037;
       x77041 <= x77040;
       x77044 <= x77043;
       x77047 <= x77046;
       x77050 <= x77049;
       x77053 <= x77052;
       x77056 <= x77055;
       x77059 <= x77058;
       x77062 <= x77061;
       x77065 <= x77064;
       x77068 <= x77067;
       x77071 <= x77070;
       x77074 <= x77073;
       x77077 <= x77076;
       x77080 <= x77079;
       x77083 <= x77082;
       x77086 <= x77085;
       x77089 <= x77088;
       x77092 <= x77091;
       x77095 <= x77094;
       x77098 <= x77097;
       x77101 <= x77100;
       x77104 <= x77103;
       x77107 <= x77106;
       x77110 <= x77109;
       x77113 <= x77112;
       x77116 <= x77115;
       x77119 <= x77118;
       x77122 <= x77121;
       x77125 <= x77124;
       x77128 <= x77127;
       x77131 <= x77130;
       x77134 <= x77133;
       x77137 <= x77136;
       x77140 <= x77139;
       x77143 <= x77142;
       x77146 <= x77145;
       x77149 <= x77148;
       x77152 <= x77151;
       x77155 <= x77154;
       x77158 <= x77157;
       x77161 <= x77160;
       x77164 <= x77163;
       x77167 <= x77166;
       x77170 <= x77169;
       x77173 <= x77172;
       x77176 <= x77175;
       x77179 <= x77178;
       x77182 <= x77181;
       x77185 <= x77184;
       x77188 <= x77187;
       x77191 <= x77190;
       x77194 <= x77193;
       x77197 <= x77196;
       x77200 <= x77199;
       x77203 <= x77202;
       x77206 <= x77205;
       x77209 <= x77208;
       x77212 <= x77211;
       x77215 <= x77214;
       x77218 <= x77217;
       x77221 <= x77220;
       x77224 <= x77223;
       x77227 <= x77226;
       x77230 <= x77229;
       x77233 <= x77232;
       x77236 <= x77235;
       x77239 <= x77238;
       x77242 <= x77241;
       x77245 <= x77244;
       x77248 <= x77247;
       x77251 <= x77250;
       x77254 <= x77253;
       x77257 <= x77256;
       x77260 <= x77259;
       x77263 <= x77262;
       x77266 <= x77265;
       x77269 <= x77268;
       x77272 <= x77271;
       x77275 <= x77274;
       x77278 <= x77277;
       x77281 <= x77280;
       x77284 <= x77283;
       x77287 <= x77286;
       x77290 <= x77289;
       x77293 <= x77292;
       x77296 <= x77295;
       x77299 <= x77298;
       x77302 <= x77301;
       x77305 <= x77304;
       x77308 <= x77307;
       x77311 <= x77310;
       x77314 <= x77313;
       x77317 <= x77316;
       x77320 <= x77319;
       x77323 <= x77322;
       x77326 <= x77325;
       x77329 <= x77328;
       x77332 <= x77331;
       x77335 <= x77334;
       x77338 <= x77337;
       x77341 <= x77340;
       x77344 <= x77343;
       x77347 <= x77346;
       x77350 <= x77349;
       x77353 <= x77352;
       x77356 <= x77355;
       x77359 <= x77358;
       x77362 <= x77361;
       x77365 <= x77364;
       x77368 <= x77367;
       x77371 <= x77370;
       x77374 <= x77373;
       x77377 <= x77376;
       x77380 <= x77379;
       x77383 <= x77382;
       x77386 <= x77385;
       x77389 <= x77388;
       x77392 <= x77391;
       x77395 <= x77394;
       x77398 <= x77397;
       x77401 <= x77400;
       x77404 <= x77403;
       x77407 <= x77406;
       x77410 <= x77409;
       x77413 <= x77412;
       x77416 <= x77415;
       x77419 <= x77418;
       x77422 <= x77421;
       x77425 <= x77424;
       x77428 <= x77427;
       x77431 <= x77430;
       x77434 <= x77433;
       x77437 <= x77436;
       x77440 <= x77439;
       x77443 <= x77442;
       x77446 <= x77445;
       x77449 <= x77448;
       x77452 <= x77451;
       x77455 <= x77454;
       x77458 <= x77457;
       x77461 <= x77460;
       x77464 <= x77463;
       x77467 <= x77466;
       x77470 <= x77469;
       x77473 <= x77472;
       x77476 <= x77475;
       x77479 <= x77478;
       x77482 <= x77481;
       x77485 <= x77484;
       x77488 <= x77487;
       x77491 <= x77490;
       x77494 <= x77493;
       x77497 <= x77496;
       x77500 <= x77499;
       x77503 <= x77502;
       x77506 <= x77505;
       x77509 <= x77508;
       x77512 <= x77511;
       x77515 <= x77514;
       x77518 <= x77517;
       x77521 <= x77520;
       x77524 <= x77523;
       x77527 <= x77526;
       x77530 <= x77529;
       x77533 <= x77532;
       x77536 <= x77535;
       x77539 <= x77538;
       x77542 <= x77541;
       x77545 <= x77544;
       x77548 <= x77547;
       x77551 <= x77550;
       x77554 <= x77553;
       x77557 <= x77556;
       x77560 <= x77559;
       x77563 <= x77562;
       x77566 <= x77565;
       x77569 <= x77568;
       x77572 <= x77571;
       x77575 <= x77574;
       x77578 <= x77577;
       x77581 <= x77580;
       x77584 <= x77583;
       x77587 <= x77586;
       x77590 <= x77589;
       x77593 <= x77592;
       x77596 <= x77595;
       x77599 <= x77598;
       x77602 <= x77601;
       x77605 <= x77604;
       x77608 <= x77607;
       x77611 <= x77610;
       x77614 <= x77613;
       x77617 <= x77616;
       x77620 <= x77619;
       x77623 <= x77622;
       x77626 <= x77625;
       x77629 <= x77628;
       x77632 <= x77631;
       x77635 <= x77634;
       x77638 <= x77637;
       x77641 <= x77640;
       x77644 <= x77643;
       x77647 <= x77646;
       x77650 <= x77649;
       x77653 <= x77652;
       x77656 <= x77655;
       x77659 <= x77658;
       x77662 <= x77661;
       x77665 <= x77664;
       x77668 <= x77667;
       x77671 <= x77670;
       x77674 <= x77673;
       x77677 <= x77676;
       x77680 <= x77679;
       x77683 <= x77682;
       x77686 <= x77685;
       x77689 <= x77688;
       x77692 <= x77691;
       x77695 <= x77694;
       x77698 <= x77697;
       x77701 <= x77700;
       x77704 <= x77703;
       x77707 <= x77706;
       x77710 <= x77709;
       x77713 <= x77712;
       x77716 <= x77715;
       x77719 <= x77718;
       x77722 <= x77721;
       x77725 <= x77724;
       x77728 <= x77727;
       x77731 <= x77730;
       x77734 <= x77733;
       x77737 <= x77736;
       x77740 <= x77739;
       x77743 <= x77742;
       x77746 <= x77745;
       x77749 <= x77748;
       x77752 <= x77751;
       x77755 <= x77754;
       x77758 <= x77757;
       x77761 <= x77760;
       x77764 <= x77763;
       x77767 <= x77766;
       x77770 <= x77769;
       x77773 <= x77772;
       x77776 <= x77775;
       x77779 <= x77778;
       x77782 <= x77781;
       x77785 <= x77784;
       x77788 <= x77787;
       x77791 <= x77790;
       x77794 <= x77793;
       x77797 <= x77796;
       x77800 <= x77799;
       x77803 <= x77802;
       x77806 <= x77805;
       x77809 <= x77808;
       x77812 <= x77811;
       x77815 <= x77814;
       x77818 <= x77817;
       x77821 <= x77820;
       x77824 <= x77823;
       x77827 <= x77826;
       x77830 <= x77829;
       x77833 <= x77832;
       x77836 <= x77835;
       x77839 <= x77838;
       x77842 <= x77841;
       x77845 <= x77844;
       x77848 <= x77847;
       x77851 <= x77850;
       x77854 <= x77853;
       x77857 <= x77856;
       x77860 <= x77859;
       x77863 <= x77862;
       x77866 <= x77865;
       x77869 <= x77868;
       x77872 <= x77871;
       x77875 <= x77874;
       x77878 <= x77877;
       x77881 <= x77880;
       x77884 <= x77883;
       x77887 <= x77886;
       x77890 <= x77889;
       x77893 <= x77892;
       x77896 <= x77895;
       x77899 <= x77898;
       x77902 <= x77901;
       x77905 <= x77904;
       x77908 <= x77907;
       x77911 <= x77910;
       x77914 <= x77913;
       x77917 <= x77916;
       x77920 <= x77919;
       x77923 <= x77922;
       x77926 <= x77925;
       x77929 <= x77928;
       x77932 <= x77931;
       x77935 <= x77934;
       x77938 <= x77937;
       x77941 <= x77940;
       x77944 <= x77943;
       x77947 <= x77946;
       x77950 <= x77949;
       x77953 <= x77952;
       x77956 <= x77955;
       x77959 <= x77958;
       x77962 <= x77961;
       x77965 <= x77964;
       x77968 <= x77967;
       x77971 <= x77970;
       x77974 <= x77973;
       x77977 <= x77976;
       x77980 <= x77979;
       x77983 <= x77982;
       x77986 <= x77985;
       x77989 <= x77988;
       x77992 <= x77991;
       x77995 <= x77994;
       x77998 <= x77997;
       x78001 <= x78000;
       x78004 <= x78003;
       x78007 <= x78006;
       x78010 <= x78009;
       x78013 <= x78012;
       x78016 <= x78015;
       x78019 <= x78018;
       x78022 <= x78021;
       x78025 <= x78024;
       x78028 <= x78027;
       x78031 <= x78030;
       x78034 <= x78033;
       x78037 <= x78036;
       x78040 <= x78039;
       x78043 <= x78042;
       x78046 <= x78045;
       x78049 <= x78048;
       x78052 <= x78051;
       x78055 <= x78054;
       x78058 <= x78057;
       x78061 <= x78060;
       x78064 <= x78063;
       x78067 <= x78066;
       x78070 <= x78069;
       x78073 <= x78072;
       x78076 <= x78075;
       x78079 <= x78078;
       x78082 <= x78081;
       x78085 <= x78084;
       x78088 <= x78087;
       x78091 <= x78090;
       x78094 <= x78093;
       x78097 <= x78096;
       x78100 <= x78099;
       x78103 <= x78102;
       x78106 <= x78105;
       x78109 <= x78108;
       x78112 <= x78111;
       x78115 <= x78114;
       x78118 <= x78117;
       x78121 <= x78120;
       x78124 <= x78123;
       x78127 <= x78126;
       x78130 <= x78129;
       x78133 <= x78132;
       x78136 <= x78135;
       x78139 <= x78138;
       x78142 <= x78141;
       x78145 <= x78144;
       x78148 <= x78147;
       x78151 <= x78150;
       x78154 <= x78153;
       x78157 <= x78156;
       x78160 <= x78159;
       x78163 <= x78162;
       x78166 <= x78165;
       x78169 <= x78168;
       x78172 <= x78171;
       x78175 <= x78174;
       x78178 <= x78177;
       x78181 <= x78180;
       x78184 <= x78183;
       x78187 <= x78186;
       x78190 <= x78189;
       x78193 <= x78192;
       x78196 <= x78195;
       x78199 <= x78198;
       x78202 <= x78201;
       x78205 <= x78204;
       x78208 <= x78207;
       x78211 <= x78210;
       x78214 <= x78213;
       x78217 <= x78216;
       x78220 <= x78219;
       x78223 <= x78222;
       x78226 <= x78225;
       x78229 <= x78228;
       x78232 <= x78231;
       x78235 <= x78234;
       x78238 <= x78237;
       x78241 <= x78240;
       x78244 <= x78243;
       x78247 <= x78246;
       x78250 <= x78249;
       x78253 <= x78252;
       x78256 <= x78255;
       x78259 <= x78258;
       x78262 <= x78261;
       x78265 <= x78264;
       x78268 <= x78267;
       x78271 <= x78270;
       x78274 <= x78273;
       x78277 <= x78276;
       x78280 <= x78279;
       x78283 <= x78282;
       x78286 <= x78285;
       x78289 <= x78288;
       x78292 <= x78291;
       x78295 <= x78294;
       x78298 <= x78297;
       x78301 <= x78300;
       x78304 <= x78303;
       x78307 <= x78306;
       x78310 <= x78309;
       x78313 <= x78312;
       x78316 <= x78315;
       x78319 <= x78318;
       x78322 <= x78321;
       x78325 <= x78324;
       x78328 <= x78327;
       x78331 <= x78330;
       x78334 <= x78333;
       x78337 <= x78336;
       x78340 <= x78339;
       x78343 <= x78342;
       x78346 <= x78345;
       x78349 <= x78348;
       x78352 <= x78351;
       x78355 <= x78354;
       x78358 <= x78357;
       x78361 <= x78360;
       x78364 <= x78363;
       x78367 <= x78366;
       x78370 <= x78369;
       x78373 <= x78372;
       x78376 <= x78375;
       x78379 <= x78378;
       x78382 <= x78381;
       x78385 <= x78384;
       x78388 <= x78387;
       x78391 <= x78390;
       x78394 <= x78393;
       x78397 <= x78396;
       x78400 <= x78399;
       x78403 <= x78402;
       x78406 <= x78405;
       x78409 <= x78408;
       x78412 <= x78411;
       x78415 <= x78414;
       x78418 <= x78417;
       x78421 <= x78420;
       x78424 <= x78423;
       x78427 <= x78426;
       x78430 <= x78429;
       x78433 <= x78432;
       x78436 <= x78435;
       x78439 <= x78438;
       x78442 <= x78441;
       x78445 <= x78444;
       x78448 <= x78447;
       x78451 <= x78450;
       x78454 <= x78453;
       x78457 <= x78456;
       x78460 <= x78459;
       x78463 <= x78462;
       x78466 <= x78465;
       x78469 <= x78468;
       x78472 <= x78471;
       x78475 <= x78474;
       x78478 <= x78477;
       x78481 <= x78480;
       x78484 <= x78483;
       x78487 <= x78486;
       x78490 <= x78489;
       x78493 <= x78492;
       x78496 <= x78495;
       x78499 <= x78498;
       x78502 <= x78501;
       x78505 <= x78504;
       x78508 <= x78507;
       x78511 <= x78510;
       x78514 <= x78513;
       x78517 <= x78516;
       x78520 <= x78519;
       x78523 <= x78522;
       x78526 <= x78525;
       x78529 <= x78528;
       x78532 <= x78531;
       x78535 <= x78534;
       x78538 <= x78537;
       x78541 <= x78540;
       x78544 <= x78543;
       x78547 <= x78546;
       x78550 <= x78549;
       x78553 <= x78552;
       x78556 <= x78555;
       x78559 <= x78558;
       x78562 <= x78561;
       x78565 <= x78564;
       x78568 <= x78567;
       x78571 <= x78570;
       x78574 <= x78573;
       x78577 <= x78576;
       x78580 <= x78579;
       x78583 <= x78582;
       x78586 <= x78585;
       x78589 <= x78588;
       x78592 <= x78591;
       x78595 <= x78594;
       x78598 <= x78597;
       x78601 <= x78600;
       x78604 <= x78603;
       x78607 <= x78606;
       x78610 <= x78609;
       x78613 <= x78612;
       x78616 <= x78615;
       x78619 <= x78618;
       x78622 <= x78621;
       x78625 <= x78624;
       x78628 <= x78627;
       x78631 <= x78630;
       x78634 <= x78633;
       x78637 <= x78636;
       x78640 <= x78639;
       x78643 <= x78642;
       x78646 <= x78645;
       x78649 <= x78648;
       x78652 <= x78651;
       x78655 <= x78654;
       x78658 <= x78657;
       x78661 <= x78660;
       x78664 <= x78663;
       x78667 <= x78666;
       x78670 <= x78669;
       x78673 <= x78672;
       x78676 <= x78675;
       x78679 <= x78678;
       x78682 <= x78681;
       x78685 <= x78684;
       x78688 <= x78687;
       x78691 <= x78690;
       x78694 <= x78693;
       x78697 <= x78696;
       x78700 <= x78699;
       x78703 <= x78702;
       x78706 <= x78705;
       x78709 <= x78708;
       x78712 <= x78711;
       x78715 <= x78714;
       x78718 <= x78717;
       x78721 <= x78720;
       x78724 <= x78723;
       x78727 <= x78726;
       x78730 <= x78729;
       x78733 <= x78732;
       x78736 <= x78735;
       x78739 <= x78738;
       x78742 <= x78741;
       x78745 <= x78744;
       x78748 <= x78747;
       x78751 <= x78750;
       x78754 <= x78753;
       x78757 <= x78756;
       x78760 <= x78759;
       x78763 <= x78762;
       x78766 <= x78765;
       x78769 <= x78768;
       x78772 <= x78771;
       x78775 <= x78774;
       x78778 <= x78777;
       x78781 <= x78780;
       x78784 <= x78783;
       x78787 <= x78786;
       x78790 <= x78789;
       x78793 <= x78792;
       x78796 <= x78795;
       x78799 <= x78798;
       x78802 <= x78801;
       x78805 <= x78804;
       x78808 <= x78807;
       x78811 <= x78810;
       x78814 <= x78813;
       x78817 <= x78816;
       x78820 <= x78819;
       x78823 <= x78822;
       x78826 <= x78825;
       x78829 <= x78828;
       x78832 <= x78831;
       x78835 <= x78834;
       x78838 <= x78837;
       x78841 <= x78840;
       x78844 <= x78843;
       x78847 <= x78846;
       x78850 <= x78849;
       x78853 <= x78852;
       x78856 <= x78855;
       x78859 <= x78858;
       x78862 <= x78861;
       x78865 <= x78864;
       x78868 <= x78867;
       x78871 <= x78870;
       x78874 <= x78873;
       x78877 <= x78876;
       x78880 <= x78879;
       x78883 <= x78882;
       x78886 <= x78885;
       x78889 <= x78888;
       x78892 <= x78891;
       x78895 <= x78894;
       x78898 <= x78897;
       x78901 <= x78900;
       x78904 <= x78903;
       x78907 <= x78906;
       x78910 <= x78909;
       x78913 <= x78912;
       x78916 <= x78915;
       x78919 <= x78918;
       x78922 <= x78921;
       x78925 <= x78924;
       x78928 <= x78927;
       x78931 <= x78930;
       x78934 <= x78933;
       x78937 <= x78936;
       x78940 <= x78939;
       x78943 <= x78942;
       x78946 <= x78945;
       x78949 <= x78948;
       x78952 <= x78951;
       x78955 <= x78954;
       x78958 <= x78957;
       x78961 <= x78960;
       x78964 <= x78963;
       x78967 <= x78966;
       x78970 <= x78969;
       x78973 <= x78972;
       x78976 <= x78975;
       x78979 <= x78978;
       x78982 <= x78981;
       x78985 <= x78984;
       x78988 <= x78987;
       x78991 <= x78990;
       x78994 <= x78993;
       x78997 <= x78996;
       x79000 <= x78999;
       x79003 <= x79002;
       x79006 <= x79005;
       x79009 <= x79008;
       x79012 <= x79011;
       x79015 <= x79014;
       x79018 <= x79017;
       x79021 <= x79020;
       x79024 <= x79023;
       x79027 <= x79026;
       x79030 <= x79029;
       x79033 <= x79032;
       x79036 <= x79035;
       x79039 <= x79038;
       x79042 <= x79041;
       x79045 <= x79044;
       x79048 <= x79047;
       x79051 <= x79050;
       x79054 <= x79053;
       x79057 <= x79056;
       x79060 <= x79059;
       x79063 <= x79062;
       x79066 <= x79065;
       x79069 <= x79068;
       x79072 <= x79071;
       x79075 <= x79074;
       x79078 <= x79077;
       x79081 <= x79080;
       x79084 <= x79083;
       x79087 <= x79086;
       x79090 <= x79089;
       x79093 <= x79092;
       x79096 <= x79095;
       x79099 <= x79098;
       x79102 <= x79101;
       x79105 <= x79104;
       x79108 <= x79107;
       x79111 <= x79110;
       x79114 <= x79113;
       x79117 <= x79116;
       x79120 <= x79119;
       x79123 <= x79122;
       x79126 <= x79125;
       x79129 <= x79128;
       x79132 <= x79131;
       x79135 <= x79134;
       x79138 <= x79137;
       x79141 <= x79140;
       x79144 <= x79143;
       x79147 <= x79146;
       x79150 <= x79149;
       x79153 <= x79152;
       x79156 <= x79155;
       x79159 <= x79158;
       x79162 <= x79161;
       x79165 <= x79164;
       x79168 <= x79167;
       x79171 <= x79170;
       x79174 <= x79173;
       x79177 <= x79176;
       x79180 <= x79179;
       x79183 <= x79182;
       x79186 <= x79185;
       x79189 <= x79188;
       x79192 <= x79191;
       x79195 <= x79194;
       x79198 <= x79197;
       x79201 <= x79200;
       x79204 <= x79203;
       x79207 <= x79206;
       x79210 <= x79209;
       x79213 <= x79212;
       x79216 <= x79215;
       x79219 <= x79218;
       x79222 <= x79221;
       x79225 <= x79224;
       x79228 <= x79227;
       x79231 <= x79230;
       x79234 <= x79233;
       x79237 <= x79236;
       x79240 <= x79239;
       x79243 <= x79242;
       x79246 <= x79245;
       x79249 <= x79248;
       x79252 <= x79251;
       x79255 <= x79254;
       x79258 <= x79257;
       x79261 <= x79260;
       x79264 <= x79263;
       x79267 <= x79266;
       x79270 <= x79269;
       x79273 <= x79272;
       x79276 <= x79275;
       x79279 <= x79278;
       x79282 <= x79281;
       x79285 <= x79284;
       x79288 <= x79287;
       x79291 <= x79290;
       x79294 <= x79293;
       x79297 <= x79296;
       x79300 <= x79299;
       x79303 <= x79302;
       x79306 <= x79305;
       x79309 <= x79308;
       x79312 <= x79311;
       x79315 <= x79314;
       x79318 <= x79317;
       x79321 <= x79320;
       x79324 <= x79323;
       x79327 <= x79326;
       x79330 <= x79329;
       x79333 <= x79332;
       x79336 <= x79335;
       x79339 <= x79338;
       x79342 <= x79341;
       x79345 <= x79344;
       x79348 <= x79347;
       x79351 <= x79350;
       x79354 <= x79353;
       x79357 <= x79356;
       x79360 <= x79359;
       x79363 <= x79362;
       x79366 <= x79365;
       x79369 <= x79368;
       x79372 <= x79371;
       x79375 <= x79374;
       x79378 <= x79377;
       x79381 <= x79380;
       x79384 <= x79383;
       x79387 <= x79386;
       x79390 <= x79389;
       x79393 <= x79392;
       x79396 <= x79395;
       x79399 <= x79398;
       x79402 <= x79401;
       x79405 <= x79404;
       x79408 <= x79407;
       x79411 <= x79410;
       x79414 <= x79413;
       x79417 <= x79416;
       x79420 <= x79419;
       x79423 <= x79422;
       x79426 <= x79425;
       x79429 <= x79428;
       x79432 <= x79431;
       x79435 <= x79434;
       x79438 <= x79437;
       x79441 <= x79440;
       x79444 <= x79443;
       x79447 <= x79446;
       x79450 <= x79449;
       x79453 <= x79452;
       x79456 <= x79455;
       x79459 <= x79458;
       x79462 <= x79461;
       x79465 <= x79464;
       x79468 <= x79467;
       x79471 <= x79470;
       x79474 <= x79473;
       x79477 <= x79476;
       x79480 <= x79479;
       x79483 <= x79482;
       x79486 <= x79485;
       x79489 <= x79488;
       x79492 <= x79491;
       x79495 <= x79494;
       x79498 <= x79497;
       x79501 <= x79500;
       x79504 <= x79503;
       x79507 <= x79506;
       x79510 <= x79509;
       x79513 <= x79512;
       x79516 <= x79515;
       x79519 <= x79518;
       x79522 <= x79521;
       x79525 <= x79524;
       x79528 <= x79527;
       x79531 <= x79530;
       x79534 <= x79533;
       x79537 <= x79536;
       x79540 <= x79539;
       x79543 <= x79542;
       x79546 <= x79545;
       x79549 <= x79548;
       x79552 <= x79551;
       x79555 <= x79554;
       x79558 <= x79557;
       x79561 <= x79560;
       x79564 <= x79563;
       x79567 <= x79566;
       x79570 <= x79569;
       x79573 <= x79572;
       x79576 <= x79575;
       x79579 <= x79578;
       x79582 <= x79581;
       x79585 <= x79584;
       x79588 <= x79587;
       x79591 <= x79590;
       x79594 <= x79593;
       x79597 <= x79596;
       x79600 <= x79599;
       x79603 <= x79602;
       x79606 <= x79605;
       x79609 <= x79608;
       x79612 <= x79611;
       x79615 <= x79614;
       x79618 <= x79617;
       x79621 <= x79620;
       x79624 <= x79623;
       x79627 <= x79626;
       x79630 <= x79629;
       x79633 <= x79632;
       x79636 <= x79635;
       x79639 <= x79638;
       x79642 <= x79641;
       x79645 <= x79644;
       x79648 <= x79647;
       x79651 <= x79650;
       x79654 <= x79653;
       x79657 <= x79656;
       x79660 <= x79659;
       x79663 <= x79662;
       x79666 <= x79665;
       x79669 <= x79668;
       x79672 <= x79671;
       x79675 <= x79674;
       x79678 <= x79677;
       x79681 <= x79680;
       x79684 <= x79683;
       x79687 <= x79686;
       x79690 <= x79689;
       x79693 <= x79692;
       x79696 <= x79695;
       x79699 <= x79698;
       x79702 <= x79701;
       x79705 <= x79704;
       x79708 <= x79707;
       x79711 <= x79710;
       x79714 <= x79713;
       x79717 <= x79716;
       x79720 <= x79719;
       x79723 <= x79722;
       x79726 <= x79725;
       x79729 <= x79728;
       x79732 <= x79731;
       x79735 <= x79734;
       x79738 <= x79737;
       x79741 <= x79740;
       x79744 <= x79743;
       x79747 <= x79746;
       x79750 <= x79749;
       x79753 <= x79752;
       x79756 <= x79755;
       x79759 <= x79758;
       x79762 <= x79761;
       x79765 <= x79764;
       x79768 <= x79767;
       x79771 <= x79770;
       x79774 <= x79773;
       x79777 <= x79776;
       x79780 <= x79779;
       x79783 <= x79782;
       x79786 <= x79785;
       x79789 <= x79788;
       x79792 <= x79791;
       x79795 <= x79794;
       x79798 <= x79797;
       x79801 <= x79800;
       x79804 <= x79803;
       x79807 <= x79806;
       x79810 <= x79809;
       x79813 <= x79812;
       x79816 <= x79815;
       x79819 <= x79818;
       x79822 <= x79821;
       x79825 <= x79824;
       x79828 <= x79827;
       x79831 <= x79830;
       x79834 <= x79833;
       x79837 <= x79836;
       x79840 <= x79839;
       x79843 <= x79842;
       x79846 <= x79845;
       x79849 <= x79848;
       x79852 <= x79851;
       x79855 <= x79854;
       x79858 <= x79857;
       x79861 <= x79860;
       x79864 <= x79863;
       x79867 <= x79866;
       x79870 <= x79869;
       x79873 <= x79872;
       x79876 <= x79875;
       x79879 <= x79878;
       x79882 <= x79881;
       x79885 <= x79884;
       x79888 <= x79887;
       x79891 <= x79890;
       x79894 <= x79893;
       x79897 <= x79896;
       x79900 <= x79899;
       x79903 <= x79902;
       x79906 <= x79905;
       x79909 <= x79908;
       x79912 <= x79911;
       x79915 <= x79914;
       x79918 <= x79917;
       x79921 <= x79920;
       x79924 <= x79923;
       x79927 <= x79926;
       x79930 <= x79929;
       x79933 <= x79932;
       x79936 <= x79935;
       x79939 <= x79938;
       x79942 <= x79941;
       x79945 <= x79944;
       x79948 <= x79947;
       x79951 <= x79950;
       x79954 <= x79953;
       x79957 <= x79956;
       x79960 <= x79959;
       x79963 <= x79962;
       x79966 <= x79965;
       x79969 <= x79968;
       x79972 <= x79971;
       x79975 <= x79974;
       x79978 <= x79977;
       x79981 <= x79980;
       x79984 <= x79983;
       x79987 <= x79986;
       x79990 <= x79989;
       x79993 <= x79992;
       x79996 <= x79995;
       x79999 <= x79998;
       x80002 <= x80001;
       x80005 <= x80004;
       x80008 <= x80007;
       x80011 <= x80010;
       x80014 <= x80013;
       x80017 <= x80016;
       x80020 <= x80019;
       x80023 <= x80022;
       x80026 <= x80025;
       x80029 <= x80028;
       x80032 <= x80031;
       x80035 <= x80034;
       x80038 <= x80037;
       x80041 <= x80040;
       x80044 <= x80043;
       x80047 <= x80046;
       x80050 <= x80049;
       x80053 <= x80052;
       x80056 <= x80055;
       x80059 <= x80058;
       x80062 <= x80061;
       x80065 <= x80064;
       x80068 <= x80067;
       x80071 <= x80070;
       x80074 <= x80073;
       x80077 <= x80076;
       x80080 <= x80079;
       x80083 <= x80082;
       x80086 <= x80085;
       x80089 <= x80088;
       x80092 <= x80091;
       x80095 <= x80094;
       x80098 <= x80097;
       x80101 <= x80100;
       x80104 <= x80103;
       x80107 <= x80106;
       x80110 <= x80109;
       x80113 <= x80112;
       x80116 <= x80115;
       x80119 <= x80118;
       x80122 <= x80121;
       x80125 <= x80124;
       x80128 <= x80127;
       x80131 <= x80130;
       x80134 <= x80133;
       x80137 <= x80136;
       x80140 <= x80139;
       x80143 <= x80142;
       x80146 <= x80145;
       x80149 <= x80148;
       x80152 <= x80151;
       x80155 <= x80154;
       x80158 <= x80157;
       x80161 <= x80160;
       x80164 <= x80163;
       x80167 <= x80166;
       x80170 <= x80169;
       x80173 <= x80172;
       x80176 <= x80175;
       x80179 <= x80178;
       x80182 <= x80181;
       x80185 <= x80184;
       x80188 <= x80187;
       x80191 <= x80190;
       x80194 <= x80193;
       x80197 <= x80196;
       x80200 <= x80199;
       x80203 <= x80202;
       x80206 <= x80205;
       x80209 <= x80208;
       x80212 <= x80211;
       x80215 <= x80214;
       x80218 <= x80217;
       x80221 <= x80220;
       x80224 <= x80223;
       x80227 <= x80226;
       x80230 <= x80229;
       x80233 <= x80232;
       x80236 <= x80235;
       x80239 <= x80238;
       x80242 <= x80241;
       x80245 <= x80244;
       x80248 <= x80247;
       x80251 <= x80250;
       x80254 <= x80253;
       x80257 <= x80256;
       x80260 <= x80259;
       x80263 <= x80262;
       x80266 <= x80265;
       x80269 <= x80268;
       x80272 <= x80271;
       x80275 <= x80274;
       x80278 <= x80277;
       x80281 <= x80280;
       x80284 <= x80283;
       x80287 <= x80286;
       x80290 <= x80289;
       x80293 <= x80292;
       x80296 <= x80295;
       x80299 <= x80298;
       x80302 <= x80301;
       x80305 <= x80304;
       x80308 <= x80307;
       x80311 <= x80310;
       x80314 <= x80313;
       x80317 <= x80316;
       x80320 <= x80319;
       x80323 <= x80322;
       x80326 <= x80325;
       x80329 <= x80328;
       x80332 <= x80331;
       x80335 <= x80334;
       x80338 <= x80337;
       x80341 <= x80340;
       x80344 <= x80343;
       x80347 <= x80346;
       x80350 <= x80349;
       x80353 <= x80352;
       x80356 <= x80355;
       x80359 <= x80358;
       x80362 <= x80361;
       x80365 <= x80364;
       x80368 <= x80367;
       x80371 <= x80370;
       x80374 <= x80373;
       x80377 <= x80376;
       x80380 <= x80379;
       x80383 <= x80382;
       x80386 <= x80385;
       x80389 <= x80388;
       x80392 <= x80391;
       x80395 <= x80394;
       x80398 <= x80397;
       x80401 <= x80400;
       x80404 <= x80403;
       x80407 <= x80406;
       x80410 <= x80409;
       x80413 <= x80412;
       x80416 <= x80415;
       x80419 <= x80418;
       x80422 <= x80421;
       x80425 <= x80424;
       x80428 <= x80427;
       x80431 <= x80430;
       x80434 <= x80433;
       x80437 <= x80436;
       x80440 <= x80439;
       x80443 <= x80442;
       x80446 <= x80445;
       x80449 <= x80448;
       x80452 <= x80451;
       x80455 <= x80454;
       x80458 <= x80457;
       x80461 <= x80460;
       x80464 <= x80463;
       x80467 <= x80466;
       x80470 <= x80469;
       x80473 <= x80472;
       x80476 <= x80475;
       x80479 <= x80478;
       x80482 <= x80481;
       x80485 <= x80484;
       x80488 <= x80487;
       x80491 <= x80490;
       x80494 <= x80493;
       x80497 <= x80496;
       x80500 <= x80499;
       x80503 <= x80502;
       x80506 <= x80505;
       x80509 <= x80508;
       x80512 <= x80511;
       x80515 <= x80514;
       x80518 <= x80517;
       x80521 <= x80520;
       x80524 <= x80523;
       x80527 <= x80526;
       x80530 <= x80529;
       x80533 <= x80532;
       x80536 <= x80535;
       x80539 <= x80538;
       x80542 <= x80541;
       x80545 <= x80544;
       x80548 <= x80547;
       x80551 <= x80550;
       x80554 <= x80553;
       x80557 <= x80556;
       x80560 <= x80559;
       x80563 <= x80562;
       x80566 <= x80565;
       x80569 <= x80568;
       x80572 <= x80571;
       x80575 <= x80574;
       x80578 <= x80577;
       x80581 <= x80580;
       x80584 <= x80583;
       x80587 <= x80586;
       x80590 <= x80589;
       x80593 <= x80592;
       x80596 <= x80595;
       x80599 <= x80598;
       x80602 <= x80601;
       x80605 <= x80604;
       x80608 <= x80607;
       x80611 <= x80610;
       x80614 <= x80613;
       x80617 <= x80616;
       x80620 <= x80619;
       x80623 <= x80622;
       x80626 <= x80625;
       x80629 <= x80628;
       x80632 <= x80631;
       x80635 <= x80634;
       x80638 <= x80637;
       x80641 <= x80640;
       x80644 <= x80643;
       x80647 <= x80646;
       x80650 <= x80649;
       x80653 <= x80652;
       x80656 <= x80655;
       x80659 <= x80658;
       x80662 <= x80661;
       x80665 <= x80664;
       x80668 <= x80667;
       x80671 <= x80670;
       x80674 <= x80673;
       x80677 <= x80676;
       x80680 <= x80679;
       x80683 <= x80682;
       x80686 <= x80685;
       x80689 <= x80688;
       x80692 <= x80691;
       x80695 <= x80694;
       x80698 <= x80697;
       x80701 <= x80700;
       x80704 <= x80703;
       x80707 <= x80706;
       x80710 <= x80709;
       x80713 <= x80712;
       x80716 <= x80715;
       x80719 <= x80718;
       x80722 <= x80721;
       x80725 <= x80724;
       x80728 <= x80727;
       x80731 <= x80730;
       x80734 <= x80733;
       x80737 <= x80736;
       x80740 <= x80739;
       x80743 <= x80742;
       x80746 <= x80745;
       x80749 <= x80748;
       x80752 <= x80751;
       x80755 <= x80754;
       x80758 <= x80757;
       x80761 <= x80760;
       x80764 <= x80763;
       x80767 <= x80766;
       x80770 <= x80769;
       x80773 <= x80772;
       x80776 <= x80775;
       x80779 <= x80778;
       x80782 <= x80781;
       x80785 <= x80784;
       x80788 <= x80787;
       x80791 <= x80790;
       x80794 <= x80793;
       x80797 <= x80796;
       x80800 <= x80799;
       x80803 <= x80802;
       x80806 <= x80805;
       x80809 <= x80808;
       x80812 <= x80811;
       x80815 <= x80814;
       x80818 <= x80817;
       x80821 <= x80820;
       x80824 <= x80823;
       x80827 <= x80826;
       x80830 <= x80829;
       x80833 <= x80832;
       x80836 <= x80835;
       x80839 <= x80838;
       x80842 <= x80841;
       x80845 <= x80844;
       x80848 <= x80847;
       x80851 <= x80850;
       x80854 <= x80853;
       x80857 <= x80856;
       x80860 <= x80859;
       x80863 <= x80862;
       x80866 <= x80865;
       x80869 <= x80868;
       x80872 <= x80871;
       x80875 <= x80874;
       x80878 <= x80877;
       x80881 <= x80880;
       x80884 <= x80883;
       x80887 <= x80886;
       x80890 <= x80889;
       x80893 <= x80892;
       x80896 <= x80895;
       x80899 <= x80898;
       x80902 <= x80901;
       x80905 <= x80904;
       x80908 <= x80907;
       x80911 <= x80910;
       x80914 <= x80913;
       x80917 <= x80916;
       x80920 <= x80919;
       x80923 <= x80922;
       x80926 <= x80925;
       x80929 <= x80928;
       x80932 <= x80931;
       x80935 <= x80934;
       x80938 <= x80937;
       x80941 <= x80940;
       x80944 <= x80943;
       x80947 <= x80946;
       x80950 <= x80949;
       x80953 <= x80952;
       x80956 <= x80955;
       x80959 <= x80958;
       x80962 <= x80961;
       x80965 <= x80964;
       x80968 <= x80967;
       x80971 <= x80970;
       x80974 <= x80973;
       x80977 <= x80976;
       x80980 <= x80979;
       x80983 <= x80982;
       x80986 <= x80985;
       x80989 <= x80988;
       x80992 <= x80991;
       x80995 <= x80994;
       x80998 <= x80997;
       x81001 <= x81000;
       x81004 <= x81003;
       x81007 <= x81006;
       x81010 <= x81009;
       x81013 <= x81012;
       x81016 <= x81015;
       x81019 <= x81018;
       x81022 <= x81021;
       x81025 <= x81024;
       x81028 <= x81027;
       x81031 <= x81030;
       x81034 <= x81033;
       x81037 <= x81036;
       x81040 <= x81039;
       x81043 <= x81042;
       x81046 <= x81045;
       x81049 <= x81048;
       x81052 <= x81051;
       x81055 <= x81054;
       x81058 <= x81057;
       x81061 <= x81060;
       x81064 <= x81063;
       x81067 <= x81066;
       x81070 <= x81069;
       x81073 <= x81072;
       x81076 <= x81075;
       x81079 <= x81078;
       x81082 <= x81081;
       x81085 <= x81084;
       x81088 <= x81087;
       x81091 <= x81090;
       x81094 <= x81093;
       x81097 <= x81096;
       x81100 <= x81099;
       x81103 <= x81102;
       x81106 <= x81105;
       x81109 <= x81108;
       x81112 <= x81111;
       x81115 <= x81114;
       x81118 <= x81117;
       x81121 <= x81120;
       x81124 <= x81123;
       x81127 <= x81126;
       x81130 <= x81129;
       x81133 <= x81132;
       x81136 <= x81135;
       x81139 <= x81138;
       x81142 <= x81141;
       x81145 <= x81144;
       x81148 <= x81147;
       x81151 <= x81150;
       x81154 <= x81153;
       x81157 <= x81156;
       x81160 <= x81159;
       x81163 <= x81162;
       x81166 <= x81165;
       x81169 <= x81168;
       x81172 <= x81171;
       x81175 <= x81174;
       x81178 <= x81177;
       x81181 <= x81180;
       x81184 <= x81183;
       x81187 <= x81186;
       x81190 <= x81189;
       x81193 <= x81192;
       x81196 <= x81195;
       x81199 <= x81198;
       x81202 <= x81201;
       x81205 <= x81204;
       x81208 <= x81207;
       x81211 <= x81210;
       x81214 <= x81213;
       x81217 <= x81216;
       x81220 <= x81219;
       x81223 <= x81222;
       x81226 <= x81225;
       x81229 <= x81228;
       x81232 <= x81231;
       x81235 <= x81234;
       x81238 <= x81237;
       x81241 <= x81240;
       x81244 <= x81243;
       x81247 <= x81246;
       x81250 <= x81249;
       x81253 <= x81252;
       x81256 <= x81255;
       x81259 <= x81258;
       x81262 <= x81261;
       x81265 <= x81264;
       x81268 <= x81267;
       x81271 <= x81270;
       x81274 <= x81273;
       x81277 <= x81276;
       x81280 <= x81279;
       x81283 <= x81282;
       x81286 <= x81285;
       x81289 <= x81288;
       x81292 <= x81291;
       x81295 <= x81294;
       x81298 <= x81297;
       x81301 <= x81300;
       x81304 <= x81303;
       x81307 <= x81306;
       x81310 <= x81309;
       x81313 <= x81312;
       x81316 <= x81315;
       x81319 <= x81318;
       x81322 <= x81321;
       x81325 <= x81324;
       x81328 <= x81327;
       x81331 <= x81330;
       x81334 <= x81333;
       x81337 <= x81336;
       x81340 <= x81339;
       x81343 <= x81342;
       x81346 <= x81345;
       x81349 <= x81348;
       x81352 <= x81351;
       x81355 <= x81354;
       x81358 <= x81357;
       x81361 <= x81360;
       x81364 <= x81363;
       x81367 <= x81366;
       x81370 <= x81369;
       x81373 <= x81372;
       x81376 <= x81375;
       x81379 <= x81378;
       x81382 <= x81381;
       x81385 <= x81384;
       x81388 <= x81387;
       x81391 <= x81390;
       x81394 <= x81393;
       x81397 <= x81396;
       x81400 <= x81399;
       x81403 <= x81402;
       x81406 <= x81405;
       x81409 <= x81408;
       x81412 <= x81411;
       x81415 <= x81414;
       x81418 <= x81417;
       x81421 <= x81420;
       x81424 <= x81423;
       x81427 <= x81426;
       x81430 <= x81429;
       x81433 <= x81432;
       x81436 <= x81435;
       x81439 <= x81438;
       x81442 <= x81441;
       x81445 <= x81444;
       x81448 <= x81447;
       x81451 <= x81450;
       x81454 <= x81453;
       x81457 <= x81456;
       x81460 <= x81459;
       x81463 <= x81462;
       x81466 <= x81465;
       x81469 <= x81468;
       x81472 <= x81471;
       x81475 <= x81474;
       x81478 <= x81477;
       x81481 <= x81480;
       x81484 <= x81483;
       x81487 <= x81486;
       x81490 <= x81489;
       x81493 <= x81492;
       x81496 <= x81495;
       x81499 <= x81498;
       x81502 <= x81501;
       x81505 <= x81504;
       x81508 <= x81507;
       x81511 <= x81510;
       x81514 <= x81513;
       x81517 <= x81516;
       x81520 <= x81519;
       x81523 <= x81522;
       x81526 <= x81525;
       x81529 <= x81528;
       x81532 <= x81531;
       x81535 <= x81534;
       x81538 <= x81537;
       x81541 <= x81540;
       x81544 <= x81543;
       x81547 <= x81546;
       x81550 <= x81549;
       x81553 <= x81552;
       x81556 <= x81555;
       x81559 <= x81558;
       x81562 <= x81561;
       x81565 <= x81564;
       x81568 <= x81567;
       x81571 <= x81570;
       x81574 <= x81573;
       x81577 <= x81576;
       x81580 <= x81579;
       x81583 <= x81582;
       x81586 <= x81585;
       x81589 <= x81588;
       x81592 <= x81591;
       x81595 <= x81594;
       x81598 <= x81597;
       x81601 <= x81600;
       x81604 <= x81603;
       x81607 <= x81606;
       x81610 <= x81609;
       x81613 <= x81612;
       x81616 <= x81615;
       x81619 <= x81618;
       x81622 <= x81621;
       x81625 <= x81624;
       x81628 <= x81627;
       x81631 <= x81630;
       x81634 <= x81633;
       x81637 <= x81636;
       x81640 <= x81639;
       x81643 <= x81642;
       x81646 <= x81645;
       x81649 <= x81648;
       x81652 <= x81651;
       x81655 <= x81654;
       x81658 <= x81657;
       x81661 <= x81660;
       x81664 <= x81663;
       x81667 <= x81666;
       x81670 <= x81669;
       x81673 <= x81672;
       x81676 <= x81675;
       x81679 <= x81678;
       x81682 <= x81681;
       x81685 <= x81684;
       x81688 <= x81687;
       x81691 <= x81690;
       x81694 <= x81693;
       x81697 <= x81696;
       x81700 <= x81699;
       x81703 <= x81702;
       x81706 <= x81705;
       x81709 <= x81708;
       x81712 <= x81711;
       x81715 <= x81714;
       x81718 <= x81717;
       x81721 <= x81720;
       x81724 <= x81723;
       x81727 <= x81726;
       x81730 <= x81729;
       x81733 <= x81732;
       x81736 <= x81735;
       x81739 <= x81738;
       x81742 <= x81741;
       x81745 <= x81744;
       x81748 <= x81747;
       x81751 <= x81750;
       x81754 <= x81753;
       x81757 <= x81756;
       x81760 <= x81759;
       x81763 <= x81762;
       x81766 <= x81765;
       x81769 <= x81768;
       x81772 <= x81771;
       x81775 <= x81774;
       x81778 <= x81777;
       x81781 <= x81780;
       x81784 <= x81783;
       x81787 <= x81786;
       x81790 <= x81789;
       x81793 <= x81792;
       x81796 <= x81795;
       x81799 <= x81798;
       x81802 <= x81801;
       x81805 <= x81804;
       x81808 <= x81807;
       x81811 <= x81810;
       x81814 <= x81813;
       x81817 <= x81816;
       x81820 <= x81819;
       x81823 <= x81822;
       x81826 <= x81825;
       x81829 <= x81828;
       x81832 <= x81831;
       x81835 <= x81834;
       x81838 <= x81837;
       x81841 <= x81840;
       x81844 <= x81843;
       x81847 <= x81846;
       x81850 <= x81849;
       x81853 <= x81852;
       x81856 <= x81855;
       x81859 <= x81858;
       x81862 <= x81861;
       x81865 <= x81864;
       x81868 <= x81867;
       x81871 <= x81870;
       x81874 <= x81873;
       x81877 <= x81876;
       x81880 <= x81879;
       x81883 <= x81882;
       x81886 <= x81885;
       x81889 <= x81888;
       x81892 <= x81891;
       x81895 <= x81894;
       x81898 <= x81897;
       x81901 <= x81900;
       x81904 <= x81903;
       x81907 <= x81906;
       x81910 <= x81909;
       x81913 <= x81912;
       x81916 <= x81915;
       x81919 <= x81918;
       x81922 <= x81921;
       x81925 <= x81924;
       x81928 <= x81927;
       x81931 <= x81930;
       x81934 <= x81933;
       x81937 <= x81936;
       x81940 <= x81939;
       x81943 <= x81942;
       x81946 <= x81945;
       x81949 <= x81948;
       x81952 <= x81951;
       x81955 <= x81954;
       x81958 <= x81957;
       x81961 <= x81960;
       x81964 <= x81963;
       x81967 <= x81966;
       x81970 <= x81969;
       x81973 <= x81972;
       x81976 <= x81975;
       x81979 <= x81978;
       x81982 <= x81981;
       x81985 <= x81984;
       x81988 <= x81987;
       x81991 <= x81990;
       x81994 <= x81993;
       x81997 <= x81996;
       x82000 <= x81999;
       x82003 <= x82002;
       x82006 <= x82005;
       x82009 <= x82008;
       x82012 <= x82011;
       x82015 <= x82014;
       x82018 <= x82017;
       x82021 <= x82020;
       x82024 <= x82023;
       x82027 <= x82026;
       x82030 <= x82029;
       x82033 <= x82032;
       x82036 <= x82035;
       x82039 <= x82038;
       x82042 <= x82041;
       x82045 <= x82044;
       x82048 <= x82047;
       x82051 <= x82050;
       x82054 <= x82053;
       x82057 <= x82056;
       x82060 <= x82059;
       x82063 <= x82062;
       x82066 <= x82065;
       x82069 <= x82068;
       x82072 <= x82071;
       x82075 <= x82074;
       x82078 <= x82077;
       x82081 <= x82080;
       x82084 <= x82083;
       x82087 <= x82086;
       x82090 <= x82089;
       x82093 <= x82092;
       x82096 <= x82095;
       x82099 <= x82098;
       x82102 <= x82101;
       x82105 <= x82104;
       x82108 <= x82107;
       x82111 <= x82110;
       x82114 <= x82113;
       x82117 <= x82116;
       x82120 <= x82119;
       x82123 <= x82122;
       x82126 <= x82125;
       x82129 <= x82128;
       x82132 <= x82131;
       x82135 <= x82134;
       x82138 <= x82137;
       x82141 <= x82140;
       x82144 <= x82143;
       x82147 <= x82146;
       x82150 <= x82149;
       x82153 <= x82152;
       x82156 <= x82155;
       x82159 <= x82158;
       x82162 <= x82161;
       x82165 <= x82164;
       x82168 <= x82167;
       x82171 <= x82170;
       x82174 <= x82173;
       x82177 <= x82176;
       x82180 <= x82179;
       x82183 <= x82182;
       x82186 <= x82185;
       x82189 <= x82188;
       x82192 <= x82191;
       x82195 <= x82194;
       x82198 <= x82197;
       x82201 <= x82200;
       x82204 <= x82203;
       x82207 <= x82206;
       x82210 <= x82209;
       x82213 <= x82212;
       x82216 <= x82215;
       x82219 <= x82218;
       x82222 <= x82221;
       x82225 <= x82224;
       x82228 <= x82227;
       x82231 <= x82230;
       x82234 <= x82233;
       x82237 <= x82236;
       x82240 <= x82239;
       x82243 <= x82242;
       x82246 <= x82245;
       x82249 <= x82248;
       x82252 <= x82251;
       x82255 <= x82254;
       x82258 <= x82257;
       x82261 <= x82260;
       x82264 <= x82263;
       x82267 <= x82266;
       x82270 <= x82269;
       x82273 <= x82272;
       x82276 <= x82275;
       x82279 <= x82278;
       x82282 <= x82281;
       x82285 <= x82284;
       x82288 <= x82287;
       x82291 <= x82290;
       x82294 <= x82293;
       x82297 <= x82296;
       x82300 <= x82299;
       x82303 <= x82302;
       x82306 <= x82305;
       x82309 <= x82308;
       x82312 <= x82311;
       x82315 <= x82314;
       x82318 <= x82317;
       x82321 <= x82320;
       x82324 <= x82323;
       x82327 <= x82326;
       x82330 <= x82329;
       x82333 <= x82332;
       x82336 <= x82335;
       x82339 <= x82338;
       x82342 <= x82341;
       x82345 <= x82344;
       x82348 <= x82347;
       x82351 <= x82350;
       x82354 <= x82353;
       x82357 <= x82356;
       x82360 <= x82359;
       x82363 <= x82362;
       x82366 <= x82365;
       x82369 <= x82368;
       x82372 <= x82371;
       x82375 <= x82374;
       x82378 <= x82377;
       x82381 <= x82380;
       x82384 <= x82383;
       x82387 <= x82386;
       x82390 <= x82389;
       x82393 <= x82392;
       x82396 <= x82395;
       x82399 <= x82398;
       x82402 <= x82401;
       x82405 <= x82404;
       x82408 <= x82407;
       x82411 <= x82410;
       x82414 <= x82413;
       x82417 <= x82416;
       x82420 <= x82419;
       x82423 <= x82422;
       x82426 <= x82425;
       x82429 <= x82428;
       x82432 <= x82431;
       x82435 <= x82434;
       x82438 <= x82437;
       x82441 <= x82440;
       x82444 <= x82443;
       x82447 <= x82446;
       x82450 <= x82449;
       x82453 <= x82452;
       x82456 <= x82455;
       x82459 <= x82458;
       x82462 <= x82461;
       x82465 <= x82464;
       x82468 <= x82467;
       x82471 <= x82470;
       x82474 <= x82473;
       x82477 <= x82476;
       x82480 <= x82479;
       x82483 <= x82482;
       x82486 <= x82485;
       x82489 <= x82488;
       x82492 <= x82491;
       x82495 <= x82494;
       x82498 <= x82497;
       x82501 <= x82500;
       x82504 <= x82503;
       x82507 <= x82506;
       x82510 <= x82509;
       x82513 <= x82512;
       x82516 <= x82515;
       x82519 <= x82518;
       x82522 <= x82521;
       x82525 <= x82524;
       x82528 <= x82527;
       x82531 <= x82530;
       x82534 <= x82533;
       x82537 <= x82536;
       x82540 <= x82539;
       x82543 <= x82542;
       x82546 <= x82545;
       x82549 <= x82548;
       x82552 <= x82551;
       x82555 <= x82554;
       x82558 <= x82557;
       x82561 <= x82560;
       x82564 <= x82563;
       x82567 <= x82566;
       x82570 <= x82569;
       x82573 <= x82572;
       x82576 <= x82575;
       x82579 <= x82578;
       x82582 <= x82581;
       x82585 <= x82584;
       x82588 <= x82587;
       x82591 <= x82590;
       x82594 <= x82593;
       x82597 <= x82596;
       x82600 <= x82599;
       x82603 <= x82602;
       x82606 <= x82605;
       x82609 <= x82608;
       x82612 <= x82611;
       x82615 <= x82614;
       x82618 <= x82617;
       x82621 <= x82620;
       x82624 <= x82623;
       x82627 <= x82626;
       x82630 <= x82629;
       x82633 <= x82632;
       x82636 <= x82635;
       x82639 <= x82638;
       x82642 <= x82641;
       x82645 <= x82644;
       x82648 <= x82647;
       x82651 <= x82650;
       x82654 <= x82653;
       x82657 <= x82656;
       x82660 <= x82659;
       x82663 <= x82662;
       x82666 <= x82665;
       x82669 <= x82668;
       x82672 <= x82671;
       x82675 <= x82674;
       x82678 <= x82677;
       x82681 <= x82680;
       x82684 <= x82683;
       x82687 <= x82686;
       x82690 <= x82689;
       x82693 <= x82692;
       x82696 <= x82695;
       x82699 <= x82698;
       x82702 <= x82701;
       x82705 <= x82704;
       x82708 <= x82707;
       x82711 <= x82710;
       x82714 <= x82713;
       x82717 <= x82716;
       x82720 <= x82719;
       x82723 <= x82722;
       x82726 <= x82725;
       x82729 <= x82728;
       x82732 <= x82731;
       x82735 <= x82734;
       x82738 <= x82737;
       x82741 <= x82740;
       x82744 <= x82743;
       x82747 <= x82746;
       x82750 <= x82749;
       x82753 <= x82752;
       x82756 <= x82755;
       x82759 <= x82758;
       x82762 <= x82761;
       x82765 <= x82764;
       x82768 <= x82767;
       x82771 <= x82770;
       x82774 <= x82773;
       x82777 <= x82776;
       x82780 <= x82779;
       x82783 <= x82782;
       x82786 <= x82785;
       x82789 <= x82788;
       x82792 <= x82791;
       x82795 <= x82794;
       x82798 <= x82797;
       x82801 <= x82800;
       x82804 <= x82803;
       x82807 <= x82806;
       x82810 <= x82809;
       x82813 <= x82812;
       x82816 <= x82815;
       x82819 <= x82818;
       x82822 <= x82821;
       x82825 <= x82824;
       x82828 <= x82827;
       x82831 <= x82830;
       x82834 <= x82833;
       x82837 <= x82836;
       x82840 <= x82839;
       x82843 <= x82842;
       x82846 <= x82845;
       x82849 <= x82848;
       x82852 <= x82851;
       x82855 <= x82854;
       x82858 <= x82857;
       x82861 <= x82860;
       x82864 <= x82863;
       x82867 <= x82866;
       x82870 <= x82869;
       x82873 <= x82872;
       x82876 <= x82875;
       x82879 <= x82878;
       x82882 <= x82881;
       x82885 <= x82884;
       x82888 <= x82887;
       x82891 <= x82890;
       x82894 <= x82893;
       x82897 <= x82896;
       x82900 <= x82899;
       x82903 <= x82902;
       x82906 <= x82905;
       x82909 <= x82908;
       x82912 <= x82911;
       x82915 <= x82914;
       x82918 <= x82917;
       x82921 <= x82920;
       x82924 <= x82923;
       x82927 <= x82926;
       x82930 <= x82929;
       x82933 <= x82932;
       x82936 <= x82935;
       x82939 <= x82938;
       x82942 <= x82941;
       x82945 <= x82944;
       x82948 <= x82947;
       x82951 <= x82950;
       x82954 <= x82953;
       x82957 <= x82956;
       x82960 <= x82959;
       x82963 <= x82962;
       x82966 <= x82965;
       x82969 <= x82968;
       x82972 <= x82971;
       x82975 <= x82974;
       x82978 <= x82977;
       x82981 <= x82980;
       x82984 <= x82983;
       x82987 <= x82986;
       x82990 <= x82989;
       x82993 <= x82992;
       x82996 <= x82995;
       x82999 <= x82998;
       x83002 <= x83001;
       x83005 <= x83004;
       x83008 <= x83007;
       x83011 <= x83010;
       x83014 <= x83013;
       x83017 <= x83016;
       x83020 <= x83019;
       x83023 <= x83022;
       x83026 <= x83025;
       x83029 <= x83028;
       x83032 <= x83031;
       x83035 <= x83034;
       x83038 <= x83037;
       x83041 <= x83040;
       x83044 <= x83043;
       x83047 <= x83046;
       x83050 <= x83049;
       x83053 <= x83052;
       x83056 <= x83055;
       x83059 <= x83058;
       x83062 <= x83061;
       x83065 <= x83064;
       x83068 <= x83067;
       x83071 <= x83070;
       x83074 <= x83073;
       x83077 <= x83076;
       x83080 <= x83079;
       x83083 <= x83082;
       x83086 <= x83085;
       x83089 <= x83088;
       x83092 <= x83091;
       x83095 <= x83094;
       x83098 <= x83097;
       x83101 <= x83100;
       x83104 <= x83103;
       x83107 <= x83106;
       x83110 <= x83109;
       x83113 <= x83112;
       x83116 <= x83115;
       x83119 <= x83118;
       x83122 <= x83121;
       x83125 <= x83124;
       x83128 <= x83127;
       x83131 <= x83130;
       x83134 <= x83133;
       x83137 <= x83136;
       x83140 <= x83139;
       x83143 <= x83142;
       x83146 <= x83145;
       x83149 <= x83148;
       x83152 <= x83151;
       x83155 <= x83154;
       x83158 <= x83157;
       x83161 <= x83160;
       x83164 <= x83163;
       x83167 <= x83166;
       x83170 <= x83169;
       x83173 <= x83172;
       x83176 <= x83175;
       x83179 <= x83178;
       x83182 <= x83181;
       x83185 <= x83184;
       x83188 <= x83187;
       x83191 <= x83190;
       x83194 <= x83193;
       x83197 <= x83196;
       x83200 <= x83199;
       x83203 <= x83202;
       x83206 <= x83205;
       x83209 <= x83208;
       x83212 <= x83211;
       x83215 <= x83214;
       x83218 <= x83217;
       x83221 <= x83220;
       x83224 <= x83223;
       x83227 <= x83226;
       x83230 <= x83229;
       x83233 <= x83232;
       x83236 <= x83235;
       x83239 <= x83238;
       x83242 <= x83241;
       x83245 <= x83244;
       x83248 <= x83247;
       x83251 <= x83250;
       x83254 <= x83253;
       x83257 <= x83256;
       x83260 <= x83259;
       x83263 <= x83262;
       x83266 <= x83265;
       x83269 <= x83268;
       x83272 <= x83271;
       x83275 <= x83274;
       x83278 <= x83277;
       x83281 <= x83280;
       x83284 <= x83283;
       x83287 <= x83286;
       x83290 <= x83289;
       x83293 <= x83292;
       x83296 <= x83295;
       x83299 <= x83298;
       x83302 <= x83301;
       x83305 <= x83304;
       x83308 <= x83307;
       x83311 <= x83310;
       x83314 <= x83313;
       x83317 <= x83316;
       x83320 <= x83319;
       x83323 <= x83322;
       x83326 <= x83325;
       x83329 <= x83328;
       x83332 <= x83331;
       x83335 <= x83334;
       x83338 <= x83337;
       x83341 <= x83340;
       x83344 <= x83343;
       x83347 <= x83346;
       x83352 <= x83351;
       x83357 <= x83356;
       x83362 <= x83361;
       x83367 <= x83366;
       x83372 <= x83371;
       x83377 <= x83376;
       x83382 <= x83381;

       ram_q0 <= ram_array0[ram_qa0];
       if (ram_w0) ram_array0[ram_da0] <= ram_d0;
       ram_q1 <= ram_array1[ram_qa1];
       if (ram_w1) ram_array1[ram_da1] <= ram_d1;
       ram_q2 <= ram_array2[ram_qa2];
       if (ram_w2) ram_array2[ram_da2] <= ram_d2;
       ram_q3 <= ram_array3[ram_qa3];
       if (ram_w3) ram_array3[ram_da3] <= ram_d3;
    end
endmodule
